`timescale 1 ns / 1 ps

`include "settings.vh"

module RISCV_Rocket_Core_RV64G #(

    parameter integer C_DRAM_BASE             = `RISCV_DRAM_BASE,
    parameter integer C_DRAM_BITS             = `RISCV_DRAM_BITS,

    // AXI Master
    parameter integer C_M_AXI_ID_WIDTH        = 6,
    parameter integer C_M_AXI_ADDR_WIDTH      = 32,
    parameter integer C_M_AXI_DATA_WIDTH      = 64,

    // AXI Slave
    parameter integer C_S_AXI_ID_WIDTH        = 12,
    parameter integer C_S_AXI_DATA_WIDTH      = 32,
    parameter integer C_S_AXI_ADDR_WIDTH      = 32
)
(
    // AXI Master
    input  wire                                m_axi_aclk,
    input  wire                                m_axi_aresetn,
    output wire [C_M_AXI_ID_WIDTH-1 : 0]       m_axi_awid,
    output wire [C_M_AXI_ADDR_WIDTH-1 : 0]     m_axi_awaddr,
    output wire [7 : 0]                        m_axi_awlen,
    output wire [2 : 0]                        m_axi_awsize,
    output wire [1 : 0]                        m_axi_awburst,
    output wire                                m_axi_awlock,
    output wire [3 : 0]                        m_axi_awcache,
    output wire [2 : 0]                        m_axi_awprot,
    output wire [3 : 0]                        m_axi_awqos,
    output wire [3 : 0]                        m_axi_awregion,
    output wire                                m_axi_awvalid,
    input  wire                                m_axi_awready,
    output wire [C_M_AXI_DATA_WIDTH-1 : 0]     m_axi_wdata,
    output wire [C_M_AXI_DATA_WIDTH/8-1 : 0]   m_axi_wstrb,
    output wire                                m_axi_wlast,
    output wire                                m_axi_wvalid,
    input  wire                                m_axi_wready,
    input  wire [C_M_AXI_ID_WIDTH-1 : 0]       m_axi_bid,
    input  wire [1 : 0]                        m_axi_bresp,
    input  wire                                m_axi_bvalid,
    output wire                                m_axi_bready,
    output wire [C_M_AXI_ID_WIDTH-1 : 0]       m_axi_arid,
    output wire [C_M_AXI_ADDR_WIDTH-1 : 0]     m_axi_araddr,
    output wire [7 : 0]                        m_axi_arlen,
    output wire [2 : 0]                        m_axi_arsize,
    output wire [1 : 0]                        m_axi_arburst,
    output wire                                m_axi_arlock,
    output wire [3 : 0]                        m_axi_arcache,
    output wire [2 : 0]                        m_axi_arprot,
    output wire [3 : 0]                        m_axi_arqos,
    output wire [3 : 0]                        m_axi_arregion,
    output wire                                m_axi_arvalid,
    input  wire                                m_axi_arready,
    input  wire [C_M_AXI_ID_WIDTH-1 : 0]       m_axi_rid,
    input  wire [C_M_AXI_DATA_WIDTH-1 : 0]     m_axi_rdata,
    input  wire [1 : 0]                        m_axi_rresp,
    input  wire                                m_axi_rlast,
    input  wire                                m_axi_rvalid,
    output wire                                m_axi_rready,

    // AXI Slave
    input  wire                                s_axi_aclk,
    input  wire                                s_axi_aresetn,
    input  wire [C_S_AXI_ID_WIDTH-1 : 0]       s_axi_awid,
    input  wire [C_S_AXI_ADDR_WIDTH-1 : 0]     s_axi_awaddr,
    input  wire [7 : 0]                        s_axi_awlen,
    input  wire [2 : 0]                        s_axi_awsize,
    input  wire [1 : 0]                        s_axi_awburst,
    input  wire                                s_axi_awlock,
    input  wire [3 : 0]                        s_axi_awcache,
    input  wire [2 : 0]                        s_axi_awprot,
    input  wire [3 : 0]                        s_axi_awqos,
    input  wire [3 : 0]                        s_axi_awregion,
    input  wire                                s_axi_awvalid,
    output wire                                s_axi_awready,
    input  wire [C_S_AXI_DATA_WIDTH-1 : 0]     s_axi_wdata,
    input  wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] s_axi_wstrb,
    input  wire                                s_axi_wlast,
    input  wire                                s_axi_wvalid,
    output wire                                s_axi_wready,
    output wire [C_S_AXI_ID_WIDTH-1 : 0]       s_axi_bid,
    output wire [1 : 0]                        s_axi_bresp,
    output wire                                s_axi_bvalid,
    input  wire                                s_axi_bready,
    input  wire [C_S_AXI_ID_WIDTH-1 : 0]       s_axi_arid,
    input  wire [C_S_AXI_ADDR_WIDTH-1 : 0]     s_axi_araddr,
    input  wire [7 : 0]                        s_axi_arlen,
    input  wire [2 : 0]                        s_axi_arsize,
    input  wire [1 : 0]                        s_axi_arburst,
    input  wire                                s_axi_arlock,
    input  wire [3 : 0]                        s_axi_arcache,
    input  wire [2 : 0]                        s_axi_arprot,
    input  wire [3 : 0]                        s_axi_arqos,
    input  wire [3 : 0]                        s_axi_arregion,
    input  wire                                s_axi_arvalid,
    output wire                                s_axi_arready,
    output wire [C_S_AXI_ID_WIDTH-1 : 0]       s_axi_rid,
    output wire [C_S_AXI_DATA_WIDTH-1 : 0]     s_axi_rdata,
    output wire [1 : 0]                        s_axi_rresp,
    output wire                                s_axi_rlast,
    output wire                                s_axi_rvalid,
    input  wire                                s_axi_rready
);

    RISCV_Rocket_Core_RV64G_AXI #(
        .C_DRAM_BASE            (C_DRAM_BASE),
        .C_DRAM_BITS            (C_DRAM_BITS),

        // AXI Master
        .C_M_AXI_ID_WIDTH       (C_M_AXI_ID_WIDTH),
        .C_M_AXI_ADDR_WIDTH     (C_M_AXI_ADDR_WIDTH),
        .C_M_AXI_DATA_WIDTH     (C_M_AXI_DATA_WIDTH),
        
        // AXI Slave            
        .C_S_AXI_ID_WIDTH       (C_S_AXI_ID_WIDTH),
        .C_S_AXI_DATA_WIDTH     (C_S_AXI_DATA_WIDTH),
        .C_S_AXI_ADDR_WIDTH     (C_S_AXI_ADDR_WIDTH)
    )
    RISCV_Rocket_Core_RV64G_AXI_inst (
        // AXI Master
        .M_AXI_ACLK     (m_axi_aclk),
        .M_AXI_ARESETN  (m_axi_aresetn),
        .M_AXI_AWID     (m_axi_awid),
        .M_AXI_AWADDR   (m_axi_awaddr),
        .M_AXI_AWLEN    (m_axi_awlen),
        .M_AXI_AWSIZE   (m_axi_awsize),
        .M_AXI_AWREGION (m_axi_awregion),
        .M_AXI_AWBURST  (m_axi_awburst),
        .M_AXI_AWLOCK   (m_axi_awlock),
        .M_AXI_AWCACHE  (m_axi_awcache),
        .M_AXI_AWPROT   (m_axi_awprot),
        .M_AXI_AWQOS    (m_axi_awqos),
        .M_AXI_AWVALID  (m_axi_awvalid),
        .M_AXI_AWREADY  (m_axi_awready),
        .M_AXI_WDATA    (m_axi_wdata),
        .M_AXI_WSTRB    (m_axi_wstrb),
        .M_AXI_WLAST    (m_axi_wlast),
        .M_AXI_WVALID   (m_axi_wvalid),
        .M_AXI_WREADY   (m_axi_wready),
        .M_AXI_BID      (m_axi_bid),
        .M_AXI_BRESP    (m_axi_bresp),
        .M_AXI_BVALID   (m_axi_bvalid),
        .M_AXI_BREADY   (m_axi_bready),
        .M_AXI_ARID     (m_axi_arid),
        .M_AXI_ARADDR   (m_axi_araddr),
        .M_AXI_ARLEN    (m_axi_arlen),
        .M_AXI_ARSIZE   (m_axi_arsize),
        .M_AXI_ARREGION (m_axi_arregion),
        .M_AXI_ARBURST  (m_axi_arburst),
        .M_AXI_ARLOCK   (m_axi_arlock),
        .M_AXI_ARCACHE  (m_axi_arcache),
        .M_AXI_ARPROT   (m_axi_arprot),
        .M_AXI_ARQOS    (m_axi_arqos),
        .M_AXI_ARVALID  (m_axi_arvalid),
        .M_AXI_ARREADY  (m_axi_arready),
        .M_AXI_RID      (m_axi_rid),
        .M_AXI_RDATA    (m_axi_rdata),
        .M_AXI_RRESP    (m_axi_rresp),
        .M_AXI_RLAST    (m_axi_rlast),
        .M_AXI_RVALID   (m_axi_rvalid),
        .M_AXI_RREADY   (m_axi_rready),

        // AXI Slave
        .S_AXI_ACLK     (s_axi_aclk),
        .S_AXI_ARESETN  (s_axi_aresetn),
        .S_AXI_AWID     (s_axi_awid),
        .S_AXI_AWADDR   (s_axi_awaddr),
        .S_AXI_AWLEN    (s_axi_awlen),
        .S_AXI_AWSIZE   (s_axi_awsize),
        .S_AXI_AWBURST  (s_axi_awburst),
        .S_AXI_AWLOCK   (s_axi_awlock),
        .S_AXI_AWCACHE  (),
        .S_AXI_AWPROT   (s_axi_awprot),
        .S_AXI_AWQOS    (s_axi_awqos),
        .S_AXI_AWREGION (s_axi_awregion),
        .S_AXI_AWVALID  (s_axi_awvalid),
        .S_AXI_AWREADY  (s_axi_awready),
        .S_AXI_WDATA    (s_axi_wdata),
        .S_AXI_WSTRB    (s_axi_wstrb),
        .S_AXI_WLAST    (s_axi_wlast),
        .S_AXI_WVALID   (s_axi_wvalid),
        .S_AXI_WREADY   (s_axi_wready),
        .S_AXI_BID      (s_axi_bid),
        .S_AXI_BRESP    (2'b00),
        .S_AXI_BVALID   (s_axi_bvalid),
        .S_AXI_BREADY   (s_axi_bready),
        .S_AXI_ARID     (s_axi_arid),
        .S_AXI_ARADDR   (s_axi_araddr),
        .S_AXI_ARLEN    (s_axi_arlen),
        .S_AXI_ARSIZE   (s_axi_arsize),
        .S_AXI_ARBURST  (s_axi_arburst),
        .S_AXI_ARLOCK   (s_axi_arlock),
        .S_AXI_ARCACHE  (),
        .S_AXI_ARPROT   (s_axi_arprot),
        .S_AXI_ARQOS    (s_axi_arqos),
        .S_AXI_ARREGION (s_axi_arregion),
        .S_AXI_ARVALID  (s_axi_arvalid),
        .S_AXI_ARREADY  (s_axi_arready),
        .S_AXI_RID      (s_axi_rid),
        .S_AXI_RDATA    (s_axi_rdata),
        .S_AXI_RRESP    (),
        .S_AXI_RLAST    (s_axi_rlast),
        .S_AXI_RVALID   (s_axi_rvalid),
        .S_AXI_RREADY   (s_axi_rready)
    );

endmodule
