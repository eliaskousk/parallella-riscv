module Htif(
  input   clk,
  input   reset,
  output  io_host_clk,
  output  io_host_clk_edge,
  output  io_host_in_ready,
  input   io_host_in_valid,
  input  [15:0] io_host_in_bits,
  input   io_host_out_ready,
  output  io_host_out_valid,
  output [15:0] io_host_out_bits,
  output  io_cpu_0_reset,
  output  io_cpu_0_id,
  input   io_cpu_0_csr_req_ready,
  output  io_cpu_0_csr_req_valid,
  output  io_cpu_0_csr_req_bits_rw,
  output [11:0] io_cpu_0_csr_req_bits_addr,
  output [63:0] io_cpu_0_csr_req_bits_data,
  output  io_cpu_0_csr_resp_ready,
  input   io_cpu_0_csr_resp_valid,
  input  [63:0] io_cpu_0_csr_resp_bits,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_scr_req_ready,
  output  io_scr_req_valid,
  output  io_scr_req_bits_rw,
  output [5:0] io_scr_req_bits_addr,
  output [63:0] io_scr_req_bits_data,
  output  io_scr_resp_ready,
  input   io_scr_resp_valid,
  input  [63:0] io_scr_resp_bits
);
  reg [14:0] rx_count;
  reg [31:0] GEN_15;
  reg [63:0] rx_shifter;
  reg [63:0] GEN_16;
  wire [47:0] T_1195;
  wire [63:0] rx_shifter_in;
  wire [3:0] next_cmd;
  reg [3:0] cmd;
  reg [31:0] GEN_35;
  reg [11:0] size;
  reg [31:0] GEN_36;
  reg [8:0] pos;
  reg [31:0] GEN_37;
  reg [7:0] seqno;
  reg [31:0] GEN_38;
  reg [39:0] addr;
  reg [63:0] GEN_39;
  wire  T_1201;
  wire [14:0] GEN_50;
  wire [15:0] T_1203;
  wire [14:0] T_1204;
  wire [14:0] GEN_51;
  wire  T_1206;
  wire [11:0] T_1207;
  wire [8:0] T_1208;
  wire [7:0] T_1209;
  wire [39:0] T_1210;
  wire [3:0] GEN_0;
  wire [11:0] GEN_1;
  wire [8:0] GEN_2;
  wire [7:0] GEN_3;
  wire [39:0] GEN_4;
  wire [63:0] GEN_5;
  wire [14:0] GEN_6;
  wire [3:0] GEN_7;
  wire [11:0] GEN_8;
  wire [8:0] GEN_9;
  wire [7:0] GEN_10;
  wire [39:0] GEN_11;
  wire [12:0] rx_word_count;
  wire [1:0] T_1211;
  wire [1:0] T_1212;
  wire [1:0] GEN_52;
  wire  T_1214;
  wire  rx_word_done;
  reg [63:0] packet_ram [0:7];
  reg [63:0] GEN_55;
  wire [63:0] packet_ram_csr_wdata_data;
  wire [2:0] packet_ram_csr_wdata_addr;
  wire  packet_ram_csr_wdata_en;
  wire [63:0] packet_ram_mem_req_data_data;
  wire [2:0] packet_ram_mem_req_data_addr;
  wire  packet_ram_mem_req_data_en;
  wire [63:0] packet_ram_T_1725_data;
  wire [2:0] packet_ram_T_1725_addr;
  wire  packet_ram_T_1725_en;
  wire [63:0] packet_ram_T_1222_data;
  wire [2:0] packet_ram_T_1222_addr;
  wire  packet_ram_T_1222_mask;
  wire  packet_ram_T_1222_en;
  wire [63:0] packet_ram_T_1345_data;
  wire [2:0] packet_ram_T_1345_addr;
  wire  packet_ram_T_1345_mask;
  wire  packet_ram_T_1345_en;
  wire  T_1217;
  wire [2:0] T_1218;
  wire [2:0] GEN_53;
  wire [3:0] T_1220;
  wire [2:0] T_1221;
  wire [11:0] csr_addr;
  wire [1:0] csr_coreid;
  wire [2:0] T_1225;
  wire [2:0] GEN_54;
  wire  T_1227;
  wire [2:0] T_1228;
  wire  T_1230;
  wire  bad_mem_packet;
  wire [3:0] GEN_56;
  wire  T_1231;
  wire [3:0] GEN_57;
  wire  T_1232;
  wire  T_1233;
  wire [3:0] GEN_58;
  wire  T_1234;
  wire [3:0] GEN_59;
  wire  T_1235;
  wire  T_1236;
  wire [11:0] GEN_60;
  wire  T_1238;
  wire  T_1240;
  wire  nack;
  reg [14:0] tx_count;
  reg [31:0] GEN_61;
  wire [1:0] tx_subword_count;
  wire [12:0] tx_word_count;
  wire [2:0] T_1242;
  wire [3:0] T_1244;
  wire [2:0] packet_ram_raddr;
  wire  T_1245;
  wire [15:0] T_1247;
  wire [14:0] T_1248;
  wire [14:0] GEN_17;
  wire [12:0] GEN_63;
  wire  T_1250;
  wire  T_1251;
  wire  T_1252;
  wire  T_1253;
  wire [12:0] GEN_66;
  wire  T_1254;
  wire  T_1257;
  wire  T_1258;
  wire  T_1259;
  wire  rx_done;
  wire  T_1261;
  wire  T_1264;
  wire  T_1266;
  wire  T_1267;
  wire [11:0] tx_size;
  wire [1:0] T_1269;
  wire  T_1271;
  wire  T_1272;
  wire [12:0] GEN_72;
  wire  T_1273;
  wire  T_1275;
  wire [2:0] T_1276;
  wire  T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  tx_done;
  reg [2:0] state;
  reg [31:0] GEN_62;
  wire  T_1282;
  wire  T_1283;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  reg [2:0] cnt;
  reg [31:0] GEN_64;
  wire  T_1289;
  wire [3:0] T_1291;
  wire [2:0] T_1292;
  wire [2:0] GEN_18;
  wire  cnt_done;
  wire [3:0] rx_cmd;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire  T_1298;
  wire  T_1299;
  wire  T_1300;
  wire  T_1301;
  wire [2:0] T_1302;
  wire [2:0] T_1303;
  wire [2:0] T_1304;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire  T_1306;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire  T_1307;
  wire  T_1308;
  wire [8:0] GEN_82;
  wire  T_1311;
  wire  T_1312;
  wire [2:0] T_1313;
  wire [9:0] T_1315;
  wire [8:0] T_1316;
  wire [39:0] GEN_84;
  wire [40:0] T_1318;
  wire [39:0] T_1319;
  wire [2:0] GEN_24;
  wire [8:0] GEN_25;
  wire [39:0] GEN_26;
  wire  T_1321;
  wire [2:0] GEN_27;
  wire [8:0] GEN_28;
  wire [39:0] GEN_29;
  wire  T_1333;
  wire  T_1334;
  wire [14:0] GEN_30;
  wire [14:0] GEN_31;
  wire [8:0] GEN_91;
  wire  T_1340;
  wire  T_1341;
  wire [2:0] T_1342;
  wire [14:0] GEN_32;
  wire [14:0] GEN_33;
  wire [2:0] GEN_34;
  wire [36:0] init_addr;
  wire  T_1349;
  wire [7:0] GEN_93;
  wire [7:0] T_1378;
  wire [8:0] T_1426;
  wire [11:0] T_1444;
  wire [25:0] T_1482_addr_block;
  wire [1:0] T_1482_client_xact_id;
  wire [2:0] T_1482_addr_beat;
  wire  T_1482_is_builtin_type;
  wire [2:0] T_1482_a_type;
  wire [11:0] T_1482_union;
  wire [63:0] T_1482_data;
  wire [25:0] T_1621_addr_block;
  wire [1:0] T_1621_client_xact_id;
  wire [2:0] T_1621_addr_beat;
  wire  T_1621_is_builtin_type;
  wire [2:0] T_1621_a_type;
  wire [11:0] T_1621_union;
  wire [63:0] T_1621_data;
  wire [25:0] T_1652_addr_block;
  wire [1:0] T_1652_client_xact_id;
  wire [2:0] T_1652_addr_beat;
  wire  T_1652_is_builtin_type;
  wire [2:0] T_1652_a_type;
  wire [11:0] T_1652_union;
  wire [63:0] T_1652_data;
  reg [63:0] csrReadData;
  reg [63:0] GEN_65;
  reg  T_1686;
  reg [31:0] GEN_67;
  wire  T_1688;
  wire  T_1689;
  wire  T_1690;
  wire [11:0] GEN_95;
  wire  T_1692;
  wire  T_1693;
  wire  T_1695;
  wire [2:0] GEN_40;
  wire  T_1699;
  wire  T_1700;
  wire  T_1702;
  wire  GEN_41;
  wire  GEN_42;
  wire [63:0] GEN_43;
  wire [2:0] GEN_44;
  wire  T_1704;
  wire  T_1705;
  wire [63:0] GEN_45;
  wire [2:0] GEN_46;
  wire [1:0] T_1707;
  wire  T_1709;
  wire  T_1710;
  wire [5:0] T_1711;
  wire  T_1714;
  wire [2:0] GEN_47;
  wire  T_1716;
  wire [63:0] GEN_48;
  wire [2:0] GEN_49;
  wire [2:0] tx_cmd;
  wire [3:0] tx_cmd_ext;
  wire [15:0] T_1718;
  wire [47:0] T_1719;
  wire [63:0] tx_header;
  wire  T_1721;
  wire [63:0] T_1726;
  wire [63:0] tx_data;
  wire [5:0] T_1731;
  wire [63:0] T_1732;
  reg  GEN_12;
  reg [31:0] GEN_68;
  reg  GEN_13;
  reg [31:0] GEN_69;
  reg  GEN_14;
  reg [31:0] GEN_70;
  assign io_host_clk = GEN_12;
  assign io_host_clk_edge = GEN_13;
  assign io_host_in_ready = T_1295;
  assign io_host_out_valid = T_1333;
  assign io_host_out_bits = T_1732[15:0];
  assign io_cpu_0_reset = T_1686;
  assign io_cpu_0_id = GEN_14;
  assign io_cpu_0_csr_req_valid = T_1693;
  assign io_cpu_0_csr_req_bits_rw = T_1235;
  assign io_cpu_0_csr_req_bits_addr = csr_addr;
  assign io_cpu_0_csr_req_bits_data = packet_ram_csr_wdata_data;
  assign io_cpu_0_csr_resp_ready = 1'h1;
  assign io_mem_acquire_valid = T_1349;
  assign io_mem_acquire_bits_addr_block = T_1652_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1652_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1652_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1652_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1652_a_type;
  assign io_mem_acquire_bits_union = T_1652_union;
  assign io_mem_acquire_bits_data = T_1652_data;
  assign io_mem_grant_ready = 1'h1;
  assign io_scr_req_valid = T_1710;
  assign io_scr_req_bits_rw = T_1235;
  assign io_scr_req_bits_addr = T_1711;
  assign io_scr_req_bits_data = packet_ram_csr_wdata_data;
  assign io_scr_resp_ready = 1'h1;
  assign T_1195 = rx_shifter[63:16];
  assign rx_shifter_in = {io_host_in_bits,T_1195};
  assign next_cmd = rx_shifter_in[3:0];
  assign T_1201 = io_host_in_valid & io_host_in_ready;
  assign GEN_50 = {{14'd0}, 1'h1};
  assign T_1203 = rx_count + GEN_50;
  assign T_1204 = T_1203[14:0];
  assign GEN_51 = {{13'd0}, 2'h3};
  assign T_1206 = rx_count == GEN_51;
  assign T_1207 = rx_shifter_in[15:4];
  assign T_1208 = rx_shifter_in[15:7];
  assign T_1209 = rx_shifter_in[23:16];
  assign T_1210 = rx_shifter_in[63:24];
  assign GEN_0 = T_1206 ? next_cmd : cmd;
  assign GEN_1 = T_1206 ? T_1207 : size;
  assign GEN_2 = T_1206 ? T_1208 : pos;
  assign GEN_3 = T_1206 ? T_1209 : seqno;
  assign GEN_4 = T_1206 ? T_1210 : addr;
  assign GEN_5 = T_1201 ? rx_shifter_in : rx_shifter;
  assign GEN_6 = T_1201 ? T_1204 : rx_count;
  assign GEN_7 = T_1201 ? GEN_0 : cmd;
  assign GEN_8 = T_1201 ? GEN_1 : size;
  assign GEN_9 = T_1201 ? GEN_2 : pos;
  assign GEN_10 = T_1201 ? GEN_3 : seqno;
  assign GEN_11 = T_1201 ? GEN_4 : addr;
  assign rx_word_count = rx_count[14:2];
  assign T_1211 = rx_count[1:0];
  assign T_1212 = ~ T_1211;
  assign GEN_52 = {{1'd0}, 1'h0};
  assign T_1214 = T_1212 == GEN_52;
  assign rx_word_done = io_host_in_valid & T_1214;
  assign packet_ram_csr_wdata_addr = {{2'd0}, 1'h0};
  assign packet_ram_csr_wdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign packet_ram_csr_wdata_data = packet_ram[packet_ram_csr_wdata_addr];
  `else
  assign packet_ram_csr_wdata_data = packet_ram_csr_wdata_addr >= 4'h8 ? $random : packet_ram[packet_ram_csr_wdata_addr];
  `endif
  assign packet_ram_mem_req_data_addr = cnt;
  assign packet_ram_mem_req_data_en = 1'h1;
  `ifdef SYNTHESIS
  assign packet_ram_mem_req_data_data = packet_ram[packet_ram_mem_req_data_addr];
  `else
  assign packet_ram_mem_req_data_data = packet_ram_mem_req_data_addr >= 4'h8 ? $random : packet_ram[packet_ram_mem_req_data_addr];
  `endif
  assign packet_ram_T_1725_addr = packet_ram_raddr;
  assign packet_ram_T_1725_en = 1'h1;
  `ifdef SYNTHESIS
  assign packet_ram_T_1725_data = packet_ram[packet_ram_T_1725_addr];
  `else
  assign packet_ram_T_1725_data = packet_ram_T_1725_addr >= 4'h8 ? $random : packet_ram[packet_ram_T_1725_addr];
  `endif
  assign packet_ram_T_1222_data = rx_shifter_in;
  assign packet_ram_T_1222_addr = T_1221;
  assign packet_ram_T_1222_mask = T_1217;
  assign packet_ram_T_1222_en = T_1217;
  assign packet_ram_T_1345_data = io_mem_grant_bits_data;
  assign packet_ram_T_1345_addr = io_mem_grant_bits_addr_beat;
  assign packet_ram_T_1345_mask = T_1285;
  assign packet_ram_T_1345_en = T_1285;
  assign T_1217 = rx_word_done & io_host_in_ready;
  assign T_1218 = rx_word_count[2:0];
  assign GEN_53 = {{2'd0}, 1'h1};
  assign T_1220 = T_1218 - GEN_53;
  assign T_1221 = T_1220[2:0];
  assign csr_addr = addr[11:0];
  assign csr_coreid = addr[21:20];
  assign T_1225 = size[2:0];
  assign GEN_54 = {{2'd0}, 1'h0};
  assign T_1227 = T_1225 != GEN_54;
  assign T_1228 = addr[2:0];
  assign T_1230 = T_1228 != GEN_54;
  assign bad_mem_packet = T_1227 | T_1230;
  assign GEN_56 = {{1'd0}, 3'h0};
  assign T_1231 = cmd == GEN_56;
  assign GEN_57 = {{1'd0}, 3'h1};
  assign T_1232 = cmd == GEN_57;
  assign T_1233 = T_1231 | T_1232;
  assign GEN_58 = {{1'd0}, 3'h2};
  assign T_1234 = cmd == GEN_58;
  assign GEN_59 = {{1'd0}, 3'h3};
  assign T_1235 = cmd == GEN_59;
  assign T_1236 = T_1234 | T_1235;
  assign GEN_60 = {{11'd0}, 1'h1};
  assign T_1238 = size != GEN_60;
  assign T_1240 = T_1236 ? T_1238 : 1'h1;
  assign nack = T_1233 ? bad_mem_packet : T_1240;
  assign tx_subword_count = tx_count[1:0];
  assign tx_word_count = tx_count[14:2];
  assign T_1242 = tx_word_count[2:0];
  assign T_1244 = T_1242 - GEN_53;
  assign packet_ram_raddr = T_1244[2:0];
  assign T_1245 = io_host_out_valid & io_host_out_ready;
  assign T_1247 = tx_count + GEN_50;
  assign T_1248 = T_1247[14:0];
  assign GEN_17 = T_1245 ? T_1248 : tx_count;
  assign GEN_63 = {{12'd0}, 1'h0};
  assign T_1250 = rx_word_count == GEN_63;
  assign T_1251 = next_cmd != GEN_57;
  assign T_1252 = next_cmd != GEN_59;
  assign T_1253 = T_1251 & T_1252;
  assign GEN_66 = {{1'd0}, size};
  assign T_1254 = rx_word_count == GEN_66;
  assign T_1257 = T_1218 == GEN_54;
  assign T_1258 = T_1254 | T_1257;
  assign T_1259 = T_1250 ? T_1253 : T_1258;
  assign rx_done = rx_word_done & T_1259;
  assign T_1261 = nack == 1'h0;
  assign T_1264 = T_1231 | T_1234;
  assign T_1266 = T_1264 | T_1235;
  assign T_1267 = T_1261 & T_1266;
  assign tx_size = T_1267 ? size : {{11'd0}, 1'h0};
  assign T_1269 = ~ tx_subword_count;
  assign T_1271 = T_1269 == GEN_52;
  assign T_1272 = io_host_out_ready & T_1271;
  assign GEN_72 = {{1'd0}, tx_size};
  assign T_1273 = tx_word_count == GEN_72;
  assign T_1275 = tx_word_count > GEN_63;
  assign T_1276 = ~ packet_ram_raddr;
  assign T_1278 = T_1276 == GEN_54;
  assign T_1279 = T_1275 & T_1278;
  assign T_1280 = T_1273 | T_1279;
  assign tx_done = T_1272 & T_1280;
  assign T_1282 = state == 3'h4;
  assign T_1283 = T_1282 & io_mem_acquire_ready;
  assign T_1284 = state == 3'h5;
  assign T_1285 = T_1284 & io_mem_grant_valid;
  assign T_1286 = T_1283 | T_1285;
  assign T_1289 = cnt == 3'h7;
  assign T_1291 = cnt + GEN_53;
  assign T_1292 = T_1291[2:0];
  assign GEN_18 = T_1286 ? T_1292 : cnt;
  assign cnt_done = T_1286 & T_1289;
  assign rx_cmd = T_1250 ? next_cmd : cmd;
  assign T_1295 = state == 3'h0;
  assign T_1296 = T_1295 & rx_done;
  assign T_1297 = rx_cmd == GEN_56;
  assign T_1298 = rx_cmd == GEN_57;
  assign T_1299 = rx_cmd == GEN_58;
  assign T_1300 = rx_cmd == GEN_59;
  assign T_1301 = T_1299 | T_1300;
  assign T_1302 = T_1301 ? 3'h1 : 3'h7;
  assign T_1303 = T_1298 ? 3'h4 : T_1302;
  assign T_1304 = T_1297 ? 3'h3 : T_1303;
  assign GEN_19 = T_1296 ? T_1304 : state;
  assign GEN_20 = cnt_done ? 3'h6 : GEN_19;
  assign GEN_21 = T_1282 ? GEN_20 : GEN_19;
  assign T_1306 = state == 3'h3;
  assign GEN_22 = io_mem_acquire_ready ? 3'h5 : GEN_21;
  assign GEN_23 = T_1306 ? GEN_22 : GEN_21;
  assign T_1307 = state == 3'h6;
  assign T_1308 = T_1307 & io_mem_grant_valid;
  assign GEN_82 = {{8'd0}, 1'h1};
  assign T_1311 = pos == GEN_82;
  assign T_1312 = T_1231 | T_1311;
  assign T_1313 = T_1312 ? 3'h7 : 3'h0;
  assign T_1315 = pos - GEN_82;
  assign T_1316 = T_1315[8:0];
  assign GEN_84 = {{36'd0}, 4'h8};
  assign T_1318 = addr + GEN_84;
  assign T_1319 = T_1318[39:0];
  assign GEN_24 = T_1308 ? T_1313 : GEN_23;
  assign GEN_25 = T_1308 ? T_1316 : GEN_9;
  assign GEN_26 = T_1308 ? T_1319 : GEN_11;
  assign T_1321 = T_1284 & cnt_done;
  assign GEN_27 = T_1321 ? T_1313 : GEN_24;
  assign GEN_28 = T_1321 ? T_1316 : GEN_25;
  assign GEN_29 = T_1321 ? T_1319 : GEN_26;
  assign T_1333 = state == 3'h7;
  assign T_1334 = T_1333 & tx_done;
  assign GEN_30 = T_1273 ? {{14'd0}, 1'h0} : GEN_6;
  assign GEN_31 = T_1273 ? {{14'd0}, 1'h0} : GEN_17;
  assign GEN_91 = {{8'd0}, 1'h0};
  assign T_1340 = pos != GEN_91;
  assign T_1341 = T_1231 & T_1340;
  assign T_1342 = T_1341 ? 3'h3 : 3'h0;
  assign GEN_32 = T_1334 ? GEN_30 : GEN_6;
  assign GEN_33 = T_1334 ? GEN_31 : GEN_17;
  assign GEN_34 = T_1334 ? T_1342 : GEN_27;
  assign init_addr = addr[39:3];
  assign T_1349 = T_1306 | T_1282;
  assign GEN_93 = $signed(8'hff);
  assign T_1378 = $unsigned(GEN_93);
  assign T_1426 = {T_1378,1'h1};
  assign T_1444 = 1'h1 ? {{3'd0}, T_1426} : 12'h0;
  assign T_1482_addr_block = init_addr[25:0];
  assign T_1482_client_xact_id = {{1'd0}, 1'h0};
  assign T_1482_addr_beat = cnt;
  assign T_1482_is_builtin_type = 1'h1;
  assign T_1482_a_type = 3'h3;
  assign T_1482_union = T_1444;
  assign T_1482_data = packet_ram_mem_req_data_data;
  assign T_1621_addr_block = init_addr[25:0];
  assign T_1621_client_xact_id = {{1'd0}, 1'h0};
  assign T_1621_addr_beat = {{2'd0}, 1'h0};
  assign T_1621_is_builtin_type = 1'h1;
  assign T_1621_a_type = 3'h1;
  assign T_1621_union = 12'h1c1;
  assign T_1621_data = {{63'd0}, 1'h0};
  assign T_1652_addr_block = T_1232 ? T_1482_addr_block : T_1621_addr_block;
  assign T_1652_client_xact_id = T_1232 ? T_1482_client_xact_id : T_1621_client_xact_id;
  assign T_1652_addr_beat = T_1232 ? T_1482_addr_beat : T_1621_addr_beat;
  assign T_1652_is_builtin_type = T_1232 ? T_1482_is_builtin_type : T_1621_is_builtin_type;
  assign T_1652_a_type = T_1232 ? T_1482_a_type : T_1621_a_type;
  assign T_1652_union = T_1232 ? T_1482_union : T_1621_union;
  assign T_1652_data = T_1232 ? T_1482_data : T_1621_data;
  assign T_1688 = csr_coreid == GEN_52;
  assign T_1689 = state == 3'h1;
  assign T_1690 = T_1689 & T_1688;
  assign GEN_95 = {{1'd0}, 11'h7c2};
  assign T_1692 = csr_addr != GEN_95;
  assign T_1693 = T_1690 & T_1692;
  assign T_1695 = io_cpu_0_csr_req_ready & io_cpu_0_csr_req_valid;
  assign GEN_40 = T_1695 ? 3'h2 : GEN_34;
  assign T_1699 = csr_addr == GEN_95;
  assign T_1700 = T_1690 & T_1699;
  assign T_1702 = packet_ram_csr_wdata_data[0];
  assign GEN_41 = T_1235 ? T_1702 : T_1686;
  assign GEN_42 = T_1700 ? GEN_41 : T_1686;
  assign GEN_43 = T_1700 ? {{63'd0}, T_1686} : csrReadData;
  assign GEN_44 = T_1700 ? 3'h7 : GEN_40;
  assign T_1704 = state == 3'h2;
  assign T_1705 = T_1704 & io_cpu_0_csr_resp_valid;
  assign GEN_45 = T_1705 ? io_cpu_0_csr_resp_bits : GEN_43;
  assign GEN_46 = T_1705 ? 3'h7 : GEN_44;
  assign T_1707 = ~ csr_coreid;
  assign T_1709 = T_1707 == GEN_52;
  assign T_1710 = T_1689 & T_1709;
  assign T_1711 = addr[5:0];
  assign T_1714 = io_scr_req_ready & io_scr_req_valid;
  assign GEN_47 = T_1714 ? 3'h2 : GEN_46;
  assign T_1716 = T_1704 & io_scr_resp_valid;
  assign GEN_48 = T_1716 ? io_scr_resp_bits : GEN_45;
  assign GEN_49 = T_1716 ? 3'h7 : GEN_47;
  assign tx_cmd = nack ? 3'h5 : 3'h4;
  assign tx_cmd_ext = {1'h0,tx_cmd};
  assign T_1718 = {tx_size,tx_cmd_ext};
  assign T_1719 = {addr,seqno};
  assign tx_header = {T_1719,T_1718};
  assign T_1721 = tx_word_count == GEN_63;
  assign T_1726 = T_1236 ? csrReadData : packet_ram_T_1725_data;
  assign tx_data = T_1721 ? tx_header : T_1726;
  assign T_1731 = {tx_subword_count,4'h0};
  assign T_1732 = tx_data >> T_1731;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  rx_count = GEN_15[14:0];
  GEN_16 = {2{$random}};
  rx_shifter = GEN_16[63:0];
  GEN_35 = {1{$random}};
  cmd = GEN_35[3:0];
  GEN_36 = {1{$random}};
  size = GEN_36[11:0];
  GEN_37 = {1{$random}};
  pos = GEN_37[8:0];
  GEN_38 = {1{$random}};
  seqno = GEN_38[7:0];
  GEN_39 = {2{$random}};
  addr = GEN_39[39:0];
  GEN_55 = {2{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    packet_ram[initvar] = GEN_55[63:0];
  GEN_61 = {1{$random}};
  tx_count = GEN_61[14:0];
  GEN_62 = {1{$random}};
  state = GEN_62[2:0];
  GEN_64 = {1{$random}};
  cnt = GEN_64[2:0];
  GEN_65 = {2{$random}};
  csrReadData = GEN_65[63:0];
  GEN_67 = {1{$random}};
  T_1686 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  GEN_12 = GEN_68[0:0];
  GEN_69 = {1{$random}};
  GEN_13 = GEN_69[0:0];
  GEN_70 = {1{$random}};
  GEN_14 = GEN_70[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rx_count <= 15'h0;
    end else begin
      rx_count <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      rx_shifter <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      cmd <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      size <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      pos <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      seqno <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      addr <= GEN_29;
    end
    if(packet_ram_T_1222_en & packet_ram_T_1222_mask) begin
      packet_ram[packet_ram_T_1222_addr] <= packet_ram_T_1222_data;
    end
    if(packet_ram_T_1345_en & packet_ram_T_1345_mask) begin
      packet_ram[packet_ram_T_1345_addr] <= packet_ram_T_1345_data;
    end
    if(reset) begin
      tx_count <= 15'h0;
    end else begin
      tx_count <= GEN_33;
    end
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_49;
    end
    if(reset) begin
      cnt <= 3'h0;
    end else begin
      cnt <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      csrReadData <= GEN_48;
    end
    if(reset) begin
      T_1686 <= 1'h1;
    end else begin
      T_1686 <= GEN_42;
    end
  end
endmodule
module Queue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_header_src,
  input  [2:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input   io_enq_bits_payload_is_builtin_type,
  input  [2:0] io_enq_bits_payload_a_type,
  input  [11:0] io_enq_bits_payload_union,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_header_src,
  output [2:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_addr_beat,
  output  io_deq_bits_payload_is_builtin_type,
  output [2:0] io_deq_bits_payload_a_type,
  output [11:0] io_deq_bits_payload_union,
  output [63:0] io_deq_bits_payload_data,
  output  io_count
);
  reg [2:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [2:0] ram_header_src_T_1160_data;
  wire  ram_header_src_T_1160_addr;
  wire  ram_header_src_T_1160_mask;
  wire  ram_header_src_T_1160_en;
  reg [2:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [2:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [2:0] ram_header_dst_T_1160_data;
  wire  ram_header_dst_T_1160_addr;
  wire  ram_header_dst_T_1160_mask;
  wire  ram_header_dst_T_1160_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1294_data;
  wire  ram_payload_addr_block_T_1294_addr;
  wire  ram_payload_addr_block_T_1294_en;
  wire [25:0] ram_payload_addr_block_T_1160_data;
  wire  ram_payload_addr_block_T_1160_addr;
  wire  ram_payload_addr_block_T_1160_mask;
  wire  ram_payload_addr_block_T_1160_en;
  reg [1:0] ram_payload_client_xact_id [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1160_data;
  wire  ram_payload_client_xact_id_T_1160_addr;
  wire  ram_payload_client_xact_id_T_1160_mask;
  wire  ram_payload_client_xact_id_T_1160_en;
  reg [2:0] ram_payload_addr_beat [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1160_data;
  wire  ram_payload_addr_beat_T_1160_addr;
  wire  ram_payload_addr_beat_T_1160_mask;
  wire  ram_payload_addr_beat_T_1160_en;
  reg  ram_payload_is_builtin_type [0:0];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1294_data;
  wire  ram_payload_is_builtin_type_T_1294_addr;
  wire  ram_payload_is_builtin_type_T_1294_en;
  wire  ram_payload_is_builtin_type_T_1160_data;
  wire  ram_payload_is_builtin_type_T_1160_addr;
  wire  ram_payload_is_builtin_type_T_1160_mask;
  wire  ram_payload_is_builtin_type_T_1160_en;
  reg [2:0] ram_payload_a_type [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_a_type_T_1294_data;
  wire  ram_payload_a_type_T_1294_addr;
  wire  ram_payload_a_type_T_1294_en;
  wire [2:0] ram_payload_a_type_T_1160_data;
  wire  ram_payload_a_type_T_1160_addr;
  wire  ram_payload_a_type_T_1160_mask;
  wire  ram_payload_a_type_T_1160_en;
  reg [11:0] ram_payload_union [0:0];
  reg [31:0] GEN_7;
  wire [11:0] ram_payload_union_T_1294_data;
  wire  ram_payload_union_T_1294_addr;
  wire  ram_payload_union_T_1294_en;
  wire [11:0] ram_payload_union_T_1160_data;
  wire  ram_payload_union_T_1160_addr;
  wire  ram_payload_union_T_1160_mask;
  wire  ram_payload_union_T_1160_en;
  reg [63:0] ram_payload_data [0:0];
  reg [63:0] GEN_8;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1160_data;
  wire  ram_payload_data_T_1160_addr;
  wire  ram_payload_data_T_1160_mask;
  wire  ram_payload_data_T_1160_en;
  reg  maybe_full;
  reg [31:0] GEN_9;
  wire  T_1157;
  wire  T_1158;
  wire  do_enq;
  wire  T_1159;
  wire  do_deq;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire [1:0] T_1421;
  wire  ptr_diff;
  wire [1:0] T_1423;
  assign io_enq_ready = T_1157;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1294_data;
  assign io_deq_bits_payload_a_type = ram_payload_a_type_T_1294_data;
  assign io_deq_bits_payload_union = ram_payload_union_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1423[0];
  assign ram_header_src_T_1294_addr = 1'h0;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 1'h1 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1160_data = io_enq_bits_header_src;
  assign ram_header_src_T_1160_addr = 1'h0;
  assign ram_header_src_T_1160_mask = do_enq;
  assign ram_header_src_T_1160_en = do_enq;
  assign ram_header_dst_T_1294_addr = 1'h0;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 1'h1 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1160_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1160_addr = 1'h0;
  assign ram_header_dst_T_1160_mask = do_enq;
  assign ram_header_dst_T_1160_en = do_enq;
  assign ram_payload_addr_block_T_1294_addr = 1'h0;
  assign ram_payload_addr_block_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `else
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block_T_1294_addr >= 1'h1 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `endif
  assign ram_payload_addr_block_T_1160_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1160_addr = 1'h0;
  assign ram_payload_addr_block_T_1160_mask = do_enq;
  assign ram_payload_addr_block_T_1160_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 1'h1 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1160_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1160_addr = 1'h0;
  assign ram_payload_client_xact_id_T_1160_mask = do_enq;
  assign ram_payload_client_xact_id_T_1160_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = 1'h0;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 1'h1 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1160_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1160_addr = 1'h0;
  assign ram_payload_addr_beat_T_1160_mask = do_enq;
  assign ram_payload_addr_beat_T_1160_en = do_enq;
  assign ram_payload_is_builtin_type_T_1294_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `else
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type_T_1294_addr >= 1'h1 ? $random : ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `endif
  assign ram_payload_is_builtin_type_T_1160_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1160_addr = 1'h0;
  assign ram_payload_is_builtin_type_T_1160_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1160_en = do_enq;
  assign ram_payload_a_type_T_1294_addr = 1'h0;
  assign ram_payload_a_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_a_type_T_1294_data = ram_payload_a_type[ram_payload_a_type_T_1294_addr];
  `else
  assign ram_payload_a_type_T_1294_data = ram_payload_a_type_T_1294_addr >= 1'h1 ? $random : ram_payload_a_type[ram_payload_a_type_T_1294_addr];
  `endif
  assign ram_payload_a_type_T_1160_data = io_enq_bits_payload_a_type;
  assign ram_payload_a_type_T_1160_addr = 1'h0;
  assign ram_payload_a_type_T_1160_mask = do_enq;
  assign ram_payload_a_type_T_1160_en = do_enq;
  assign ram_payload_union_T_1294_addr = 1'h0;
  assign ram_payload_union_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_union_T_1294_data = ram_payload_union[ram_payload_union_T_1294_addr];
  `else
  assign ram_payload_union_T_1294_data = ram_payload_union_T_1294_addr >= 1'h1 ? $random : ram_payload_union[ram_payload_union_T_1294_addr];
  `endif
  assign ram_payload_union_T_1160_data = io_enq_bits_payload_union;
  assign ram_payload_union_T_1160_addr = 1'h0;
  assign ram_payload_union_T_1160_mask = do_enq;
  assign ram_payload_union_T_1160_en = do_enq;
  assign ram_payload_data_T_1294_addr = 1'h0;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 1'h1 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1160_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1160_addr = 1'h0;
  assign ram_payload_data_T_1160_mask = do_enq;
  assign ram_payload_data_T_1160_en = do_enq;
  assign T_1157 = maybe_full == 1'h0;
  assign T_1158 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1158;
  assign T_1159 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1159;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = T_1157 == 1'h0;
  assign T_1421 = 1'h0 - 1'h0;
  assign ptr_diff = T_1421[0:0];
  assign T_1423 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[2:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_a_type[initvar] = GEN_6[2:0];
  GEN_7 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_union[initvar] = GEN_7[11:0];
  GEN_8 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_8[63:0];
  GEN_9 = {1{$random}};
  maybe_full = GEN_9[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1160_en & ram_header_src_T_1160_mask) begin
      ram_header_src[ram_header_src_T_1160_addr] <= ram_header_src_T_1160_data;
    end
    if(ram_header_dst_T_1160_en & ram_header_dst_T_1160_mask) begin
      ram_header_dst[ram_header_dst_T_1160_addr] <= ram_header_dst_T_1160_data;
    end
    if(ram_payload_addr_block_T_1160_en & ram_payload_addr_block_T_1160_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1160_addr] <= ram_payload_addr_block_T_1160_data;
    end
    if(ram_payload_client_xact_id_T_1160_en & ram_payload_client_xact_id_T_1160_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1160_addr] <= ram_payload_client_xact_id_T_1160_data;
    end
    if(ram_payload_addr_beat_T_1160_en & ram_payload_addr_beat_T_1160_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1160_addr] <= ram_payload_addr_beat_T_1160_data;
    end
    if(ram_payload_is_builtin_type_T_1160_en & ram_payload_is_builtin_type_T_1160_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1160_addr] <= ram_payload_is_builtin_type_T_1160_data;
    end
    if(ram_payload_a_type_T_1160_en & ram_payload_a_type_T_1160_mask) begin
      ram_payload_a_type[ram_payload_a_type_T_1160_addr] <= ram_payload_a_type_T_1160_data;
    end
    if(ram_payload_union_T_1160_en & ram_payload_union_T_1160_mask) begin
      ram_payload_union[ram_payload_union_T_1160_addr] <= ram_payload_union_T_1160_data;
    end
    if(ram_payload_data_T_1160_en & ram_payload_data_T_1160_mask) begin
      ram_payload_data[ram_payload_data_T_1160_addr] <= ram_payload_data_T_1160_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_21;
    end
  end
endmodule
module Queue_1(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_header_src,
  input  [2:0] io_enq_bits_header_dst,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_p_type,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_header_src,
  output [2:0] io_deq_bits_header_dst,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_p_type,
  output  io_count
);
  reg [2:0] ram_header_src [0:0];
  reg [31:0] GEN_0;
  wire [2:0] ram_header_src_T_1244_data;
  wire  ram_header_src_T_1244_addr;
  wire  ram_header_src_T_1244_en;
  wire [2:0] ram_header_src_T_1115_data;
  wire  ram_header_src_T_1115_addr;
  wire  ram_header_src_T_1115_mask;
  wire  ram_header_src_T_1115_en;
  reg [2:0] ram_header_dst [0:0];
  reg [31:0] GEN_1;
  wire [2:0] ram_header_dst_T_1244_data;
  wire  ram_header_dst_T_1244_addr;
  wire  ram_header_dst_T_1244_en;
  wire [2:0] ram_header_dst_T_1115_data;
  wire  ram_header_dst_T_1115_addr;
  wire  ram_header_dst_T_1115_mask;
  wire  ram_header_dst_T_1115_en;
  reg [25:0] ram_payload_addr_block [0:0];
  reg [31:0] GEN_2;
  wire [25:0] ram_payload_addr_block_T_1244_data;
  wire  ram_payload_addr_block_T_1244_addr;
  wire  ram_payload_addr_block_T_1244_en;
  wire [25:0] ram_payload_addr_block_T_1115_data;
  wire  ram_payload_addr_block_T_1115_addr;
  wire  ram_payload_addr_block_T_1115_mask;
  wire  ram_payload_addr_block_T_1115_en;
  reg [1:0] ram_payload_p_type [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_p_type_T_1244_data;
  wire  ram_payload_p_type_T_1244_addr;
  wire  ram_payload_p_type_T_1244_en;
  wire [1:0] ram_payload_p_type_T_1115_data;
  wire  ram_payload_p_type_T_1115_addr;
  wire  ram_payload_p_type_T_1115_mask;
  wire  ram_payload_p_type_T_1115_en;
  reg  maybe_full;
  reg [31:0] GEN_4;
  wire  T_1112;
  wire  T_1113;
  wire  do_enq;
  wire  T_1114;
  wire  do_deq;
  wire  T_1239;
  wire  GEN_11;
  wire  T_1241;
  wire [1:0] T_1366;
  wire  ptr_diff;
  wire [1:0] T_1368;
  assign io_enq_ready = T_1112;
  assign io_deq_valid = T_1241;
  assign io_deq_bits_header_src = ram_header_src_T_1244_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1244_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1244_data;
  assign io_deq_bits_payload_p_type = ram_payload_p_type_T_1244_data;
  assign io_count = T_1368[0];
  assign ram_header_src_T_1244_addr = 1'h0;
  assign ram_header_src_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1244_data = ram_header_src[ram_header_src_T_1244_addr];
  `else
  assign ram_header_src_T_1244_data = ram_header_src_T_1244_addr >= 1'h1 ? $random : ram_header_src[ram_header_src_T_1244_addr];
  `endif
  assign ram_header_src_T_1115_data = io_enq_bits_header_src;
  assign ram_header_src_T_1115_addr = 1'h0;
  assign ram_header_src_T_1115_mask = do_enq;
  assign ram_header_src_T_1115_en = do_enq;
  assign ram_header_dst_T_1244_addr = 1'h0;
  assign ram_header_dst_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1244_data = ram_header_dst[ram_header_dst_T_1244_addr];
  `else
  assign ram_header_dst_T_1244_data = ram_header_dst_T_1244_addr >= 1'h1 ? $random : ram_header_dst[ram_header_dst_T_1244_addr];
  `endif
  assign ram_header_dst_T_1115_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1115_addr = 1'h0;
  assign ram_header_dst_T_1115_mask = do_enq;
  assign ram_header_dst_T_1115_en = do_enq;
  assign ram_payload_addr_block_T_1244_addr = 1'h0;
  assign ram_payload_addr_block_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1244_data = ram_payload_addr_block[ram_payload_addr_block_T_1244_addr];
  `else
  assign ram_payload_addr_block_T_1244_data = ram_payload_addr_block_T_1244_addr >= 1'h1 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1244_addr];
  `endif
  assign ram_payload_addr_block_T_1115_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1115_addr = 1'h0;
  assign ram_payload_addr_block_T_1115_mask = do_enq;
  assign ram_payload_addr_block_T_1115_en = do_enq;
  assign ram_payload_p_type_T_1244_addr = 1'h0;
  assign ram_payload_p_type_T_1244_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_p_type_T_1244_data = ram_payload_p_type[ram_payload_p_type_T_1244_addr];
  `else
  assign ram_payload_p_type_T_1244_data = ram_payload_p_type_T_1244_addr >= 1'h1 ? $random : ram_payload_p_type[ram_payload_p_type_T_1244_addr];
  `endif
  assign ram_payload_p_type_T_1115_data = io_enq_bits_payload_p_type;
  assign ram_payload_p_type_T_1115_addr = 1'h0;
  assign ram_payload_p_type_T_1115_mask = do_enq;
  assign ram_payload_p_type_T_1115_en = do_enq;
  assign T_1112 = maybe_full == 1'h0;
  assign T_1113 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1113;
  assign T_1114 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1114;
  assign T_1239 = do_enq != do_deq;
  assign GEN_11 = T_1239 ? do_enq : maybe_full;
  assign T_1241 = T_1112 == 1'h0;
  assign T_1366 = 1'h0 - 1'h0;
  assign ptr_diff = T_1366[0:0];
  assign T_1368 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[2:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_2[25:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_payload_p_type[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  maybe_full = GEN_4[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1115_en & ram_header_src_T_1115_mask) begin
      ram_header_src[ram_header_src_T_1115_addr] <= ram_header_src_T_1115_data;
    end
    if(ram_header_dst_T_1115_en & ram_header_dst_T_1115_mask) begin
      ram_header_dst[ram_header_dst_T_1115_addr] <= ram_header_dst_T_1115_data;
    end
    if(ram_payload_addr_block_T_1115_en & ram_payload_addr_block_T_1115_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1115_addr] <= ram_payload_addr_block_T_1115_data;
    end
    if(ram_payload_p_type_T_1115_en & ram_payload_p_type_T_1115_mask) begin
      ram_payload_p_type[ram_payload_p_type_T_1115_addr] <= ram_payload_p_type_T_1115_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_11;
    end
  end
endmodule
module Queue_2(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_header_src,
  input  [2:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [25:0] io_enq_bits_payload_addr_block,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input   io_enq_bits_payload_voluntary,
  input  [2:0] io_enq_bits_payload_r_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_header_src,
  output [2:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [25:0] io_deq_bits_payload_addr_block,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output  io_deq_bits_payload_voluntary,
  output [2:0] io_deq_bits_payload_r_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [2:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [2:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [2:0] ram_header_src_T_1153_data;
  wire  ram_header_src_T_1153_addr;
  wire  ram_header_src_T_1153_mask;
  wire  ram_header_src_T_1153_en;
  reg [2:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [2:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [2:0] ram_header_dst_T_1153_data;
  wire  ram_header_dst_T_1153_addr;
  wire  ram_header_dst_T_1153_mask;
  wire  ram_header_dst_T_1153_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1153_data;
  wire  ram_payload_addr_beat_T_1153_addr;
  wire  ram_payload_addr_beat_T_1153_mask;
  wire  ram_payload_addr_beat_T_1153_en;
  reg [25:0] ram_payload_addr_block [0:1];
  reg [31:0] GEN_3;
  wire [25:0] ram_payload_addr_block_T_1294_data;
  wire  ram_payload_addr_block_T_1294_addr;
  wire  ram_payload_addr_block_T_1294_en;
  wire [25:0] ram_payload_addr_block_T_1153_data;
  wire  ram_payload_addr_block_T_1153_addr;
  wire  ram_payload_addr_block_T_1153_mask;
  wire  ram_payload_addr_block_T_1153_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1153_data;
  wire  ram_payload_client_xact_id_T_1153_addr;
  wire  ram_payload_client_xact_id_T_1153_mask;
  wire  ram_payload_client_xact_id_T_1153_en;
  reg  ram_payload_voluntary [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_voluntary_T_1294_data;
  wire  ram_payload_voluntary_T_1294_addr;
  wire  ram_payload_voluntary_T_1294_en;
  wire  ram_payload_voluntary_T_1153_data;
  wire  ram_payload_voluntary_T_1153_addr;
  wire  ram_payload_voluntary_T_1153_mask;
  wire  ram_payload_voluntary_T_1153_en;
  reg [2:0] ram_payload_r_type [0:1];
  reg [31:0] GEN_6;
  wire [2:0] ram_payload_r_type_T_1294_data;
  wire  ram_payload_r_type_T_1294_addr;
  wire  ram_payload_r_type_T_1294_en;
  wire [2:0] ram_payload_r_type_T_1153_data;
  wire  ram_payload_r_type_T_1153_addr;
  wire  ram_payload_r_type_T_1153_mask;
  wire  ram_payload_r_type_T_1153_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1153_data;
  wire  ram_payload_data_T_1153_addr;
  wire  ram_payload_data_T_1153_mask;
  wire  ram_payload_data_T_1153_en;
  reg  T_1145;
  reg [31:0] GEN_8;
  reg  T_1147;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1150;
  wire  empty;
  wire  full;
  wire  T_1151;
  wire  do_enq;
  wire  T_1152;
  wire  do_deq;
  wire [1:0] T_1282;
  wire  T_1283;
  wire  GEN_19;
  wire [1:0] T_1287;
  wire  T_1288;
  wire  GEN_20;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire  T_1293;
  wire [1:0] T_1420;
  wire  ptr_diff;
  wire  T_1421;
  wire [1:0] T_1422;
  assign io_enq_ready = T_1293;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_addr_block = ram_payload_addr_block_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_voluntary = ram_payload_voluntary_T_1294_data;
  assign io_deq_bits_payload_r_type = ram_payload_r_type_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1422;
  assign ram_header_src_T_1294_addr = T_1147;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 2'h2 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1153_data = io_enq_bits_header_src;
  assign ram_header_src_T_1153_addr = T_1145;
  assign ram_header_src_T_1153_mask = do_enq;
  assign ram_header_src_T_1153_en = do_enq;
  assign ram_header_dst_T_1294_addr = T_1147;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 2'h2 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1153_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1153_addr = T_1145;
  assign ram_header_dst_T_1153_mask = do_enq;
  assign ram_header_dst_T_1153_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = T_1147;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1153_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1153_addr = T_1145;
  assign ram_payload_addr_beat_T_1153_mask = do_enq;
  assign ram_payload_addr_beat_T_1153_en = do_enq;
  assign ram_payload_addr_block_T_1294_addr = T_1147;
  assign ram_payload_addr_block_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `else
  assign ram_payload_addr_block_T_1294_data = ram_payload_addr_block_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_block[ram_payload_addr_block_T_1294_addr];
  `endif
  assign ram_payload_addr_block_T_1153_data = io_enq_bits_payload_addr_block;
  assign ram_payload_addr_block_T_1153_addr = T_1145;
  assign ram_payload_addr_block_T_1153_mask = do_enq;
  assign ram_payload_addr_block_T_1153_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = T_1147;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1153_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1153_addr = T_1145;
  assign ram_payload_client_xact_id_T_1153_mask = do_enq;
  assign ram_payload_client_xact_id_T_1153_en = do_enq;
  assign ram_payload_voluntary_T_1294_addr = T_1147;
  assign ram_payload_voluntary_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_voluntary_T_1294_data = ram_payload_voluntary[ram_payload_voluntary_T_1294_addr];
  `else
  assign ram_payload_voluntary_T_1294_data = ram_payload_voluntary_T_1294_addr >= 2'h2 ? $random : ram_payload_voluntary[ram_payload_voluntary_T_1294_addr];
  `endif
  assign ram_payload_voluntary_T_1153_data = io_enq_bits_payload_voluntary;
  assign ram_payload_voluntary_T_1153_addr = T_1145;
  assign ram_payload_voluntary_T_1153_mask = do_enq;
  assign ram_payload_voluntary_T_1153_en = do_enq;
  assign ram_payload_r_type_T_1294_addr = T_1147;
  assign ram_payload_r_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_r_type_T_1294_data = ram_payload_r_type[ram_payload_r_type_T_1294_addr];
  `else
  assign ram_payload_r_type_T_1294_data = ram_payload_r_type_T_1294_addr >= 2'h2 ? $random : ram_payload_r_type[ram_payload_r_type_T_1294_addr];
  `endif
  assign ram_payload_r_type_T_1153_data = io_enq_bits_payload_r_type;
  assign ram_payload_r_type_T_1153_addr = T_1145;
  assign ram_payload_r_type_T_1153_mask = do_enq;
  assign ram_payload_r_type_T_1153_en = do_enq;
  assign ram_payload_data_T_1294_addr = T_1147;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 2'h2 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1153_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1153_addr = T_1145;
  assign ram_payload_data_T_1153_mask = do_enq;
  assign ram_payload_data_T_1153_en = do_enq;
  assign ptr_match = T_1145 == T_1147;
  assign T_1150 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1150;
  assign full = ptr_match & maybe_full;
  assign T_1151 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1151;
  assign T_1152 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1152;
  assign T_1282 = T_1145 + 1'h1;
  assign T_1283 = T_1282[0:0];
  assign GEN_19 = do_enq ? T_1283 : T_1145;
  assign T_1287 = T_1147 + 1'h1;
  assign T_1288 = T_1287[0:0];
  assign GEN_20 = do_deq ? T_1288 : T_1147;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = empty == 1'h0;
  assign T_1293 = full == 1'h0;
  assign T_1420 = T_1145 - T_1147;
  assign ptr_diff = T_1420[0:0];
  assign T_1421 = maybe_full & ptr_match;
  assign T_1422 = {T_1421,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[2:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_block[initvar] = GEN_3[25:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_4[1:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_voluntary[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_r_type[initvar] = GEN_6[2:0];
  GEN_7 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  GEN_8 = {1{$random}};
  T_1145 = GEN_8[0:0];
  GEN_9 = {1{$random}};
  T_1147 = GEN_9[0:0];
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1153_en & ram_header_src_T_1153_mask) begin
      ram_header_src[ram_header_src_T_1153_addr] <= ram_header_src_T_1153_data;
    end
    if(ram_header_dst_T_1153_en & ram_header_dst_T_1153_mask) begin
      ram_header_dst[ram_header_dst_T_1153_addr] <= ram_header_dst_T_1153_data;
    end
    if(ram_payload_addr_beat_T_1153_en & ram_payload_addr_beat_T_1153_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1153_addr] <= ram_payload_addr_beat_T_1153_data;
    end
    if(ram_payload_addr_block_T_1153_en & ram_payload_addr_block_T_1153_mask) begin
      ram_payload_addr_block[ram_payload_addr_block_T_1153_addr] <= ram_payload_addr_block_T_1153_data;
    end
    if(ram_payload_client_xact_id_T_1153_en & ram_payload_client_xact_id_T_1153_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1153_addr] <= ram_payload_client_xact_id_T_1153_data;
    end
    if(ram_payload_voluntary_T_1153_en & ram_payload_voluntary_T_1153_mask) begin
      ram_payload_voluntary[ram_payload_voluntary_T_1153_addr] <= ram_payload_voluntary_T_1153_data;
    end
    if(ram_payload_r_type_T_1153_en & ram_payload_r_type_T_1153_mask) begin
      ram_payload_r_type[ram_payload_r_type_T_1153_addr] <= ram_payload_r_type_T_1153_data;
    end
    if(ram_payload_data_T_1153_en & ram_payload_data_T_1153_mask) begin
      ram_payload_data[ram_payload_data_T_1153_addr] <= ram_payload_data_T_1153_data;
    end
    if(reset) begin
      T_1145 <= 1'h0;
    end else begin
      T_1145 <= GEN_19;
    end
    if(reset) begin
      T_1147 <= 1'h0;
    end else begin
      T_1147 <= GEN_20;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_21;
    end
  end
endmodule
module Queue_3(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_header_src,
  input  [2:0] io_enq_bits_header_dst,
  input  [2:0] io_enq_bits_payload_addr_beat,
  input  [1:0] io_enq_bits_payload_client_xact_id,
  input  [2:0] io_enq_bits_payload_manager_xact_id,
  input   io_enq_bits_payload_is_builtin_type,
  input  [3:0] io_enq_bits_payload_g_type,
  input  [63:0] io_enq_bits_payload_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_header_src,
  output [2:0] io_deq_bits_header_dst,
  output [2:0] io_deq_bits_payload_addr_beat,
  output [1:0] io_deq_bits_payload_client_xact_id,
  output [2:0] io_deq_bits_payload_manager_xact_id,
  output  io_deq_bits_payload_is_builtin_type,
  output [3:0] io_deq_bits_payload_g_type,
  output [63:0] io_deq_bits_payload_data,
  output [1:0] io_count
);
  reg [2:0] ram_header_src [0:1];
  reg [31:0] GEN_0;
  wire [2:0] ram_header_src_T_1294_data;
  wire  ram_header_src_T_1294_addr;
  wire  ram_header_src_T_1294_en;
  wire [2:0] ram_header_src_T_1153_data;
  wire  ram_header_src_T_1153_addr;
  wire  ram_header_src_T_1153_mask;
  wire  ram_header_src_T_1153_en;
  reg [2:0] ram_header_dst [0:1];
  reg [31:0] GEN_1;
  wire [2:0] ram_header_dst_T_1294_data;
  wire  ram_header_dst_T_1294_addr;
  wire  ram_header_dst_T_1294_en;
  wire [2:0] ram_header_dst_T_1153_data;
  wire  ram_header_dst_T_1153_addr;
  wire  ram_header_dst_T_1153_mask;
  wire  ram_header_dst_T_1153_en;
  reg [2:0] ram_payload_addr_beat [0:1];
  reg [31:0] GEN_2;
  wire [2:0] ram_payload_addr_beat_T_1294_data;
  wire  ram_payload_addr_beat_T_1294_addr;
  wire  ram_payload_addr_beat_T_1294_en;
  wire [2:0] ram_payload_addr_beat_T_1153_data;
  wire  ram_payload_addr_beat_T_1153_addr;
  wire  ram_payload_addr_beat_T_1153_mask;
  wire  ram_payload_addr_beat_T_1153_en;
  reg [1:0] ram_payload_client_xact_id [0:1];
  reg [31:0] GEN_3;
  wire [1:0] ram_payload_client_xact_id_T_1294_data;
  wire  ram_payload_client_xact_id_T_1294_addr;
  wire  ram_payload_client_xact_id_T_1294_en;
  wire [1:0] ram_payload_client_xact_id_T_1153_data;
  wire  ram_payload_client_xact_id_T_1153_addr;
  wire  ram_payload_client_xact_id_T_1153_mask;
  wire  ram_payload_client_xact_id_T_1153_en;
  reg [2:0] ram_payload_manager_xact_id [0:1];
  reg [31:0] GEN_4;
  wire [2:0] ram_payload_manager_xact_id_T_1294_data;
  wire  ram_payload_manager_xact_id_T_1294_addr;
  wire  ram_payload_manager_xact_id_T_1294_en;
  wire [2:0] ram_payload_manager_xact_id_T_1153_data;
  wire  ram_payload_manager_xact_id_T_1153_addr;
  wire  ram_payload_manager_xact_id_T_1153_mask;
  wire  ram_payload_manager_xact_id_T_1153_en;
  reg  ram_payload_is_builtin_type [0:1];
  reg [31:0] GEN_5;
  wire  ram_payload_is_builtin_type_T_1294_data;
  wire  ram_payload_is_builtin_type_T_1294_addr;
  wire  ram_payload_is_builtin_type_T_1294_en;
  wire  ram_payload_is_builtin_type_T_1153_data;
  wire  ram_payload_is_builtin_type_T_1153_addr;
  wire  ram_payload_is_builtin_type_T_1153_mask;
  wire  ram_payload_is_builtin_type_T_1153_en;
  reg [3:0] ram_payload_g_type [0:1];
  reg [31:0] GEN_6;
  wire [3:0] ram_payload_g_type_T_1294_data;
  wire  ram_payload_g_type_T_1294_addr;
  wire  ram_payload_g_type_T_1294_en;
  wire [3:0] ram_payload_g_type_T_1153_data;
  wire  ram_payload_g_type_T_1153_addr;
  wire  ram_payload_g_type_T_1153_mask;
  wire  ram_payload_g_type_T_1153_en;
  reg [63:0] ram_payload_data [0:1];
  reg [63:0] GEN_7;
  wire [63:0] ram_payload_data_T_1294_data;
  wire  ram_payload_data_T_1294_addr;
  wire  ram_payload_data_T_1294_en;
  wire [63:0] ram_payload_data_T_1153_data;
  wire  ram_payload_data_T_1153_addr;
  wire  ram_payload_data_T_1153_mask;
  wire  ram_payload_data_T_1153_en;
  reg  T_1145;
  reg [31:0] GEN_8;
  reg  T_1147;
  reg [31:0] GEN_9;
  reg  maybe_full;
  reg [31:0] GEN_10;
  wire  ptr_match;
  wire  T_1150;
  wire  empty;
  wire  full;
  wire  T_1151;
  wire  do_enq;
  wire  T_1152;
  wire  do_deq;
  wire [1:0] T_1282;
  wire  T_1283;
  wire  GEN_19;
  wire [1:0] T_1287;
  wire  T_1288;
  wire  GEN_20;
  wire  T_1289;
  wire  GEN_21;
  wire  T_1291;
  wire  T_1293;
  wire [1:0] T_1420;
  wire  ptr_diff;
  wire  T_1421;
  wire [1:0] T_1422;
  assign io_enq_ready = T_1293;
  assign io_deq_valid = T_1291;
  assign io_deq_bits_header_src = ram_header_src_T_1294_data;
  assign io_deq_bits_header_dst = ram_header_dst_T_1294_data;
  assign io_deq_bits_payload_addr_beat = ram_payload_addr_beat_T_1294_data;
  assign io_deq_bits_payload_client_xact_id = ram_payload_client_xact_id_T_1294_data;
  assign io_deq_bits_payload_manager_xact_id = ram_payload_manager_xact_id_T_1294_data;
  assign io_deq_bits_payload_is_builtin_type = ram_payload_is_builtin_type_T_1294_data;
  assign io_deq_bits_payload_g_type = ram_payload_g_type_T_1294_data;
  assign io_deq_bits_payload_data = ram_payload_data_T_1294_data;
  assign io_count = T_1422;
  assign ram_header_src_T_1294_addr = T_1147;
  assign ram_header_src_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_src_T_1294_data = ram_header_src[ram_header_src_T_1294_addr];
  `else
  assign ram_header_src_T_1294_data = ram_header_src_T_1294_addr >= 2'h2 ? $random : ram_header_src[ram_header_src_T_1294_addr];
  `endif
  assign ram_header_src_T_1153_data = io_enq_bits_header_src;
  assign ram_header_src_T_1153_addr = T_1145;
  assign ram_header_src_T_1153_mask = do_enq;
  assign ram_header_src_T_1153_en = do_enq;
  assign ram_header_dst_T_1294_addr = T_1147;
  assign ram_header_dst_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_header_dst_T_1294_data = ram_header_dst[ram_header_dst_T_1294_addr];
  `else
  assign ram_header_dst_T_1294_data = ram_header_dst_T_1294_addr >= 2'h2 ? $random : ram_header_dst[ram_header_dst_T_1294_addr];
  `endif
  assign ram_header_dst_T_1153_data = io_enq_bits_header_dst;
  assign ram_header_dst_T_1153_addr = T_1145;
  assign ram_header_dst_T_1153_mask = do_enq;
  assign ram_header_dst_T_1153_en = do_enq;
  assign ram_payload_addr_beat_T_1294_addr = T_1147;
  assign ram_payload_addr_beat_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `else
  assign ram_payload_addr_beat_T_1294_data = ram_payload_addr_beat_T_1294_addr >= 2'h2 ? $random : ram_payload_addr_beat[ram_payload_addr_beat_T_1294_addr];
  `endif
  assign ram_payload_addr_beat_T_1153_data = io_enq_bits_payload_addr_beat;
  assign ram_payload_addr_beat_T_1153_addr = T_1145;
  assign ram_payload_addr_beat_T_1153_mask = do_enq;
  assign ram_payload_addr_beat_T_1153_en = do_enq;
  assign ram_payload_client_xact_id_T_1294_addr = T_1147;
  assign ram_payload_client_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `else
  assign ram_payload_client_xact_id_T_1294_data = ram_payload_client_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_client_xact_id[ram_payload_client_xact_id_T_1294_addr];
  `endif
  assign ram_payload_client_xact_id_T_1153_data = io_enq_bits_payload_client_xact_id;
  assign ram_payload_client_xact_id_T_1153_addr = T_1145;
  assign ram_payload_client_xact_id_T_1153_mask = do_enq;
  assign ram_payload_client_xact_id_T_1153_en = do_enq;
  assign ram_payload_manager_xact_id_T_1294_addr = T_1147;
  assign ram_payload_manager_xact_id_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_manager_xact_id_T_1294_data = ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1294_addr];
  `else
  assign ram_payload_manager_xact_id_T_1294_data = ram_payload_manager_xact_id_T_1294_addr >= 2'h2 ? $random : ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1294_addr];
  `endif
  assign ram_payload_manager_xact_id_T_1153_data = io_enq_bits_payload_manager_xact_id;
  assign ram_payload_manager_xact_id_T_1153_addr = T_1145;
  assign ram_payload_manager_xact_id_T_1153_mask = do_enq;
  assign ram_payload_manager_xact_id_T_1153_en = do_enq;
  assign ram_payload_is_builtin_type_T_1294_addr = T_1147;
  assign ram_payload_is_builtin_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `else
  assign ram_payload_is_builtin_type_T_1294_data = ram_payload_is_builtin_type_T_1294_addr >= 2'h2 ? $random : ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1294_addr];
  `endif
  assign ram_payload_is_builtin_type_T_1153_data = io_enq_bits_payload_is_builtin_type;
  assign ram_payload_is_builtin_type_T_1153_addr = T_1145;
  assign ram_payload_is_builtin_type_T_1153_mask = do_enq;
  assign ram_payload_is_builtin_type_T_1153_en = do_enq;
  assign ram_payload_g_type_T_1294_addr = T_1147;
  assign ram_payload_g_type_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_g_type_T_1294_data = ram_payload_g_type[ram_payload_g_type_T_1294_addr];
  `else
  assign ram_payload_g_type_T_1294_data = ram_payload_g_type_T_1294_addr >= 2'h2 ? $random : ram_payload_g_type[ram_payload_g_type_T_1294_addr];
  `endif
  assign ram_payload_g_type_T_1153_data = io_enq_bits_payload_g_type;
  assign ram_payload_g_type_T_1153_addr = T_1145;
  assign ram_payload_g_type_T_1153_mask = do_enq;
  assign ram_payload_g_type_T_1153_en = do_enq;
  assign ram_payload_data_T_1294_addr = T_1147;
  assign ram_payload_data_T_1294_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_payload_data_T_1294_data = ram_payload_data[ram_payload_data_T_1294_addr];
  `else
  assign ram_payload_data_T_1294_data = ram_payload_data_T_1294_addr >= 2'h2 ? $random : ram_payload_data[ram_payload_data_T_1294_addr];
  `endif
  assign ram_payload_data_T_1153_data = io_enq_bits_payload_data;
  assign ram_payload_data_T_1153_addr = T_1145;
  assign ram_payload_data_T_1153_mask = do_enq;
  assign ram_payload_data_T_1153_en = do_enq;
  assign ptr_match = T_1145 == T_1147;
  assign T_1150 = maybe_full == 1'h0;
  assign empty = ptr_match & T_1150;
  assign full = ptr_match & maybe_full;
  assign T_1151 = io_enq_ready & io_enq_valid;
  assign do_enq = T_1151;
  assign T_1152 = io_deq_ready & io_deq_valid;
  assign do_deq = T_1152;
  assign T_1282 = T_1145 + 1'h1;
  assign T_1283 = T_1282[0:0];
  assign GEN_19 = do_enq ? T_1283 : T_1145;
  assign T_1287 = T_1147 + 1'h1;
  assign T_1288 = T_1287[0:0];
  assign GEN_20 = do_deq ? T_1288 : T_1147;
  assign T_1289 = do_enq != do_deq;
  assign GEN_21 = T_1289 ? do_enq : maybe_full;
  assign T_1291 = empty == 1'h0;
  assign T_1293 = full == 1'h0;
  assign T_1420 = T_1145 - T_1147;
  assign ptr_diff = T_1420[0:0];
  assign T_1421 = maybe_full & ptr_match;
  assign T_1422 = {T_1421,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_src[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_header_dst[initvar] = GEN_1[2:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_client_xact_id[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_manager_xact_id[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_is_builtin_type[initvar] = GEN_5[0:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_g_type[initvar] = GEN_6[3:0];
  GEN_7 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_payload_data[initvar] = GEN_7[63:0];
  GEN_8 = {1{$random}};
  T_1145 = GEN_8[0:0];
  GEN_9 = {1{$random}};
  T_1147 = GEN_9[0:0];
  GEN_10 = {1{$random}};
  maybe_full = GEN_10[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_header_src_T_1153_en & ram_header_src_T_1153_mask) begin
      ram_header_src[ram_header_src_T_1153_addr] <= ram_header_src_T_1153_data;
    end
    if(ram_header_dst_T_1153_en & ram_header_dst_T_1153_mask) begin
      ram_header_dst[ram_header_dst_T_1153_addr] <= ram_header_dst_T_1153_data;
    end
    if(ram_payload_addr_beat_T_1153_en & ram_payload_addr_beat_T_1153_mask) begin
      ram_payload_addr_beat[ram_payload_addr_beat_T_1153_addr] <= ram_payload_addr_beat_T_1153_data;
    end
    if(ram_payload_client_xact_id_T_1153_en & ram_payload_client_xact_id_T_1153_mask) begin
      ram_payload_client_xact_id[ram_payload_client_xact_id_T_1153_addr] <= ram_payload_client_xact_id_T_1153_data;
    end
    if(ram_payload_manager_xact_id_T_1153_en & ram_payload_manager_xact_id_T_1153_mask) begin
      ram_payload_manager_xact_id[ram_payload_manager_xact_id_T_1153_addr] <= ram_payload_manager_xact_id_T_1153_data;
    end
    if(ram_payload_is_builtin_type_T_1153_en & ram_payload_is_builtin_type_T_1153_mask) begin
      ram_payload_is_builtin_type[ram_payload_is_builtin_type_T_1153_addr] <= ram_payload_is_builtin_type_T_1153_data;
    end
    if(ram_payload_g_type_T_1153_en & ram_payload_g_type_T_1153_mask) begin
      ram_payload_g_type[ram_payload_g_type_T_1153_addr] <= ram_payload_g_type_T_1153_data;
    end
    if(ram_payload_data_T_1153_en & ram_payload_data_T_1153_mask) begin
      ram_payload_data[ram_payload_data_T_1153_addr] <= ram_payload_data_T_1153_data;
    end
    if(reset) begin
      T_1145 <= 1'h0;
    end else begin
      T_1145 <= GEN_19;
    end
    if(reset) begin
      T_1147 <= 1'h0;
    end else begin
      T_1147 <= GEN_20;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_21;
    end
  end
endmodule
module TileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [2:0] io_client_acquire_bits_header_src,
  input  [2:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_header_src,
  output [2:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_header_src,
  input  [2:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [2:0] io_client_probe_bits_header_src,
  output [2:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_header_src,
  input  [2:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [2:0] io_manager_acquire_bits_header_src,
  output [2:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_header_src,
  input  [2:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_header_src,
  output [2:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [2:0] io_manager_probe_bits_header_src,
  input  [2:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_header_src,
  output [2:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_7774_clk;
  wire  Queue_7774_reset;
  wire  Queue_7774_io_enq_ready;
  wire  Queue_7774_io_enq_valid;
  wire [2:0] Queue_7774_io_enq_bits_header_src;
  wire [2:0] Queue_7774_io_enq_bits_header_dst;
  wire [25:0] Queue_7774_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_7774_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_7774_io_enq_bits_payload_addr_beat;
  wire  Queue_7774_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_7774_io_enq_bits_payload_a_type;
  wire [11:0] Queue_7774_io_enq_bits_payload_union;
  wire [63:0] Queue_7774_io_enq_bits_payload_data;
  wire  Queue_7774_io_deq_ready;
  wire  Queue_7774_io_deq_valid;
  wire [2:0] Queue_7774_io_deq_bits_header_src;
  wire [2:0] Queue_7774_io_deq_bits_header_dst;
  wire [25:0] Queue_7774_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_7774_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_7774_io_deq_bits_payload_addr_beat;
  wire  Queue_7774_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_7774_io_deq_bits_payload_a_type;
  wire [11:0] Queue_7774_io_deq_bits_payload_union;
  wire [63:0] Queue_7774_io_deq_bits_payload_data;
  wire  Queue_7774_io_count;
  wire  Queue_1_7897_clk;
  wire  Queue_1_7897_reset;
  wire  Queue_1_7897_io_enq_ready;
  wire  Queue_1_7897_io_enq_valid;
  wire [2:0] Queue_1_7897_io_enq_bits_header_src;
  wire [2:0] Queue_1_7897_io_enq_bits_header_dst;
  wire [25:0] Queue_1_7897_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_1_7897_io_enq_bits_payload_p_type;
  wire  Queue_1_7897_io_deq_ready;
  wire  Queue_1_7897_io_deq_valid;
  wire [2:0] Queue_1_7897_io_deq_bits_header_src;
  wire [2:0] Queue_1_7897_io_deq_bits_header_dst;
  wire [25:0] Queue_1_7897_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_1_7897_io_deq_bits_payload_p_type;
  wire  Queue_1_7897_io_count;
  wire  Queue_2_8024_clk;
  wire  Queue_2_8024_reset;
  wire  Queue_2_8024_io_enq_ready;
  wire  Queue_2_8024_io_enq_valid;
  wire [2:0] Queue_2_8024_io_enq_bits_header_src;
  wire [2:0] Queue_2_8024_io_enq_bits_header_dst;
  wire [2:0] Queue_2_8024_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_2_8024_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_2_8024_io_enq_bits_payload_client_xact_id;
  wire  Queue_2_8024_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_2_8024_io_enq_bits_payload_r_type;
  wire [63:0] Queue_2_8024_io_enq_bits_payload_data;
  wire  Queue_2_8024_io_deq_ready;
  wire  Queue_2_8024_io_deq_valid;
  wire [2:0] Queue_2_8024_io_deq_bits_header_src;
  wire [2:0] Queue_2_8024_io_deq_bits_header_dst;
  wire [2:0] Queue_2_8024_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_2_8024_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_2_8024_io_deq_bits_payload_client_xact_id;
  wire  Queue_2_8024_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_2_8024_io_deq_bits_payload_r_type;
  wire [63:0] Queue_2_8024_io_deq_bits_payload_data;
  wire [1:0] Queue_2_8024_io_count;
  wire  Queue_3_8151_clk;
  wire  Queue_3_8151_reset;
  wire  Queue_3_8151_io_enq_ready;
  wire  Queue_3_8151_io_enq_valid;
  wire [2:0] Queue_3_8151_io_enq_bits_header_src;
  wire [2:0] Queue_3_8151_io_enq_bits_header_dst;
  wire [2:0] Queue_3_8151_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_3_8151_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_3_8151_io_enq_bits_payload_manager_xact_id;
  wire  Queue_3_8151_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_8151_io_enq_bits_payload_g_type;
  wire [63:0] Queue_3_8151_io_enq_bits_payload_data;
  wire  Queue_3_8151_io_deq_ready;
  wire  Queue_3_8151_io_deq_valid;
  wire [2:0] Queue_3_8151_io_deq_bits_header_src;
  wire [2:0] Queue_3_8151_io_deq_bits_header_dst;
  wire [2:0] Queue_3_8151_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_3_8151_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_3_8151_io_deq_bits_payload_manager_xact_id;
  wire  Queue_3_8151_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_3_8151_io_deq_bits_payload_g_type;
  wire [63:0] Queue_3_8151_io_deq_bits_payload_data;
  wire [1:0] Queue_3_8151_io_count;
  Queue Queue_7774 (
    .clk(Queue_7774_clk),
    .reset(Queue_7774_reset),
    .io_enq_ready(Queue_7774_io_enq_ready),
    .io_enq_valid(Queue_7774_io_enq_valid),
    .io_enq_bits_header_src(Queue_7774_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7774_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_7774_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_7774_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_7774_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_7774_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_7774_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_7774_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_7774_io_enq_bits_payload_data),
    .io_deq_ready(Queue_7774_io_deq_ready),
    .io_deq_valid(Queue_7774_io_deq_valid),
    .io_deq_bits_header_src(Queue_7774_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7774_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_7774_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_7774_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_7774_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_7774_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_7774_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_7774_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_7774_io_deq_bits_payload_data),
    .io_count(Queue_7774_io_count)
  );
  Queue_1 Queue_1_7897 (
    .clk(Queue_1_7897_clk),
    .reset(Queue_1_7897_reset),
    .io_enq_ready(Queue_1_7897_io_enq_ready),
    .io_enq_valid(Queue_1_7897_io_enq_valid),
    .io_enq_bits_header_src(Queue_1_7897_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_1_7897_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_1_7897_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_1_7897_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_1_7897_io_deq_ready),
    .io_deq_valid(Queue_1_7897_io_deq_valid),
    .io_deq_bits_header_src(Queue_1_7897_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_1_7897_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_1_7897_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_1_7897_io_deq_bits_payload_p_type),
    .io_count(Queue_1_7897_io_count)
  );
  Queue_2 Queue_2_8024 (
    .clk(Queue_2_8024_clk),
    .reset(Queue_2_8024_reset),
    .io_enq_ready(Queue_2_8024_io_enq_ready),
    .io_enq_valid(Queue_2_8024_io_enq_valid),
    .io_enq_bits_header_src(Queue_2_8024_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_2_8024_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_2_8024_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_2_8024_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_2_8024_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_2_8024_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_2_8024_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_2_8024_io_enq_bits_payload_data),
    .io_deq_ready(Queue_2_8024_io_deq_ready),
    .io_deq_valid(Queue_2_8024_io_deq_valid),
    .io_deq_bits_header_src(Queue_2_8024_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_2_8024_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_2_8024_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_2_8024_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_2_8024_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_2_8024_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_2_8024_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_2_8024_io_deq_bits_payload_data),
    .io_count(Queue_2_8024_io_count)
  );
  Queue_3 Queue_3_8151 (
    .clk(Queue_3_8151_clk),
    .reset(Queue_3_8151_reset),
    .io_enq_ready(Queue_3_8151_io_enq_ready),
    .io_enq_valid(Queue_3_8151_io_enq_valid),
    .io_enq_bits_header_src(Queue_3_8151_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_3_8151_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_3_8151_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_3_8151_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_3_8151_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_3_8151_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_3_8151_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_3_8151_io_enq_bits_payload_data),
    .io_deq_ready(Queue_3_8151_io_deq_ready),
    .io_deq_valid(Queue_3_8151_io_deq_valid),
    .io_deq_bits_header_src(Queue_3_8151_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_3_8151_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_3_8151_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_3_8151_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_3_8151_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_3_8151_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_3_8151_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_3_8151_io_deq_bits_payload_data),
    .io_count(Queue_3_8151_io_count)
  );
  assign io_client_acquire_ready = Queue_7774_io_enq_ready;
  assign io_client_grant_valid = Queue_3_8151_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_3_8151_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_3_8151_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_3_8151_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_3_8151_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_3_8151_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_3_8151_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_3_8151_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_3_8151_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_1_7897_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_1_7897_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_1_7897_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_1_7897_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_1_7897_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_2_8024_io_enq_ready;
  assign io_manager_acquire_valid = Queue_7774_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_7774_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_7774_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_7774_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_7774_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_7774_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_7774_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_7774_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_7774_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_7774_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_3_8151_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_1_7897_io_enq_ready;
  assign io_manager_release_valid = Queue_2_8024_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_2_8024_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_2_8024_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_2_8024_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_2_8024_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_2_8024_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_2_8024_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_2_8024_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_2_8024_io_deq_bits_payload_data;
  assign Queue_7774_clk = clk;
  assign Queue_7774_reset = reset;
  assign Queue_7774_io_enq_valid = io_client_acquire_valid;
  assign Queue_7774_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_7774_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_7774_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_7774_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_7774_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_7774_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_7774_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_7774_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_7774_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_7774_io_deq_ready = io_manager_acquire_ready;
  assign Queue_1_7897_clk = clk;
  assign Queue_1_7897_reset = reset;
  assign Queue_1_7897_io_enq_valid = io_manager_probe_valid;
  assign Queue_1_7897_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_1_7897_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_1_7897_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_1_7897_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_1_7897_io_deq_ready = io_client_probe_ready;
  assign Queue_2_8024_clk = clk;
  assign Queue_2_8024_reset = reset;
  assign Queue_2_8024_io_enq_valid = io_client_release_valid;
  assign Queue_2_8024_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_2_8024_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_2_8024_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_2_8024_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_2_8024_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_2_8024_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_2_8024_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_2_8024_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_2_8024_io_deq_ready = io_manager_release_ready;
  assign Queue_3_8151_clk = clk;
  assign Queue_3_8151_reset = reset;
  assign Queue_3_8151_io_enq_valid = io_manager_grant_valid;
  assign Queue_3_8151_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_3_8151_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_3_8151_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_3_8151_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_3_8151_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_3_8151_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_3_8151_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_3_8151_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_3_8151_io_deq_ready = io_client_grant_ready;
endmodule
module ClientTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [25:0] io_client_probe_bits_addr_block,
  output [1:0] io_client_probe_bits_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_addr_beat,
  input  [25:0] io_client_release_bits_addr_block,
  input  [1:0] io_client_release_bits_client_xact_id,
  input   io_client_release_bits_voluntary,
  input  [2:0] io_client_release_bits_r_type,
  input  [63:0] io_client_release_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  output  io_client_grant_bits_manager_id,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_manager_xact_id,
  input   io_client_finish_bits_manager_id,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [2:0] io_network_acquire_bits_header_src,
  output [2:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [2:0] io_network_grant_bits_header_src,
  input  [2:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [2:0] io_network_finish_bits_header_src,
  output [2:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [2:0] io_network_probe_bits_header_src,
  input  [2:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [2:0] io_network_release_bits_header_src,
  output [2:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [2:0] acq_with_header_bits_header_src;
  wire [2:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_4395;
  wire  T_4397;
  wire  T_4403;
  wire  rel_with_header_ready;
  wire  rel_with_header_valid;
  wire [2:0] rel_with_header_bits_header_src;
  wire [2:0] rel_with_header_bits_header_dst;
  wire [2:0] rel_with_header_bits_payload_addr_beat;
  wire [25:0] rel_with_header_bits_payload_addr_block;
  wire [1:0] rel_with_header_bits_payload_client_xact_id;
  wire  rel_with_header_bits_payload_voluntary;
  wire [2:0] rel_with_header_bits_payload_r_type;
  wire [63:0] rel_with_header_bits_payload_data;
  wire [31:0] GEN_1;
  wire [31:0] T_5040;
  wire  T_5042;
  wire  T_5048;
  wire  fin_with_header_ready;
  wire  fin_with_header_valid;
  wire [2:0] fin_with_header_bits_header_src;
  wire [2:0] fin_with_header_bits_header_dst;
  wire [2:0] fin_with_header_bits_payload_manager_xact_id;
  wire  fin_with_header_bits_payload_manager_id;
  wire  prb_without_header_ready;
  wire  prb_without_header_valid;
  wire [25:0] prb_without_header_bits_addr_block;
  wire [1:0] prb_without_header_bits_p_type;
  wire  gnt_without_header_ready;
  wire  gnt_without_header_valid;
  wire [2:0] gnt_without_header_bits_addr_beat;
  wire [1:0] gnt_without_header_bits_client_xact_id;
  wire [2:0] gnt_without_header_bits_manager_xact_id;
  wire  gnt_without_header_bits_is_builtin_type;
  wire [3:0] gnt_without_header_bits_g_type;
  wire [63:0] gnt_without_header_bits_data;
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_probe_valid = prb_without_header_valid;
  assign io_client_probe_bits_addr_block = prb_without_header_bits_addr_block;
  assign io_client_probe_bits_p_type = prb_without_header_bits_p_type;
  assign io_client_release_ready = rel_with_header_ready;
  assign io_client_grant_valid = gnt_without_header_valid;
  assign io_client_grant_bits_addr_beat = gnt_without_header_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = gnt_without_header_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = gnt_without_header_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = gnt_without_header_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = gnt_without_header_bits_g_type;
  assign io_client_grant_bits_data = gnt_without_header_bits_data;
  assign io_client_grant_bits_manager_id = io_network_grant_bits_header_src[0];
  assign io_client_finish_ready = fin_with_header_ready;
  assign io_network_acquire_valid = acq_with_header_valid;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = gnt_without_header_ready;
  assign io_network_finish_valid = fin_with_header_valid;
  assign io_network_finish_bits_header_src = fin_with_header_bits_header_src;
  assign io_network_finish_bits_header_dst = fin_with_header_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = fin_with_header_bits_payload_manager_xact_id;
  assign io_network_probe_ready = prb_without_header_ready;
  assign io_network_release_valid = rel_with_header_valid;
  assign io_network_release_bits_header_src = rel_with_header_bits_header_src;
  assign io_network_release_bits_header_dst = rel_with_header_bits_header_dst;
  assign io_network_release_bits_payload_addr_beat = rel_with_header_bits_payload_addr_beat;
  assign io_network_release_bits_payload_addr_block = rel_with_header_bits_payload_addr_block;
  assign io_network_release_bits_payload_client_xact_id = rel_with_header_bits_payload_client_xact_id;
  assign io_network_release_bits_payload_voluntary = rel_with_header_bits_payload_voluntary;
  assign io_network_release_bits_payload_r_type = rel_with_header_bits_payload_r_type;
  assign io_network_release_bits_payload_data = rel_with_header_bits_payload_data;
  assign acq_with_header_ready = io_network_acquire_ready;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = {{2'd0}, 1'h0};
  assign acq_with_header_bits_header_dst = {{2'd0}, T_4403};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_4395 = GEN_0 << 6;
  assign T_4397 = 32'h80000000 <= T_4395;
  assign T_4403 = T_4397 ? 1'h0 : 1'h1;
  assign rel_with_header_ready = io_network_release_ready;
  assign rel_with_header_valid = io_client_release_valid;
  assign rel_with_header_bits_header_src = {{2'd0}, 1'h0};
  assign rel_with_header_bits_header_dst = {{2'd0}, T_5048};
  assign rel_with_header_bits_payload_addr_beat = io_client_release_bits_addr_beat;
  assign rel_with_header_bits_payload_addr_block = io_client_release_bits_addr_block;
  assign rel_with_header_bits_payload_client_xact_id = io_client_release_bits_client_xact_id;
  assign rel_with_header_bits_payload_voluntary = io_client_release_bits_voluntary;
  assign rel_with_header_bits_payload_r_type = io_client_release_bits_r_type;
  assign rel_with_header_bits_payload_data = io_client_release_bits_data;
  assign GEN_1 = {{6'd0}, io_client_release_bits_addr_block};
  assign T_5040 = GEN_1 << 6;
  assign T_5042 = 32'h80000000 <= T_5040;
  assign T_5048 = T_5042 ? 1'h0 : 1'h1;
  assign fin_with_header_ready = io_network_finish_ready;
  assign fin_with_header_valid = io_client_finish_valid;
  assign fin_with_header_bits_header_src = {{2'd0}, 1'h0};
  assign fin_with_header_bits_header_dst = {{2'd0}, io_client_finish_bits_manager_id};
  assign fin_with_header_bits_payload_manager_xact_id = io_client_finish_bits_manager_xact_id;
  assign fin_with_header_bits_payload_manager_id = io_client_finish_bits_manager_id;
  assign prb_without_header_ready = io_client_probe_ready;
  assign prb_without_header_valid = io_network_probe_valid;
  assign prb_without_header_bits_addr_block = io_network_probe_bits_payload_addr_block;
  assign prb_without_header_bits_p_type = io_network_probe_bits_payload_p_type;
  assign gnt_without_header_ready = io_client_grant_ready;
  assign gnt_without_header_valid = io_network_grant_valid;
  assign gnt_without_header_bits_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign gnt_without_header_bits_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign gnt_without_header_bits_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign gnt_without_header_bits_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign gnt_without_header_bits_g_type = io_network_grant_bits_payload_g_type;
  assign gnt_without_header_bits_data = io_network_grant_bits_payload_data;
endmodule
module TileLinkEnqueuer_4(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [2:0] io_client_acquire_bits_header_src,
  input  [2:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_header_src,
  output [2:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_header_src,
  input  [2:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [2:0] io_client_probe_bits_header_src,
  output [2:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_header_src,
  input  [2:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [2:0] io_manager_acquire_bits_header_src,
  output [2:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_header_src,
  input  [2:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_header_src,
  output [2:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [2:0] io_manager_probe_bits_header_src,
  input  [2:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_header_src,
  output [2:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_5_7774_clk;
  wire  Queue_5_7774_reset;
  wire  Queue_5_7774_io_enq_ready;
  wire  Queue_5_7774_io_enq_valid;
  wire [2:0] Queue_5_7774_io_enq_bits_header_src;
  wire [2:0] Queue_5_7774_io_enq_bits_header_dst;
  wire [25:0] Queue_5_7774_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_5_7774_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_5_7774_io_enq_bits_payload_addr_beat;
  wire  Queue_5_7774_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_5_7774_io_enq_bits_payload_a_type;
  wire [11:0] Queue_5_7774_io_enq_bits_payload_union;
  wire [63:0] Queue_5_7774_io_enq_bits_payload_data;
  wire  Queue_5_7774_io_deq_ready;
  wire  Queue_5_7774_io_deq_valid;
  wire [2:0] Queue_5_7774_io_deq_bits_header_src;
  wire [2:0] Queue_5_7774_io_deq_bits_header_dst;
  wire [25:0] Queue_5_7774_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_5_7774_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_5_7774_io_deq_bits_payload_addr_beat;
  wire  Queue_5_7774_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_5_7774_io_deq_bits_payload_a_type;
  wire [11:0] Queue_5_7774_io_deq_bits_payload_union;
  wire [63:0] Queue_5_7774_io_deq_bits_payload_data;
  wire  Queue_5_7774_io_count;
  wire  Queue_6_7897_clk;
  wire  Queue_6_7897_reset;
  wire  Queue_6_7897_io_enq_ready;
  wire  Queue_6_7897_io_enq_valid;
  wire [2:0] Queue_6_7897_io_enq_bits_header_src;
  wire [2:0] Queue_6_7897_io_enq_bits_header_dst;
  wire [25:0] Queue_6_7897_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_6_7897_io_enq_bits_payload_p_type;
  wire  Queue_6_7897_io_deq_ready;
  wire  Queue_6_7897_io_deq_valid;
  wire [2:0] Queue_6_7897_io_deq_bits_header_src;
  wire [2:0] Queue_6_7897_io_deq_bits_header_dst;
  wire [25:0] Queue_6_7897_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_6_7897_io_deq_bits_payload_p_type;
  wire  Queue_6_7897_io_count;
  wire  Queue_7_8024_clk;
  wire  Queue_7_8024_reset;
  wire  Queue_7_8024_io_enq_ready;
  wire  Queue_7_8024_io_enq_valid;
  wire [2:0] Queue_7_8024_io_enq_bits_header_src;
  wire [2:0] Queue_7_8024_io_enq_bits_header_dst;
  wire [2:0] Queue_7_8024_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_7_8024_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_7_8024_io_enq_bits_payload_client_xact_id;
  wire  Queue_7_8024_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_7_8024_io_enq_bits_payload_r_type;
  wire [63:0] Queue_7_8024_io_enq_bits_payload_data;
  wire  Queue_7_8024_io_deq_ready;
  wire  Queue_7_8024_io_deq_valid;
  wire [2:0] Queue_7_8024_io_deq_bits_header_src;
  wire [2:0] Queue_7_8024_io_deq_bits_header_dst;
  wire [2:0] Queue_7_8024_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_7_8024_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_7_8024_io_deq_bits_payload_client_xact_id;
  wire  Queue_7_8024_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_7_8024_io_deq_bits_payload_r_type;
  wire [63:0] Queue_7_8024_io_deq_bits_payload_data;
  wire [1:0] Queue_7_8024_io_count;
  wire  Queue_8_8151_clk;
  wire  Queue_8_8151_reset;
  wire  Queue_8_8151_io_enq_ready;
  wire  Queue_8_8151_io_enq_valid;
  wire [2:0] Queue_8_8151_io_enq_bits_header_src;
  wire [2:0] Queue_8_8151_io_enq_bits_header_dst;
  wire [2:0] Queue_8_8151_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_8_8151_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_8_8151_io_enq_bits_payload_manager_xact_id;
  wire  Queue_8_8151_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_8_8151_io_enq_bits_payload_g_type;
  wire [63:0] Queue_8_8151_io_enq_bits_payload_data;
  wire  Queue_8_8151_io_deq_ready;
  wire  Queue_8_8151_io_deq_valid;
  wire [2:0] Queue_8_8151_io_deq_bits_header_src;
  wire [2:0] Queue_8_8151_io_deq_bits_header_dst;
  wire [2:0] Queue_8_8151_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_8_8151_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_8_8151_io_deq_bits_payload_manager_xact_id;
  wire  Queue_8_8151_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_8_8151_io_deq_bits_payload_g_type;
  wire [63:0] Queue_8_8151_io_deq_bits_payload_data;
  wire [1:0] Queue_8_8151_io_count;
  Queue Queue_5_7774 (
    .clk(Queue_5_7774_clk),
    .reset(Queue_5_7774_reset),
    .io_enq_ready(Queue_5_7774_io_enq_ready),
    .io_enq_valid(Queue_5_7774_io_enq_valid),
    .io_enq_bits_header_src(Queue_5_7774_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_5_7774_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_5_7774_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_5_7774_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_5_7774_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_5_7774_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_5_7774_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_5_7774_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_5_7774_io_enq_bits_payload_data),
    .io_deq_ready(Queue_5_7774_io_deq_ready),
    .io_deq_valid(Queue_5_7774_io_deq_valid),
    .io_deq_bits_header_src(Queue_5_7774_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_5_7774_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_5_7774_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_5_7774_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_5_7774_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_5_7774_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_5_7774_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_5_7774_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_5_7774_io_deq_bits_payload_data),
    .io_count(Queue_5_7774_io_count)
  );
  Queue_1 Queue_6_7897 (
    .clk(Queue_6_7897_clk),
    .reset(Queue_6_7897_reset),
    .io_enq_ready(Queue_6_7897_io_enq_ready),
    .io_enq_valid(Queue_6_7897_io_enq_valid),
    .io_enq_bits_header_src(Queue_6_7897_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_6_7897_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_6_7897_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_6_7897_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_6_7897_io_deq_ready),
    .io_deq_valid(Queue_6_7897_io_deq_valid),
    .io_deq_bits_header_src(Queue_6_7897_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_6_7897_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_6_7897_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_6_7897_io_deq_bits_payload_p_type),
    .io_count(Queue_6_7897_io_count)
  );
  Queue_2 Queue_7_8024 (
    .clk(Queue_7_8024_clk),
    .reset(Queue_7_8024_reset),
    .io_enq_ready(Queue_7_8024_io_enq_ready),
    .io_enq_valid(Queue_7_8024_io_enq_valid),
    .io_enq_bits_header_src(Queue_7_8024_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_7_8024_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_7_8024_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_7_8024_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_7_8024_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_7_8024_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_7_8024_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_7_8024_io_enq_bits_payload_data),
    .io_deq_ready(Queue_7_8024_io_deq_ready),
    .io_deq_valid(Queue_7_8024_io_deq_valid),
    .io_deq_bits_header_src(Queue_7_8024_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_7_8024_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_7_8024_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_7_8024_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_7_8024_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_7_8024_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_7_8024_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_7_8024_io_deq_bits_payload_data),
    .io_count(Queue_7_8024_io_count)
  );
  Queue_3 Queue_8_8151 (
    .clk(Queue_8_8151_clk),
    .reset(Queue_8_8151_reset),
    .io_enq_ready(Queue_8_8151_io_enq_ready),
    .io_enq_valid(Queue_8_8151_io_enq_valid),
    .io_enq_bits_header_src(Queue_8_8151_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_8_8151_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_8_8151_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_8_8151_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_8_8151_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_8_8151_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_8_8151_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_8_8151_io_enq_bits_payload_data),
    .io_deq_ready(Queue_8_8151_io_deq_ready),
    .io_deq_valid(Queue_8_8151_io_deq_valid),
    .io_deq_bits_header_src(Queue_8_8151_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_8_8151_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_8_8151_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_8_8151_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_8_8151_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_8_8151_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_8_8151_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_8_8151_io_deq_bits_payload_data),
    .io_count(Queue_8_8151_io_count)
  );
  assign io_client_acquire_ready = Queue_5_7774_io_enq_ready;
  assign io_client_grant_valid = Queue_8_8151_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_8_8151_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_8_8151_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_8_8151_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_8_8151_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_8_8151_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_8_8151_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_8_8151_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_8_8151_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_6_7897_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_6_7897_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_6_7897_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_6_7897_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_6_7897_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_7_8024_io_enq_ready;
  assign io_manager_acquire_valid = Queue_5_7774_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_5_7774_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_5_7774_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_5_7774_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_5_7774_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_5_7774_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_5_7774_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_5_7774_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_5_7774_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_5_7774_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_8_8151_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_6_7897_io_enq_ready;
  assign io_manager_release_valid = Queue_7_8024_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_7_8024_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_7_8024_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_7_8024_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_7_8024_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_7_8024_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_7_8024_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_7_8024_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_7_8024_io_deq_bits_payload_data;
  assign Queue_5_7774_clk = clk;
  assign Queue_5_7774_reset = reset;
  assign Queue_5_7774_io_enq_valid = io_client_acquire_valid;
  assign Queue_5_7774_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_5_7774_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_5_7774_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_5_7774_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_5_7774_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_5_7774_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_5_7774_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_5_7774_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_5_7774_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_5_7774_io_deq_ready = io_manager_acquire_ready;
  assign Queue_6_7897_clk = clk;
  assign Queue_6_7897_reset = reset;
  assign Queue_6_7897_io_enq_valid = io_manager_probe_valid;
  assign Queue_6_7897_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_6_7897_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_6_7897_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_6_7897_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_6_7897_io_deq_ready = io_client_probe_ready;
  assign Queue_7_8024_clk = clk;
  assign Queue_7_8024_reset = reset;
  assign Queue_7_8024_io_enq_valid = io_client_release_valid;
  assign Queue_7_8024_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_7_8024_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_7_8024_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_7_8024_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_7_8024_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_7_8024_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_7_8024_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_7_8024_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_7_8024_io_deq_ready = io_manager_release_ready;
  assign Queue_8_8151_clk = clk;
  assign Queue_8_8151_reset = reset;
  assign Queue_8_8151_io_enq_valid = io_manager_grant_valid;
  assign Queue_8_8151_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_8_8151_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_8_8151_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_8_8151_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_8_8151_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_8_8151_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_8_8151_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_8_8151_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_8_8151_io_deq_ready = io_client_grant_ready;
endmodule
module FinishQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output [1:0] io_count
);
  reg [2:0] T_244_manager_xact_id [0:1];
  reg [31:0] GEN_0;
  wire [2:0] T_244_manager_xact_id_T_301_data;
  wire  T_244_manager_xact_id_T_301_addr;
  wire  T_244_manager_xact_id_T_301_en;
  wire [2:0] T_244_manager_xact_id_T_260_data;
  wire  T_244_manager_xact_id_T_260_addr;
  wire  T_244_manager_xact_id_T_260_mask;
  wire  T_244_manager_xact_id_T_260_en;
  reg  T_244_manager_id [0:1];
  reg [31:0] GEN_1;
  wire  T_244_manager_id_T_301_data;
  wire  T_244_manager_id_T_301_addr;
  wire  T_244_manager_id_T_301_en;
  wire  T_244_manager_id_T_260_data;
  wire  T_244_manager_id_T_260_addr;
  wire  T_244_manager_id_T_260_mask;
  wire  T_244_manager_id_T_260_en;
  reg  T_246;
  reg [31:0] GEN_2;
  reg  T_248;
  reg [31:0] GEN_3;
  reg  T_250;
  reg [31:0] GEN_4;
  wire  T_251;
  wire  T_253;
  wire  T_254;
  wire  T_255;
  wire  T_256;
  wire  T_257;
  wire  T_258;
  wire  T_259;
  wire [1:0] T_289;
  wire  T_290;
  wire  GEN_7;
  wire [1:0] T_294;
  wire  T_295;
  wire  GEN_8;
  wire  T_296;
  wire  GEN_9;
  wire  T_298;
  wire  T_300;
  wire [1:0] T_327;
  wire  T_328;
  wire  T_329;
  wire [1:0] T_330;
  assign io_enq_ready = T_300;
  assign io_deq_valid = T_298;
  assign io_deq_bits_manager_xact_id = T_244_manager_xact_id_T_301_data;
  assign io_deq_bits_manager_id = T_244_manager_id_T_301_data;
  assign io_count = T_330;
  assign T_244_manager_xact_id_T_301_addr = T_248;
  assign T_244_manager_xact_id_T_301_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_xact_id_T_301_data = T_244_manager_xact_id[T_244_manager_xact_id_T_301_addr];
  `else
  assign T_244_manager_xact_id_T_301_data = T_244_manager_xact_id_T_301_addr >= 2'h2 ? $random : T_244_manager_xact_id[T_244_manager_xact_id_T_301_addr];
  `endif
  assign T_244_manager_xact_id_T_260_data = io_enq_bits_manager_xact_id;
  assign T_244_manager_xact_id_T_260_addr = T_246;
  assign T_244_manager_xact_id_T_260_mask = T_257;
  assign T_244_manager_xact_id_T_260_en = T_257;
  assign T_244_manager_id_T_301_addr = T_248;
  assign T_244_manager_id_T_301_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_id_T_301_data = T_244_manager_id[T_244_manager_id_T_301_addr];
  `else
  assign T_244_manager_id_T_301_data = T_244_manager_id_T_301_addr >= 2'h2 ? $random : T_244_manager_id[T_244_manager_id_T_301_addr];
  `endif
  assign T_244_manager_id_T_260_data = io_enq_bits_manager_id;
  assign T_244_manager_id_T_260_addr = T_246;
  assign T_244_manager_id_T_260_mask = T_257;
  assign T_244_manager_id_T_260_en = T_257;
  assign T_251 = T_246 == T_248;
  assign T_253 = T_250 == 1'h0;
  assign T_254 = T_251 & T_253;
  assign T_255 = T_251 & T_250;
  assign T_256 = io_enq_ready & io_enq_valid;
  assign T_257 = T_256;
  assign T_258 = io_deq_ready & io_deq_valid;
  assign T_259 = T_258;
  assign T_289 = T_246 + 1'h1;
  assign T_290 = T_289[0:0];
  assign GEN_7 = T_257 ? T_290 : T_246;
  assign T_294 = T_248 + 1'h1;
  assign T_295 = T_294[0:0];
  assign GEN_8 = T_259 ? T_295 : T_248;
  assign T_296 = T_257 != T_259;
  assign GEN_9 = T_296 ? T_257 : T_250;
  assign T_298 = T_254 == 1'h0;
  assign T_300 = T_255 == 1'h0;
  assign T_327 = T_246 - T_248;
  assign T_328 = T_327[0:0];
  assign T_329 = T_250 & T_251;
  assign T_330 = {T_329,T_328};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    T_244_manager_xact_id[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    T_244_manager_id[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  T_246 = GEN_2[0:0];
  GEN_3 = {1{$random}};
  T_248 = GEN_3[0:0];
  GEN_4 = {1{$random}};
  T_250 = GEN_4[0:0];
  end
`endif
  always @(posedge clk) begin
    if(T_244_manager_xact_id_T_260_en & T_244_manager_xact_id_T_260_mask) begin
      T_244_manager_xact_id[T_244_manager_xact_id_T_260_addr] <= T_244_manager_xact_id_T_260_data;
    end
    if(T_244_manager_id_T_260_en & T_244_manager_id_T_260_mask) begin
      T_244_manager_id[T_244_manager_id_T_260_addr] <= T_244_manager_id_T_260_data;
    end
    if(reset) begin
      T_246 <= 1'h0;
    end else begin
      T_246 <= GEN_7;
    end
    if(reset) begin
      T_248 <= 1'h0;
    end else begin
      T_248 <= GEN_8;
    end
    if(reset) begin
      T_250 <= 1'h0;
    end else begin
      T_250 <= GEN_9;
    end
  end
endmodule
module FinishUnit(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [2:0] io_grant_bits_header_src,
  input  [2:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input  [1:0] io_grant_bits_payload_client_xact_id,
  input  [2:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output [1:0] io_refill_bits_client_xact_id,
  output [2:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [2:0] io_finish_bits_header_src,
  output [2:0] io_finish_bits_header_dst,
  output [2:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1173;
  wire [2:0] T_1182_0;
  wire [3:0] GEN_1;
  wire  T_1184;
  wire [1:0] T_1192_0;
  wire [1:0] T_1192_1;
  wire [3:0] GEN_2;
  wire  T_1194;
  wire [3:0] GEN_3;
  wire  T_1195;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  reg [2:0] T_1203;
  reg [31:0] GEN_9;
  wire  T_1205;
  wire [2:0] GEN_4;
  wire [3:0] T_1207;
  wire [2:0] T_1208;
  wire [2:0] GEN_0;
  wire  T_1209;
  wire  T_1211;
  wire  FinishQueue_1238_clk;
  wire  FinishQueue_1238_reset;
  wire  FinishQueue_1238_io_enq_ready;
  wire  FinishQueue_1238_io_enq_valid;
  wire [2:0] FinishQueue_1238_io_enq_bits_manager_xact_id;
  wire  FinishQueue_1238_io_enq_bits_manager_id;
  wire  FinishQueue_1238_io_deq_ready;
  wire  FinishQueue_1238_io_deq_valid;
  wire [2:0] FinishQueue_1238_io_deq_bits_manager_xact_id;
  wire  FinishQueue_1238_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_1238_io_count;
  wire [3:0] GEN_5;
  wire  T_1244;
  wire  T_1245;
  wire  T_1247;
  wire  T_1249;
  wire [2:0] T_1257_0;
  wire [3:0] GEN_6;
  wire  T_1259;
  wire [1:0] T_1267_0;
  wire [1:0] T_1267_1;
  wire [3:0] GEN_7;
  wire  T_1269;
  wire [3:0] GEN_8;
  wire  T_1270;
  wire  T_1273;
  wire  T_1274;
  wire  T_1277;
  wire  T_1278;
  wire  T_1279;
  wire [2:0] T_1305_manager_xact_id;
  wire  T_1341;
  wire  T_1342;
  wire  T_1343;
  wire  T_1356;
  FinishQueue FinishQueue_1238 (
    .clk(FinishQueue_1238_clk),
    .reset(FinishQueue_1238_reset),
    .io_enq_ready(FinishQueue_1238_io_enq_ready),
    .io_enq_valid(FinishQueue_1238_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_1238_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_1238_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_1238_io_deq_ready),
    .io_deq_valid(FinishQueue_1238_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_1238_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_1238_io_deq_bits_manager_id),
    .io_count(FinishQueue_1238_io_count)
  );
  assign io_grant_ready = T_1356;
  assign io_refill_valid = T_1343;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_1238_io_deq_valid;
  assign io_finish_bits_header_src = {{2'd0}, 1'h1};
  assign io_finish_bits_header_dst = {{2'd0}, FinishQueue_1238_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_1238_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_1238_io_enq_ready;
  assign T_1173 = io_grant_ready & io_grant_valid;
  assign T_1182_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1182_0};
  assign T_1184 = GEN_1 == io_grant_bits_payload_g_type;
  assign T_1192_0 = 2'h0;
  assign T_1192_1 = 2'h1;
  assign GEN_2 = {{2'd0}, T_1192_0};
  assign T_1194 = GEN_2 == io_grant_bits_payload_g_type;
  assign GEN_3 = {{2'd0}, T_1192_1};
  assign T_1195 = GEN_3 == io_grant_bits_payload_g_type;
  assign T_1198 = T_1194 | T_1195;
  assign T_1199 = io_grant_bits_payload_is_builtin_type ? T_1184 : T_1198;
  assign T_1201 = T_1173 & T_1199;
  assign T_1205 = T_1203 == 3'h7;
  assign GEN_4 = {{2'd0}, 1'h1};
  assign T_1207 = T_1203 + GEN_4;
  assign T_1208 = T_1207[2:0];
  assign GEN_0 = T_1201 ? T_1208 : T_1203;
  assign T_1209 = T_1201 & T_1205;
  assign T_1211 = T_1199 ? T_1209 : T_1173;
  assign FinishQueue_1238_clk = clk;
  assign FinishQueue_1238_reset = reset;
  assign FinishQueue_1238_io_enq_valid = T_1279;
  assign FinishQueue_1238_io_enq_bits_manager_xact_id = T_1305_manager_xact_id;
  assign FinishQueue_1238_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_1238_io_deq_ready = io_finish_ready;
  assign GEN_5 = {{1'd0}, 3'h0};
  assign T_1244 = io_grant_bits_payload_g_type == GEN_5;
  assign T_1245 = io_grant_bits_payload_is_builtin_type & T_1244;
  assign T_1247 = T_1245 == 1'h0;
  assign T_1249 = T_1173 & T_1247;
  assign T_1257_0 = 3'h5;
  assign GEN_6 = {{1'd0}, T_1257_0};
  assign T_1259 = GEN_6 == io_grant_bits_payload_g_type;
  assign T_1267_0 = 2'h0;
  assign T_1267_1 = 2'h1;
  assign GEN_7 = {{2'd0}, T_1267_0};
  assign T_1269 = GEN_7 == io_grant_bits_payload_g_type;
  assign GEN_8 = {{2'd0}, T_1267_1};
  assign T_1270 = GEN_8 == io_grant_bits_payload_g_type;
  assign T_1273 = T_1269 | T_1270;
  assign T_1274 = io_grant_bits_payload_is_builtin_type ? T_1259 : T_1273;
  assign T_1277 = T_1274 == 1'h0;
  assign T_1278 = T_1277 | T_1211;
  assign T_1279 = T_1249 & T_1278;
  assign T_1305_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1341 = T_1247 == 1'h0;
  assign T_1342 = FinishQueue_1238_io_enq_ready | T_1341;
  assign T_1343 = T_1342 & io_grant_valid;
  assign T_1356 = T_1342 & io_refill_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  T_1203 = GEN_9[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1203 <= 3'h0;
    end else begin
      T_1203 <= GEN_0;
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [2:0] io_network_acquire_bits_header_src,
  output [2:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [2:0] io_network_grant_bits_header_src,
  input  [2:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [2:0] io_network_finish_bits_header_src,
  output [2:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [2:0] io_network_probe_bits_header_src,
  input  [2:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [2:0] io_network_release_bits_header_src,
  output [2:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [2:0] finisher_io_grant_bits_header_src;
  wire [2:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire [1:0] finisher_io_grant_bits_payload_client_xact_id;
  wire [2:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire [1:0] finisher_io_refill_bits_client_xact_id;
  wire [2:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [2:0] finisher_io_finish_bits_header_src;
  wire [2:0] finisher_io_finish_bits_header_dst;
  wire [2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [2:0] acq_with_header_bits_header_src;
  wire [2:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3765;
  wire  T_3767;
  wire  T_3773;
  wire  T_3774;
  wire  T_3775;
  reg [2:0] GEN_1;
  reg [31:0] GEN_9;
  reg [2:0] GEN_2;
  reg [31:0] GEN_10;
  reg [2:0] GEN_3;
  reg [31:0] GEN_11;
  reg [25:0] GEN_4;
  reg [31:0] GEN_12;
  reg [1:0] GEN_5;
  reg [31:0] GEN_13;
  reg  GEN_6;
  reg [31:0] GEN_14;
  reg [2:0] GEN_7;
  reg [31:0] GEN_15;
  reg [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3774;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3775;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = {{2'd0}, 1'h1};
  assign acq_with_header_bits_header_dst = {{2'd0}, T_3773};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3765 = GEN_0 << 6;
  assign T_3767 = 32'h80000000 <= T_3765;
  assign T_3773 = T_3767 ? 1'h0 : 1'h1;
  assign T_3774 = acq_with_header_valid & finisher_io_ready;
  assign T_3775 = io_network_acquire_ready & finisher_io_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  GEN_1 = GEN_9[2:0];
  GEN_10 = {1{$random}};
  GEN_2 = GEN_10[2:0];
  GEN_11 = {1{$random}};
  GEN_3 = GEN_11[2:0];
  GEN_12 = {1{$random}};
  GEN_4 = GEN_12[25:0];
  GEN_13 = {1{$random}};
  GEN_5 = GEN_13[1:0];
  GEN_14 = {1{$random}};
  GEN_6 = GEN_14[0:0];
  GEN_15 = {1{$random}};
  GEN_7 = GEN_15[2:0];
  GEN_16 = {2{$random}};
  GEN_8 = GEN_16[63:0];
  end
`endif
endmodule
module TileLinkEnqueuer_9(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [2:0] io_client_acquire_bits_header_src,
  input  [2:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_header_src,
  output [2:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_header_src,
  input  [2:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [2:0] io_client_probe_bits_header_src,
  output [2:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_header_src,
  input  [2:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [2:0] io_manager_acquire_bits_header_src,
  output [2:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_header_src,
  input  [2:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_header_src,
  output [2:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [2:0] io_manager_probe_bits_header_src,
  input  [2:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_header_src,
  output [2:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  wire  Queue_10_7774_clk;
  wire  Queue_10_7774_reset;
  wire  Queue_10_7774_io_enq_ready;
  wire  Queue_10_7774_io_enq_valid;
  wire [2:0] Queue_10_7774_io_enq_bits_header_src;
  wire [2:0] Queue_10_7774_io_enq_bits_header_dst;
  wire [25:0] Queue_10_7774_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_10_7774_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_10_7774_io_enq_bits_payload_addr_beat;
  wire  Queue_10_7774_io_enq_bits_payload_is_builtin_type;
  wire [2:0] Queue_10_7774_io_enq_bits_payload_a_type;
  wire [11:0] Queue_10_7774_io_enq_bits_payload_union;
  wire [63:0] Queue_10_7774_io_enq_bits_payload_data;
  wire  Queue_10_7774_io_deq_ready;
  wire  Queue_10_7774_io_deq_valid;
  wire [2:0] Queue_10_7774_io_deq_bits_header_src;
  wire [2:0] Queue_10_7774_io_deq_bits_header_dst;
  wire [25:0] Queue_10_7774_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_10_7774_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_10_7774_io_deq_bits_payload_addr_beat;
  wire  Queue_10_7774_io_deq_bits_payload_is_builtin_type;
  wire [2:0] Queue_10_7774_io_deq_bits_payload_a_type;
  wire [11:0] Queue_10_7774_io_deq_bits_payload_union;
  wire [63:0] Queue_10_7774_io_deq_bits_payload_data;
  wire  Queue_10_7774_io_count;
  wire  Queue_11_7897_clk;
  wire  Queue_11_7897_reset;
  wire  Queue_11_7897_io_enq_ready;
  wire  Queue_11_7897_io_enq_valid;
  wire [2:0] Queue_11_7897_io_enq_bits_header_src;
  wire [2:0] Queue_11_7897_io_enq_bits_header_dst;
  wire [25:0] Queue_11_7897_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_11_7897_io_enq_bits_payload_p_type;
  wire  Queue_11_7897_io_deq_ready;
  wire  Queue_11_7897_io_deq_valid;
  wire [2:0] Queue_11_7897_io_deq_bits_header_src;
  wire [2:0] Queue_11_7897_io_deq_bits_header_dst;
  wire [25:0] Queue_11_7897_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_11_7897_io_deq_bits_payload_p_type;
  wire  Queue_11_7897_io_count;
  wire  Queue_12_8024_clk;
  wire  Queue_12_8024_reset;
  wire  Queue_12_8024_io_enq_ready;
  wire  Queue_12_8024_io_enq_valid;
  wire [2:0] Queue_12_8024_io_enq_bits_header_src;
  wire [2:0] Queue_12_8024_io_enq_bits_header_dst;
  wire [2:0] Queue_12_8024_io_enq_bits_payload_addr_beat;
  wire [25:0] Queue_12_8024_io_enq_bits_payload_addr_block;
  wire [1:0] Queue_12_8024_io_enq_bits_payload_client_xact_id;
  wire  Queue_12_8024_io_enq_bits_payload_voluntary;
  wire [2:0] Queue_12_8024_io_enq_bits_payload_r_type;
  wire [63:0] Queue_12_8024_io_enq_bits_payload_data;
  wire  Queue_12_8024_io_deq_ready;
  wire  Queue_12_8024_io_deq_valid;
  wire [2:0] Queue_12_8024_io_deq_bits_header_src;
  wire [2:0] Queue_12_8024_io_deq_bits_header_dst;
  wire [2:0] Queue_12_8024_io_deq_bits_payload_addr_beat;
  wire [25:0] Queue_12_8024_io_deq_bits_payload_addr_block;
  wire [1:0] Queue_12_8024_io_deq_bits_payload_client_xact_id;
  wire  Queue_12_8024_io_deq_bits_payload_voluntary;
  wire [2:0] Queue_12_8024_io_deq_bits_payload_r_type;
  wire [63:0] Queue_12_8024_io_deq_bits_payload_data;
  wire [1:0] Queue_12_8024_io_count;
  wire  Queue_13_8151_clk;
  wire  Queue_13_8151_reset;
  wire  Queue_13_8151_io_enq_ready;
  wire  Queue_13_8151_io_enq_valid;
  wire [2:0] Queue_13_8151_io_enq_bits_header_src;
  wire [2:0] Queue_13_8151_io_enq_bits_header_dst;
  wire [2:0] Queue_13_8151_io_enq_bits_payload_addr_beat;
  wire [1:0] Queue_13_8151_io_enq_bits_payload_client_xact_id;
  wire [2:0] Queue_13_8151_io_enq_bits_payload_manager_xact_id;
  wire  Queue_13_8151_io_enq_bits_payload_is_builtin_type;
  wire [3:0] Queue_13_8151_io_enq_bits_payload_g_type;
  wire [63:0] Queue_13_8151_io_enq_bits_payload_data;
  wire  Queue_13_8151_io_deq_ready;
  wire  Queue_13_8151_io_deq_valid;
  wire [2:0] Queue_13_8151_io_deq_bits_header_src;
  wire [2:0] Queue_13_8151_io_deq_bits_header_dst;
  wire [2:0] Queue_13_8151_io_deq_bits_payload_addr_beat;
  wire [1:0] Queue_13_8151_io_deq_bits_payload_client_xact_id;
  wire [2:0] Queue_13_8151_io_deq_bits_payload_manager_xact_id;
  wire  Queue_13_8151_io_deq_bits_payload_is_builtin_type;
  wire [3:0] Queue_13_8151_io_deq_bits_payload_g_type;
  wire [63:0] Queue_13_8151_io_deq_bits_payload_data;
  wire [1:0] Queue_13_8151_io_count;
  Queue Queue_10_7774 (
    .clk(Queue_10_7774_clk),
    .reset(Queue_10_7774_reset),
    .io_enq_ready(Queue_10_7774_io_enq_ready),
    .io_enq_valid(Queue_10_7774_io_enq_valid),
    .io_enq_bits_header_src(Queue_10_7774_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_10_7774_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_10_7774_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_10_7774_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_addr_beat(Queue_10_7774_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_is_builtin_type(Queue_10_7774_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_a_type(Queue_10_7774_io_enq_bits_payload_a_type),
    .io_enq_bits_payload_union(Queue_10_7774_io_enq_bits_payload_union),
    .io_enq_bits_payload_data(Queue_10_7774_io_enq_bits_payload_data),
    .io_deq_ready(Queue_10_7774_io_deq_ready),
    .io_deq_valid(Queue_10_7774_io_deq_valid),
    .io_deq_bits_header_src(Queue_10_7774_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_10_7774_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_10_7774_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_10_7774_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_addr_beat(Queue_10_7774_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_is_builtin_type(Queue_10_7774_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_a_type(Queue_10_7774_io_deq_bits_payload_a_type),
    .io_deq_bits_payload_union(Queue_10_7774_io_deq_bits_payload_union),
    .io_deq_bits_payload_data(Queue_10_7774_io_deq_bits_payload_data),
    .io_count(Queue_10_7774_io_count)
  );
  Queue_1 Queue_11_7897 (
    .clk(Queue_11_7897_clk),
    .reset(Queue_11_7897_reset),
    .io_enq_ready(Queue_11_7897_io_enq_ready),
    .io_enq_valid(Queue_11_7897_io_enq_valid),
    .io_enq_bits_header_src(Queue_11_7897_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_11_7897_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_block(Queue_11_7897_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_p_type(Queue_11_7897_io_enq_bits_payload_p_type),
    .io_deq_ready(Queue_11_7897_io_deq_ready),
    .io_deq_valid(Queue_11_7897_io_deq_valid),
    .io_deq_bits_header_src(Queue_11_7897_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_11_7897_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_block(Queue_11_7897_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_p_type(Queue_11_7897_io_deq_bits_payload_p_type),
    .io_count(Queue_11_7897_io_count)
  );
  Queue_2 Queue_12_8024 (
    .clk(Queue_12_8024_clk),
    .reset(Queue_12_8024_reset),
    .io_enq_ready(Queue_12_8024_io_enq_ready),
    .io_enq_valid(Queue_12_8024_io_enq_valid),
    .io_enq_bits_header_src(Queue_12_8024_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_12_8024_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_12_8024_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_addr_block(Queue_12_8024_io_enq_bits_payload_addr_block),
    .io_enq_bits_payload_client_xact_id(Queue_12_8024_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_voluntary(Queue_12_8024_io_enq_bits_payload_voluntary),
    .io_enq_bits_payload_r_type(Queue_12_8024_io_enq_bits_payload_r_type),
    .io_enq_bits_payload_data(Queue_12_8024_io_enq_bits_payload_data),
    .io_deq_ready(Queue_12_8024_io_deq_ready),
    .io_deq_valid(Queue_12_8024_io_deq_valid),
    .io_deq_bits_header_src(Queue_12_8024_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_12_8024_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_12_8024_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_addr_block(Queue_12_8024_io_deq_bits_payload_addr_block),
    .io_deq_bits_payload_client_xact_id(Queue_12_8024_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_voluntary(Queue_12_8024_io_deq_bits_payload_voluntary),
    .io_deq_bits_payload_r_type(Queue_12_8024_io_deq_bits_payload_r_type),
    .io_deq_bits_payload_data(Queue_12_8024_io_deq_bits_payload_data),
    .io_count(Queue_12_8024_io_count)
  );
  Queue_3 Queue_13_8151 (
    .clk(Queue_13_8151_clk),
    .reset(Queue_13_8151_reset),
    .io_enq_ready(Queue_13_8151_io_enq_ready),
    .io_enq_valid(Queue_13_8151_io_enq_valid),
    .io_enq_bits_header_src(Queue_13_8151_io_enq_bits_header_src),
    .io_enq_bits_header_dst(Queue_13_8151_io_enq_bits_header_dst),
    .io_enq_bits_payload_addr_beat(Queue_13_8151_io_enq_bits_payload_addr_beat),
    .io_enq_bits_payload_client_xact_id(Queue_13_8151_io_enq_bits_payload_client_xact_id),
    .io_enq_bits_payload_manager_xact_id(Queue_13_8151_io_enq_bits_payload_manager_xact_id),
    .io_enq_bits_payload_is_builtin_type(Queue_13_8151_io_enq_bits_payload_is_builtin_type),
    .io_enq_bits_payload_g_type(Queue_13_8151_io_enq_bits_payload_g_type),
    .io_enq_bits_payload_data(Queue_13_8151_io_enq_bits_payload_data),
    .io_deq_ready(Queue_13_8151_io_deq_ready),
    .io_deq_valid(Queue_13_8151_io_deq_valid),
    .io_deq_bits_header_src(Queue_13_8151_io_deq_bits_header_src),
    .io_deq_bits_header_dst(Queue_13_8151_io_deq_bits_header_dst),
    .io_deq_bits_payload_addr_beat(Queue_13_8151_io_deq_bits_payload_addr_beat),
    .io_deq_bits_payload_client_xact_id(Queue_13_8151_io_deq_bits_payload_client_xact_id),
    .io_deq_bits_payload_manager_xact_id(Queue_13_8151_io_deq_bits_payload_manager_xact_id),
    .io_deq_bits_payload_is_builtin_type(Queue_13_8151_io_deq_bits_payload_is_builtin_type),
    .io_deq_bits_payload_g_type(Queue_13_8151_io_deq_bits_payload_g_type),
    .io_deq_bits_payload_data(Queue_13_8151_io_deq_bits_payload_data),
    .io_count(Queue_13_8151_io_count)
  );
  assign io_client_acquire_ready = Queue_10_7774_io_enq_ready;
  assign io_client_grant_valid = Queue_13_8151_io_deq_valid;
  assign io_client_grant_bits_header_src = Queue_13_8151_io_deq_bits_header_src;
  assign io_client_grant_bits_header_dst = Queue_13_8151_io_deq_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = Queue_13_8151_io_deq_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = Queue_13_8151_io_deq_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = Queue_13_8151_io_deq_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = Queue_13_8151_io_deq_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = Queue_13_8151_io_deq_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = Queue_13_8151_io_deq_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = Queue_11_7897_io_deq_valid;
  assign io_client_probe_bits_header_src = Queue_11_7897_io_deq_bits_header_src;
  assign io_client_probe_bits_header_dst = Queue_11_7897_io_deq_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = Queue_11_7897_io_deq_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = Queue_11_7897_io_deq_bits_payload_p_type;
  assign io_client_release_ready = Queue_12_8024_io_enq_ready;
  assign io_manager_acquire_valid = Queue_10_7774_io_deq_valid;
  assign io_manager_acquire_bits_header_src = Queue_10_7774_io_deq_bits_header_src;
  assign io_manager_acquire_bits_header_dst = Queue_10_7774_io_deq_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = Queue_10_7774_io_deq_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = Queue_10_7774_io_deq_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = Queue_10_7774_io_deq_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = Queue_10_7774_io_deq_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = Queue_10_7774_io_deq_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = Queue_10_7774_io_deq_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = Queue_10_7774_io_deq_bits_payload_data;
  assign io_manager_grant_ready = Queue_13_8151_io_enq_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = Queue_11_7897_io_enq_ready;
  assign io_manager_release_valid = Queue_12_8024_io_deq_valid;
  assign io_manager_release_bits_header_src = Queue_12_8024_io_deq_bits_header_src;
  assign io_manager_release_bits_header_dst = Queue_12_8024_io_deq_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = Queue_12_8024_io_deq_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = Queue_12_8024_io_deq_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = Queue_12_8024_io_deq_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = Queue_12_8024_io_deq_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = Queue_12_8024_io_deq_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = Queue_12_8024_io_deq_bits_payload_data;
  assign Queue_10_7774_clk = clk;
  assign Queue_10_7774_reset = reset;
  assign Queue_10_7774_io_enq_valid = io_client_acquire_valid;
  assign Queue_10_7774_io_enq_bits_header_src = io_client_acquire_bits_header_src;
  assign Queue_10_7774_io_enq_bits_header_dst = io_client_acquire_bits_header_dst;
  assign Queue_10_7774_io_enq_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign Queue_10_7774_io_enq_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign Queue_10_7774_io_enq_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign Queue_10_7774_io_enq_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign Queue_10_7774_io_enq_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign Queue_10_7774_io_enq_bits_payload_union = io_client_acquire_bits_payload_union;
  assign Queue_10_7774_io_enq_bits_payload_data = io_client_acquire_bits_payload_data;
  assign Queue_10_7774_io_deq_ready = io_manager_acquire_ready;
  assign Queue_11_7897_clk = clk;
  assign Queue_11_7897_reset = reset;
  assign Queue_11_7897_io_enq_valid = io_manager_probe_valid;
  assign Queue_11_7897_io_enq_bits_header_src = io_manager_probe_bits_header_src;
  assign Queue_11_7897_io_enq_bits_header_dst = io_manager_probe_bits_header_dst;
  assign Queue_11_7897_io_enq_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign Queue_11_7897_io_enq_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign Queue_11_7897_io_deq_ready = io_client_probe_ready;
  assign Queue_12_8024_clk = clk;
  assign Queue_12_8024_reset = reset;
  assign Queue_12_8024_io_enq_valid = io_client_release_valid;
  assign Queue_12_8024_io_enq_bits_header_src = io_client_release_bits_header_src;
  assign Queue_12_8024_io_enq_bits_header_dst = io_client_release_bits_header_dst;
  assign Queue_12_8024_io_enq_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign Queue_12_8024_io_enq_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign Queue_12_8024_io_enq_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign Queue_12_8024_io_enq_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign Queue_12_8024_io_enq_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign Queue_12_8024_io_enq_bits_payload_data = io_client_release_bits_payload_data;
  assign Queue_12_8024_io_deq_ready = io_manager_release_ready;
  assign Queue_13_8151_clk = clk;
  assign Queue_13_8151_reset = reset;
  assign Queue_13_8151_io_enq_valid = io_manager_grant_valid;
  assign Queue_13_8151_io_enq_bits_header_src = io_manager_grant_bits_header_src;
  assign Queue_13_8151_io_enq_bits_header_dst = io_manager_grant_bits_header_dst;
  assign Queue_13_8151_io_enq_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign Queue_13_8151_io_enq_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign Queue_13_8151_io_enq_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign Queue_13_8151_io_enq_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign Queue_13_8151_io_enq_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign Queue_13_8151_io_enq_bits_payload_data = io_manager_grant_bits_payload_data;
  assign Queue_13_8151_io_deq_ready = io_client_grant_ready;
endmodule
module FinishUnit_15(
  input   clk,
  input   reset,
  output  io_grant_ready,
  input   io_grant_valid,
  input  [2:0] io_grant_bits_header_src,
  input  [2:0] io_grant_bits_header_dst,
  input  [2:0] io_grant_bits_payload_addr_beat,
  input  [1:0] io_grant_bits_payload_client_xact_id,
  input  [2:0] io_grant_bits_payload_manager_xact_id,
  input   io_grant_bits_payload_is_builtin_type,
  input  [3:0] io_grant_bits_payload_g_type,
  input  [63:0] io_grant_bits_payload_data,
  input   io_refill_ready,
  output  io_refill_valid,
  output [2:0] io_refill_bits_addr_beat,
  output [1:0] io_refill_bits_client_xact_id,
  output [2:0] io_refill_bits_manager_xact_id,
  output  io_refill_bits_is_builtin_type,
  output [3:0] io_refill_bits_g_type,
  output [63:0] io_refill_bits_data,
  input   io_finish_ready,
  output  io_finish_valid,
  output [2:0] io_finish_bits_header_src,
  output [2:0] io_finish_bits_header_dst,
  output [2:0] io_finish_bits_payload_manager_xact_id,
  output  io_ready
);
  wire  T_1173;
  wire [2:0] T_1182_0;
  wire [3:0] GEN_1;
  wire  T_1184;
  wire [1:0] T_1192_0;
  wire [1:0] T_1192_1;
  wire [3:0] GEN_2;
  wire  T_1194;
  wire [3:0] GEN_3;
  wire  T_1195;
  wire  T_1198;
  wire  T_1199;
  wire  T_1201;
  reg [2:0] T_1203;
  reg [31:0] GEN_9;
  wire  T_1205;
  wire [2:0] GEN_4;
  wire [3:0] T_1207;
  wire [2:0] T_1208;
  wire [2:0] GEN_0;
  wire  T_1209;
  wire  T_1211;
  wire  FinishQueue_16_1238_clk;
  wire  FinishQueue_16_1238_reset;
  wire  FinishQueue_16_1238_io_enq_ready;
  wire  FinishQueue_16_1238_io_enq_valid;
  wire [2:0] FinishQueue_16_1238_io_enq_bits_manager_xact_id;
  wire  FinishQueue_16_1238_io_enq_bits_manager_id;
  wire  FinishQueue_16_1238_io_deq_ready;
  wire  FinishQueue_16_1238_io_deq_valid;
  wire [2:0] FinishQueue_16_1238_io_deq_bits_manager_xact_id;
  wire  FinishQueue_16_1238_io_deq_bits_manager_id;
  wire [1:0] FinishQueue_16_1238_io_count;
  wire [3:0] GEN_5;
  wire  T_1244;
  wire  T_1245;
  wire  T_1247;
  wire  T_1249;
  wire [2:0] T_1257_0;
  wire [3:0] GEN_6;
  wire  T_1259;
  wire [1:0] T_1267_0;
  wire [1:0] T_1267_1;
  wire [3:0] GEN_7;
  wire  T_1269;
  wire [3:0] GEN_8;
  wire  T_1270;
  wire  T_1273;
  wire  T_1274;
  wire  T_1277;
  wire  T_1278;
  wire  T_1279;
  wire [2:0] T_1305_manager_xact_id;
  wire  T_1341;
  wire  T_1342;
  wire  T_1343;
  wire  T_1356;
  FinishQueue FinishQueue_16_1238 (
    .clk(FinishQueue_16_1238_clk),
    .reset(FinishQueue_16_1238_reset),
    .io_enq_ready(FinishQueue_16_1238_io_enq_ready),
    .io_enq_valid(FinishQueue_16_1238_io_enq_valid),
    .io_enq_bits_manager_xact_id(FinishQueue_16_1238_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(FinishQueue_16_1238_io_enq_bits_manager_id),
    .io_deq_ready(FinishQueue_16_1238_io_deq_ready),
    .io_deq_valid(FinishQueue_16_1238_io_deq_valid),
    .io_deq_bits_manager_xact_id(FinishQueue_16_1238_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(FinishQueue_16_1238_io_deq_bits_manager_id),
    .io_count(FinishQueue_16_1238_io_count)
  );
  assign io_grant_ready = T_1356;
  assign io_refill_valid = T_1343;
  assign io_refill_bits_addr_beat = io_grant_bits_payload_addr_beat;
  assign io_refill_bits_client_xact_id = io_grant_bits_payload_client_xact_id;
  assign io_refill_bits_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign io_refill_bits_is_builtin_type = io_grant_bits_payload_is_builtin_type;
  assign io_refill_bits_g_type = io_grant_bits_payload_g_type;
  assign io_refill_bits_data = io_grant_bits_payload_data;
  assign io_finish_valid = FinishQueue_16_1238_io_deq_valid;
  assign io_finish_bits_header_src = {{1'd0}, 2'h2};
  assign io_finish_bits_header_dst = {{2'd0}, FinishQueue_16_1238_io_deq_bits_manager_id};
  assign io_finish_bits_payload_manager_xact_id = FinishQueue_16_1238_io_deq_bits_manager_xact_id;
  assign io_ready = FinishQueue_16_1238_io_enq_ready;
  assign T_1173 = io_grant_ready & io_grant_valid;
  assign T_1182_0 = 3'h5;
  assign GEN_1 = {{1'd0}, T_1182_0};
  assign T_1184 = GEN_1 == io_grant_bits_payload_g_type;
  assign T_1192_0 = 2'h0;
  assign T_1192_1 = 2'h1;
  assign GEN_2 = {{2'd0}, T_1192_0};
  assign T_1194 = GEN_2 == io_grant_bits_payload_g_type;
  assign GEN_3 = {{2'd0}, T_1192_1};
  assign T_1195 = GEN_3 == io_grant_bits_payload_g_type;
  assign T_1198 = T_1194 | T_1195;
  assign T_1199 = io_grant_bits_payload_is_builtin_type ? T_1184 : T_1198;
  assign T_1201 = T_1173 & T_1199;
  assign T_1205 = T_1203 == 3'h7;
  assign GEN_4 = {{2'd0}, 1'h1};
  assign T_1207 = T_1203 + GEN_4;
  assign T_1208 = T_1207[2:0];
  assign GEN_0 = T_1201 ? T_1208 : T_1203;
  assign T_1209 = T_1201 & T_1205;
  assign T_1211 = T_1199 ? T_1209 : T_1173;
  assign FinishQueue_16_1238_clk = clk;
  assign FinishQueue_16_1238_reset = reset;
  assign FinishQueue_16_1238_io_enq_valid = T_1279;
  assign FinishQueue_16_1238_io_enq_bits_manager_xact_id = T_1305_manager_xact_id;
  assign FinishQueue_16_1238_io_enq_bits_manager_id = io_grant_bits_header_src[0];
  assign FinishQueue_16_1238_io_deq_ready = io_finish_ready;
  assign GEN_5 = {{1'd0}, 3'h0};
  assign T_1244 = io_grant_bits_payload_g_type == GEN_5;
  assign T_1245 = io_grant_bits_payload_is_builtin_type & T_1244;
  assign T_1247 = T_1245 == 1'h0;
  assign T_1249 = T_1173 & T_1247;
  assign T_1257_0 = 3'h5;
  assign GEN_6 = {{1'd0}, T_1257_0};
  assign T_1259 = GEN_6 == io_grant_bits_payload_g_type;
  assign T_1267_0 = 2'h0;
  assign T_1267_1 = 2'h1;
  assign GEN_7 = {{2'd0}, T_1267_0};
  assign T_1269 = GEN_7 == io_grant_bits_payload_g_type;
  assign GEN_8 = {{2'd0}, T_1267_1};
  assign T_1270 = GEN_8 == io_grant_bits_payload_g_type;
  assign T_1273 = T_1269 | T_1270;
  assign T_1274 = io_grant_bits_payload_is_builtin_type ? T_1259 : T_1273;
  assign T_1277 = T_1274 == 1'h0;
  assign T_1278 = T_1277 | T_1211;
  assign T_1279 = T_1249 & T_1278;
  assign T_1305_manager_xact_id = io_grant_bits_payload_manager_xact_id;
  assign T_1341 = T_1247 == 1'h0;
  assign T_1342 = FinishQueue_16_1238_io_enq_ready | T_1341;
  assign T_1343 = T_1342 & io_grant_valid;
  assign T_1356 = T_1342 & io_refill_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  T_1203 = GEN_9[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1203 <= 3'h0;
    end else begin
      T_1203 <= GEN_0;
    end
  end
endmodule
module ClientUncachedTileLinkNetworkPort_14(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [25:0] io_client_acquire_bits_addr_block,
  input  [1:0] io_client_acquire_bits_client_xact_id,
  input  [2:0] io_client_acquire_bits_addr_beat,
  input   io_client_acquire_bits_is_builtin_type,
  input  [2:0] io_client_acquire_bits_a_type,
  input  [11:0] io_client_acquire_bits_union,
  input  [63:0] io_client_acquire_bits_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_addr_beat,
  output [1:0] io_client_grant_bits_client_xact_id,
  output [2:0] io_client_grant_bits_manager_xact_id,
  output  io_client_grant_bits_is_builtin_type,
  output [3:0] io_client_grant_bits_g_type,
  output [63:0] io_client_grant_bits_data,
  input   io_network_acquire_ready,
  output  io_network_acquire_valid,
  output [2:0] io_network_acquire_bits_header_src,
  output [2:0] io_network_acquire_bits_header_dst,
  output [25:0] io_network_acquire_bits_payload_addr_block,
  output [1:0] io_network_acquire_bits_payload_client_xact_id,
  output [2:0] io_network_acquire_bits_payload_addr_beat,
  output  io_network_acquire_bits_payload_is_builtin_type,
  output [2:0] io_network_acquire_bits_payload_a_type,
  output [11:0] io_network_acquire_bits_payload_union,
  output [63:0] io_network_acquire_bits_payload_data,
  output  io_network_grant_ready,
  input   io_network_grant_valid,
  input  [2:0] io_network_grant_bits_header_src,
  input  [2:0] io_network_grant_bits_header_dst,
  input  [2:0] io_network_grant_bits_payload_addr_beat,
  input  [1:0] io_network_grant_bits_payload_client_xact_id,
  input  [2:0] io_network_grant_bits_payload_manager_xact_id,
  input   io_network_grant_bits_payload_is_builtin_type,
  input  [3:0] io_network_grant_bits_payload_g_type,
  input  [63:0] io_network_grant_bits_payload_data,
  input   io_network_finish_ready,
  output  io_network_finish_valid,
  output [2:0] io_network_finish_bits_header_src,
  output [2:0] io_network_finish_bits_header_dst,
  output [2:0] io_network_finish_bits_payload_manager_xact_id,
  output  io_network_probe_ready,
  input   io_network_probe_valid,
  input  [2:0] io_network_probe_bits_header_src,
  input  [2:0] io_network_probe_bits_header_dst,
  input  [25:0] io_network_probe_bits_payload_addr_block,
  input  [1:0] io_network_probe_bits_payload_p_type,
  input   io_network_release_ready,
  output  io_network_release_valid,
  output [2:0] io_network_release_bits_header_src,
  output [2:0] io_network_release_bits_header_dst,
  output [2:0] io_network_release_bits_payload_addr_beat,
  output [25:0] io_network_release_bits_payload_addr_block,
  output [1:0] io_network_release_bits_payload_client_xact_id,
  output  io_network_release_bits_payload_voluntary,
  output [2:0] io_network_release_bits_payload_r_type,
  output [63:0] io_network_release_bits_payload_data
);
  wire  finisher_clk;
  wire  finisher_reset;
  wire  finisher_io_grant_ready;
  wire  finisher_io_grant_valid;
  wire [2:0] finisher_io_grant_bits_header_src;
  wire [2:0] finisher_io_grant_bits_header_dst;
  wire [2:0] finisher_io_grant_bits_payload_addr_beat;
  wire [1:0] finisher_io_grant_bits_payload_client_xact_id;
  wire [2:0] finisher_io_grant_bits_payload_manager_xact_id;
  wire  finisher_io_grant_bits_payload_is_builtin_type;
  wire [3:0] finisher_io_grant_bits_payload_g_type;
  wire [63:0] finisher_io_grant_bits_payload_data;
  wire  finisher_io_refill_ready;
  wire  finisher_io_refill_valid;
  wire [2:0] finisher_io_refill_bits_addr_beat;
  wire [1:0] finisher_io_refill_bits_client_xact_id;
  wire [2:0] finisher_io_refill_bits_manager_xact_id;
  wire  finisher_io_refill_bits_is_builtin_type;
  wire [3:0] finisher_io_refill_bits_g_type;
  wire [63:0] finisher_io_refill_bits_data;
  wire  finisher_io_finish_ready;
  wire  finisher_io_finish_valid;
  wire [2:0] finisher_io_finish_bits_header_src;
  wire [2:0] finisher_io_finish_bits_header_dst;
  wire [2:0] finisher_io_finish_bits_payload_manager_xact_id;
  wire  finisher_io_ready;
  wire  acq_with_header_ready;
  wire  acq_with_header_valid;
  wire [2:0] acq_with_header_bits_header_src;
  wire [2:0] acq_with_header_bits_header_dst;
  wire [25:0] acq_with_header_bits_payload_addr_block;
  wire [1:0] acq_with_header_bits_payload_client_xact_id;
  wire [2:0] acq_with_header_bits_payload_addr_beat;
  wire  acq_with_header_bits_payload_is_builtin_type;
  wire [2:0] acq_with_header_bits_payload_a_type;
  wire [11:0] acq_with_header_bits_payload_union;
  wire [63:0] acq_with_header_bits_payload_data;
  wire [31:0] GEN_0;
  wire [31:0] T_3765;
  wire  T_3767;
  wire  T_3773;
  wire  T_3774;
  wire  T_3775;
  reg [2:0] GEN_1;
  reg [31:0] GEN_9;
  reg [2:0] GEN_2;
  reg [31:0] GEN_10;
  reg [2:0] GEN_3;
  reg [31:0] GEN_11;
  reg [25:0] GEN_4;
  reg [31:0] GEN_12;
  reg [1:0] GEN_5;
  reg [31:0] GEN_13;
  reg  GEN_6;
  reg [31:0] GEN_14;
  reg [2:0] GEN_7;
  reg [31:0] GEN_15;
  reg [63:0] GEN_8;
  reg [63:0] GEN_16;
  FinishUnit_15 finisher (
    .clk(finisher_clk),
    .reset(finisher_reset),
    .io_grant_ready(finisher_io_grant_ready),
    .io_grant_valid(finisher_io_grant_valid),
    .io_grant_bits_header_src(finisher_io_grant_bits_header_src),
    .io_grant_bits_header_dst(finisher_io_grant_bits_header_dst),
    .io_grant_bits_payload_addr_beat(finisher_io_grant_bits_payload_addr_beat),
    .io_grant_bits_payload_client_xact_id(finisher_io_grant_bits_payload_client_xact_id),
    .io_grant_bits_payload_manager_xact_id(finisher_io_grant_bits_payload_manager_xact_id),
    .io_grant_bits_payload_is_builtin_type(finisher_io_grant_bits_payload_is_builtin_type),
    .io_grant_bits_payload_g_type(finisher_io_grant_bits_payload_g_type),
    .io_grant_bits_payload_data(finisher_io_grant_bits_payload_data),
    .io_refill_ready(finisher_io_refill_ready),
    .io_refill_valid(finisher_io_refill_valid),
    .io_refill_bits_addr_beat(finisher_io_refill_bits_addr_beat),
    .io_refill_bits_client_xact_id(finisher_io_refill_bits_client_xact_id),
    .io_refill_bits_manager_xact_id(finisher_io_refill_bits_manager_xact_id),
    .io_refill_bits_is_builtin_type(finisher_io_refill_bits_is_builtin_type),
    .io_refill_bits_g_type(finisher_io_refill_bits_g_type),
    .io_refill_bits_data(finisher_io_refill_bits_data),
    .io_finish_ready(finisher_io_finish_ready),
    .io_finish_valid(finisher_io_finish_valid),
    .io_finish_bits_header_src(finisher_io_finish_bits_header_src),
    .io_finish_bits_header_dst(finisher_io_finish_bits_header_dst),
    .io_finish_bits_payload_manager_xact_id(finisher_io_finish_bits_payload_manager_xact_id),
    .io_ready(finisher_io_ready)
  );
  assign io_client_acquire_ready = acq_with_header_ready;
  assign io_client_grant_valid = finisher_io_refill_valid;
  assign io_client_grant_bits_addr_beat = finisher_io_refill_bits_addr_beat;
  assign io_client_grant_bits_client_xact_id = finisher_io_refill_bits_client_xact_id;
  assign io_client_grant_bits_manager_xact_id = finisher_io_refill_bits_manager_xact_id;
  assign io_client_grant_bits_is_builtin_type = finisher_io_refill_bits_is_builtin_type;
  assign io_client_grant_bits_g_type = finisher_io_refill_bits_g_type;
  assign io_client_grant_bits_data = finisher_io_refill_bits_data;
  assign io_network_acquire_valid = T_3774;
  assign io_network_acquire_bits_header_src = acq_with_header_bits_header_src;
  assign io_network_acquire_bits_header_dst = acq_with_header_bits_header_dst;
  assign io_network_acquire_bits_payload_addr_block = acq_with_header_bits_payload_addr_block;
  assign io_network_acquire_bits_payload_client_xact_id = acq_with_header_bits_payload_client_xact_id;
  assign io_network_acquire_bits_payload_addr_beat = acq_with_header_bits_payload_addr_beat;
  assign io_network_acquire_bits_payload_is_builtin_type = acq_with_header_bits_payload_is_builtin_type;
  assign io_network_acquire_bits_payload_a_type = acq_with_header_bits_payload_a_type;
  assign io_network_acquire_bits_payload_union = acq_with_header_bits_payload_union;
  assign io_network_acquire_bits_payload_data = acq_with_header_bits_payload_data;
  assign io_network_grant_ready = finisher_io_grant_ready;
  assign io_network_finish_valid = finisher_io_finish_valid;
  assign io_network_finish_bits_header_src = finisher_io_finish_bits_header_src;
  assign io_network_finish_bits_header_dst = finisher_io_finish_bits_header_dst;
  assign io_network_finish_bits_payload_manager_xact_id = finisher_io_finish_bits_payload_manager_xact_id;
  assign io_network_probe_ready = 1'h0;
  assign io_network_release_valid = 1'h0;
  assign io_network_release_bits_header_src = GEN_1;
  assign io_network_release_bits_header_dst = GEN_2;
  assign io_network_release_bits_payload_addr_beat = GEN_3;
  assign io_network_release_bits_payload_addr_block = GEN_4;
  assign io_network_release_bits_payload_client_xact_id = GEN_5;
  assign io_network_release_bits_payload_voluntary = GEN_6;
  assign io_network_release_bits_payload_r_type = GEN_7;
  assign io_network_release_bits_payload_data = GEN_8;
  assign finisher_clk = clk;
  assign finisher_reset = reset;
  assign finisher_io_grant_valid = io_network_grant_valid;
  assign finisher_io_grant_bits_header_src = io_network_grant_bits_header_src;
  assign finisher_io_grant_bits_header_dst = io_network_grant_bits_header_dst;
  assign finisher_io_grant_bits_payload_addr_beat = io_network_grant_bits_payload_addr_beat;
  assign finisher_io_grant_bits_payload_client_xact_id = io_network_grant_bits_payload_client_xact_id;
  assign finisher_io_grant_bits_payload_manager_xact_id = io_network_grant_bits_payload_manager_xact_id;
  assign finisher_io_grant_bits_payload_is_builtin_type = io_network_grant_bits_payload_is_builtin_type;
  assign finisher_io_grant_bits_payload_g_type = io_network_grant_bits_payload_g_type;
  assign finisher_io_grant_bits_payload_data = io_network_grant_bits_payload_data;
  assign finisher_io_refill_ready = io_client_grant_ready;
  assign finisher_io_finish_ready = io_network_finish_ready;
  assign acq_with_header_ready = T_3775;
  assign acq_with_header_valid = io_client_acquire_valid;
  assign acq_with_header_bits_header_src = {{1'd0}, 2'h2};
  assign acq_with_header_bits_header_dst = {{2'd0}, T_3773};
  assign acq_with_header_bits_payload_addr_block = io_client_acquire_bits_addr_block;
  assign acq_with_header_bits_payload_client_xact_id = io_client_acquire_bits_client_xact_id;
  assign acq_with_header_bits_payload_addr_beat = io_client_acquire_bits_addr_beat;
  assign acq_with_header_bits_payload_is_builtin_type = io_client_acquire_bits_is_builtin_type;
  assign acq_with_header_bits_payload_a_type = io_client_acquire_bits_a_type;
  assign acq_with_header_bits_payload_union = io_client_acquire_bits_union;
  assign acq_with_header_bits_payload_data = io_client_acquire_bits_data;
  assign GEN_0 = {{6'd0}, io_client_acquire_bits_addr_block};
  assign T_3765 = GEN_0 << 6;
  assign T_3767 = 32'h80000000 <= T_3765;
  assign T_3773 = T_3767 ? 1'h0 : 1'h1;
  assign T_3774 = acq_with_header_valid & finisher_io_ready;
  assign T_3775 = io_network_acquire_ready & finisher_io_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  GEN_1 = GEN_9[2:0];
  GEN_10 = {1{$random}};
  GEN_2 = GEN_10[2:0];
  GEN_11 = {1{$random}};
  GEN_3 = GEN_11[2:0];
  GEN_12 = {1{$random}};
  GEN_4 = GEN_12[25:0];
  GEN_13 = {1{$random}};
  GEN_5 = GEN_13[1:0];
  GEN_14 = {1{$random}};
  GEN_6 = GEN_14[0:0];
  GEN_15 = {1{$random}};
  GEN_7 = GEN_15[2:0];
  GEN_16 = {2{$random}};
  GEN_8 = GEN_16[63:0];
  end
`endif
endmodule
module ManagerTileLinkNetworkPort(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output [1:0] io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input  [1:0] io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input  [1:0] io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output [1:0] io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [2:0] io_network_acquire_bits_header_src,
  input  [2:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [2:0] io_network_grant_bits_header_src,
  output [2:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [2:0] io_network_finish_bits_header_src,
  input  [2:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [2:0] io_network_probe_bits_header_src,
  output [2:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [2:0] io_network_release_bits_header_src,
  input  [2:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6829_ready;
  wire  T_6829_valid;
  wire [2:0] T_6829_bits_header_src;
  wire [2:0] T_6829_bits_header_dst;
  wire [2:0] T_6829_bits_payload_addr_beat;
  wire [1:0] T_6829_bits_payload_client_xact_id;
  wire [2:0] T_6829_bits_payload_manager_xact_id;
  wire  T_6829_bits_payload_is_builtin_type;
  wire [3:0] T_6829_bits_payload_g_type;
  wire [63:0] T_6829_bits_payload_data;
  wire [1:0] T_6829_bits_payload_client_id;
  wire  T_7459_ready;
  wire  T_7459_valid;
  wire [2:0] T_7459_bits_header_src;
  wire [2:0] T_7459_bits_header_dst;
  wire [25:0] T_7459_bits_payload_addr_block;
  wire [1:0] T_7459_bits_payload_p_type;
  wire [1:0] T_7459_bits_payload_client_id;
  wire  T_7774_ready;
  wire  T_7774_valid;
  wire [25:0] T_7774_bits_addr_block;
  wire [1:0] T_7774_bits_client_xact_id;
  wire [2:0] T_7774_bits_addr_beat;
  wire  T_7774_bits_is_builtin_type;
  wire [2:0] T_7774_bits_a_type;
  wire [11:0] T_7774_bits_union;
  wire [63:0] T_7774_bits_data;
  wire  T_7902_ready;
  wire  T_7902_valid;
  wire [2:0] T_7902_bits_addr_beat;
  wire [25:0] T_7902_bits_addr_block;
  wire [1:0] T_7902_bits_client_xact_id;
  wire  T_7902_bits_voluntary;
  wire [2:0] T_7902_bits_r_type;
  wire [63:0] T_7902_bits_data;
  wire  T_8018_ready;
  wire  T_8018_valid;
  wire [2:0] T_8018_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_7774_valid;
  assign io_manager_acquire_bits_addr_block = T_7774_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_7774_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_7774_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_7774_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_7774_bits_a_type;
  assign io_manager_acquire_bits_union = T_7774_bits_union;
  assign io_manager_acquire_bits_data = T_7774_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[1:0];
  assign io_manager_grant_ready = T_6829_ready;
  assign io_manager_finish_valid = T_8018_valid;
  assign io_manager_finish_bits_manager_xact_id = T_8018_bits_manager_xact_id;
  assign io_manager_probe_ready = T_7459_ready;
  assign io_manager_release_valid = T_7902_valid;
  assign io_manager_release_bits_addr_beat = T_7902_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_7902_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_7902_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_7902_bits_voluntary;
  assign io_manager_release_bits_r_type = T_7902_bits_r_type;
  assign io_manager_release_bits_data = T_7902_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[1:0];
  assign io_network_acquire_ready = T_7774_ready;
  assign io_network_grant_valid = T_6829_valid;
  assign io_network_grant_bits_header_src = T_6829_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6829_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6829_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6829_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6829_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6829_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6829_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6829_bits_payload_data;
  assign io_network_finish_ready = T_8018_ready;
  assign io_network_probe_valid = T_7459_valid;
  assign io_network_probe_bits_header_src = T_7459_bits_header_src;
  assign io_network_probe_bits_header_dst = T_7459_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_7459_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_7459_bits_payload_p_type;
  assign io_network_release_ready = T_7902_ready;
  assign T_6829_ready = io_network_grant_ready;
  assign T_6829_valid = io_manager_grant_valid;
  assign T_6829_bits_header_src = {{2'd0}, 1'h0};
  assign T_6829_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6829_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6829_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6829_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6829_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6829_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6829_bits_payload_data = io_manager_grant_bits_data;
  assign T_6829_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_7459_ready = io_network_probe_ready;
  assign T_7459_valid = io_manager_probe_valid;
  assign T_7459_bits_header_src = {{2'd0}, 1'h0};
  assign T_7459_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_7459_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_7459_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_7459_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_7774_ready = io_manager_acquire_ready;
  assign T_7774_valid = io_network_acquire_valid;
  assign T_7774_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_7774_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_7774_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_7774_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_7774_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_7774_bits_union = io_network_acquire_bits_payload_union;
  assign T_7774_bits_data = io_network_acquire_bits_payload_data;
  assign T_7902_ready = io_manager_release_ready;
  assign T_7902_valid = io_network_release_valid;
  assign T_7902_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_7902_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_7902_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_7902_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_7902_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_7902_bits_data = io_network_release_bits_payload_data;
  assign T_8018_ready = io_manager_finish_ready;
  assign T_8018_valid = io_network_finish_valid;
  assign T_8018_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module TileLinkEnqueuer_17(
  input   clk,
  input   reset,
  output  io_client_acquire_ready,
  input   io_client_acquire_valid,
  input  [2:0] io_client_acquire_bits_header_src,
  input  [2:0] io_client_acquire_bits_header_dst,
  input  [25:0] io_client_acquire_bits_payload_addr_block,
  input  [1:0] io_client_acquire_bits_payload_client_xact_id,
  input  [2:0] io_client_acquire_bits_payload_addr_beat,
  input   io_client_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_client_acquire_bits_payload_a_type,
  input  [11:0] io_client_acquire_bits_payload_union,
  input  [63:0] io_client_acquire_bits_payload_data,
  input   io_client_grant_ready,
  output  io_client_grant_valid,
  output [2:0] io_client_grant_bits_header_src,
  output [2:0] io_client_grant_bits_header_dst,
  output [2:0] io_client_grant_bits_payload_addr_beat,
  output [1:0] io_client_grant_bits_payload_client_xact_id,
  output [2:0] io_client_grant_bits_payload_manager_xact_id,
  output  io_client_grant_bits_payload_is_builtin_type,
  output [3:0] io_client_grant_bits_payload_g_type,
  output [63:0] io_client_grant_bits_payload_data,
  output  io_client_finish_ready,
  input   io_client_finish_valid,
  input  [2:0] io_client_finish_bits_header_src,
  input  [2:0] io_client_finish_bits_header_dst,
  input  [2:0] io_client_finish_bits_payload_manager_xact_id,
  input   io_client_probe_ready,
  output  io_client_probe_valid,
  output [2:0] io_client_probe_bits_header_src,
  output [2:0] io_client_probe_bits_header_dst,
  output [25:0] io_client_probe_bits_payload_addr_block,
  output [1:0] io_client_probe_bits_payload_p_type,
  output  io_client_release_ready,
  input   io_client_release_valid,
  input  [2:0] io_client_release_bits_header_src,
  input  [2:0] io_client_release_bits_header_dst,
  input  [2:0] io_client_release_bits_payload_addr_beat,
  input  [25:0] io_client_release_bits_payload_addr_block,
  input  [1:0] io_client_release_bits_payload_client_xact_id,
  input   io_client_release_bits_payload_voluntary,
  input  [2:0] io_client_release_bits_payload_r_type,
  input  [63:0] io_client_release_bits_payload_data,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [2:0] io_manager_acquire_bits_header_src,
  output [2:0] io_manager_acquire_bits_header_dst,
  output [25:0] io_manager_acquire_bits_payload_addr_block,
  output [1:0] io_manager_acquire_bits_payload_client_xact_id,
  output [2:0] io_manager_acquire_bits_payload_addr_beat,
  output  io_manager_acquire_bits_payload_is_builtin_type,
  output [2:0] io_manager_acquire_bits_payload_a_type,
  output [11:0] io_manager_acquire_bits_payload_union,
  output [63:0] io_manager_acquire_bits_payload_data,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_header_src,
  input  [2:0] io_manager_grant_bits_header_dst,
  input  [2:0] io_manager_grant_bits_payload_addr_beat,
  input  [1:0] io_manager_grant_bits_payload_client_xact_id,
  input  [2:0] io_manager_grant_bits_payload_manager_xact_id,
  input   io_manager_grant_bits_payload_is_builtin_type,
  input  [3:0] io_manager_grant_bits_payload_g_type,
  input  [63:0] io_manager_grant_bits_payload_data,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_header_src,
  output [2:0] io_manager_finish_bits_header_dst,
  output [2:0] io_manager_finish_bits_payload_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [2:0] io_manager_probe_bits_header_src,
  input  [2:0] io_manager_probe_bits_header_dst,
  input  [25:0] io_manager_probe_bits_payload_addr_block,
  input  [1:0] io_manager_probe_bits_payload_p_type,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_header_src,
  output [2:0] io_manager_release_bits_header_dst,
  output [2:0] io_manager_release_bits_payload_addr_beat,
  output [25:0] io_manager_release_bits_payload_addr_block,
  output [1:0] io_manager_release_bits_payload_client_xact_id,
  output  io_manager_release_bits_payload_voluntary,
  output [2:0] io_manager_release_bits_payload_r_type,
  output [63:0] io_manager_release_bits_payload_data
);
  assign io_client_acquire_ready = io_manager_acquire_ready;
  assign io_client_grant_valid = io_manager_grant_valid;
  assign io_client_grant_bits_header_src = io_manager_grant_bits_header_src;
  assign io_client_grant_bits_header_dst = io_manager_grant_bits_header_dst;
  assign io_client_grant_bits_payload_addr_beat = io_manager_grant_bits_payload_addr_beat;
  assign io_client_grant_bits_payload_client_xact_id = io_manager_grant_bits_payload_client_xact_id;
  assign io_client_grant_bits_payload_manager_xact_id = io_manager_grant_bits_payload_manager_xact_id;
  assign io_client_grant_bits_payload_is_builtin_type = io_manager_grant_bits_payload_is_builtin_type;
  assign io_client_grant_bits_payload_g_type = io_manager_grant_bits_payload_g_type;
  assign io_client_grant_bits_payload_data = io_manager_grant_bits_payload_data;
  assign io_client_finish_ready = io_manager_finish_ready;
  assign io_client_probe_valid = io_manager_probe_valid;
  assign io_client_probe_bits_header_src = io_manager_probe_bits_header_src;
  assign io_client_probe_bits_header_dst = io_manager_probe_bits_header_dst;
  assign io_client_probe_bits_payload_addr_block = io_manager_probe_bits_payload_addr_block;
  assign io_client_probe_bits_payload_p_type = io_manager_probe_bits_payload_p_type;
  assign io_client_release_ready = io_manager_release_ready;
  assign io_manager_acquire_valid = io_client_acquire_valid;
  assign io_manager_acquire_bits_header_src = io_client_acquire_bits_header_src;
  assign io_manager_acquire_bits_header_dst = io_client_acquire_bits_header_dst;
  assign io_manager_acquire_bits_payload_addr_block = io_client_acquire_bits_payload_addr_block;
  assign io_manager_acquire_bits_payload_client_xact_id = io_client_acquire_bits_payload_client_xact_id;
  assign io_manager_acquire_bits_payload_addr_beat = io_client_acquire_bits_payload_addr_beat;
  assign io_manager_acquire_bits_payload_is_builtin_type = io_client_acquire_bits_payload_is_builtin_type;
  assign io_manager_acquire_bits_payload_a_type = io_client_acquire_bits_payload_a_type;
  assign io_manager_acquire_bits_payload_union = io_client_acquire_bits_payload_union;
  assign io_manager_acquire_bits_payload_data = io_client_acquire_bits_payload_data;
  assign io_manager_grant_ready = io_client_grant_ready;
  assign io_manager_finish_valid = io_client_finish_valid;
  assign io_manager_finish_bits_header_src = io_client_finish_bits_header_src;
  assign io_manager_finish_bits_header_dst = io_client_finish_bits_header_dst;
  assign io_manager_finish_bits_payload_manager_xact_id = io_client_finish_bits_payload_manager_xact_id;
  assign io_manager_probe_ready = io_client_probe_ready;
  assign io_manager_release_valid = io_client_release_valid;
  assign io_manager_release_bits_header_src = io_client_release_bits_header_src;
  assign io_manager_release_bits_header_dst = io_client_release_bits_header_dst;
  assign io_manager_release_bits_payload_addr_beat = io_client_release_bits_payload_addr_beat;
  assign io_manager_release_bits_payload_addr_block = io_client_release_bits_payload_addr_block;
  assign io_manager_release_bits_payload_client_xact_id = io_client_release_bits_payload_client_xact_id;
  assign io_manager_release_bits_payload_voluntary = io_client_release_bits_payload_voluntary;
  assign io_manager_release_bits_payload_r_type = io_client_release_bits_payload_r_type;
  assign io_manager_release_bits_payload_data = io_client_release_bits_payload_data;
endmodule
module ManagerTileLinkNetworkPort_18(
  input   clk,
  input   reset,
  input   io_manager_acquire_ready,
  output  io_manager_acquire_valid,
  output [25:0] io_manager_acquire_bits_addr_block,
  output [1:0] io_manager_acquire_bits_client_xact_id,
  output [2:0] io_manager_acquire_bits_addr_beat,
  output  io_manager_acquire_bits_is_builtin_type,
  output [2:0] io_manager_acquire_bits_a_type,
  output [11:0] io_manager_acquire_bits_union,
  output [63:0] io_manager_acquire_bits_data,
  output [1:0] io_manager_acquire_bits_client_id,
  output  io_manager_grant_ready,
  input   io_manager_grant_valid,
  input  [2:0] io_manager_grant_bits_addr_beat,
  input  [1:0] io_manager_grant_bits_client_xact_id,
  input  [2:0] io_manager_grant_bits_manager_xact_id,
  input   io_manager_grant_bits_is_builtin_type,
  input  [3:0] io_manager_grant_bits_g_type,
  input  [63:0] io_manager_grant_bits_data,
  input  [1:0] io_manager_grant_bits_client_id,
  input   io_manager_finish_ready,
  output  io_manager_finish_valid,
  output [2:0] io_manager_finish_bits_manager_xact_id,
  output  io_manager_probe_ready,
  input   io_manager_probe_valid,
  input  [25:0] io_manager_probe_bits_addr_block,
  input  [1:0] io_manager_probe_bits_p_type,
  input  [1:0] io_manager_probe_bits_client_id,
  input   io_manager_release_ready,
  output  io_manager_release_valid,
  output [2:0] io_manager_release_bits_addr_beat,
  output [25:0] io_manager_release_bits_addr_block,
  output [1:0] io_manager_release_bits_client_xact_id,
  output  io_manager_release_bits_voluntary,
  output [2:0] io_manager_release_bits_r_type,
  output [63:0] io_manager_release_bits_data,
  output [1:0] io_manager_release_bits_client_id,
  output  io_network_acquire_ready,
  input   io_network_acquire_valid,
  input  [2:0] io_network_acquire_bits_header_src,
  input  [2:0] io_network_acquire_bits_header_dst,
  input  [25:0] io_network_acquire_bits_payload_addr_block,
  input  [1:0] io_network_acquire_bits_payload_client_xact_id,
  input  [2:0] io_network_acquire_bits_payload_addr_beat,
  input   io_network_acquire_bits_payload_is_builtin_type,
  input  [2:0] io_network_acquire_bits_payload_a_type,
  input  [11:0] io_network_acquire_bits_payload_union,
  input  [63:0] io_network_acquire_bits_payload_data,
  input   io_network_grant_ready,
  output  io_network_grant_valid,
  output [2:0] io_network_grant_bits_header_src,
  output [2:0] io_network_grant_bits_header_dst,
  output [2:0] io_network_grant_bits_payload_addr_beat,
  output [1:0] io_network_grant_bits_payload_client_xact_id,
  output [2:0] io_network_grant_bits_payload_manager_xact_id,
  output  io_network_grant_bits_payload_is_builtin_type,
  output [3:0] io_network_grant_bits_payload_g_type,
  output [63:0] io_network_grant_bits_payload_data,
  output  io_network_finish_ready,
  input   io_network_finish_valid,
  input  [2:0] io_network_finish_bits_header_src,
  input  [2:0] io_network_finish_bits_header_dst,
  input  [2:0] io_network_finish_bits_payload_manager_xact_id,
  input   io_network_probe_ready,
  output  io_network_probe_valid,
  output [2:0] io_network_probe_bits_header_src,
  output [2:0] io_network_probe_bits_header_dst,
  output [25:0] io_network_probe_bits_payload_addr_block,
  output [1:0] io_network_probe_bits_payload_p_type,
  output  io_network_release_ready,
  input   io_network_release_valid,
  input  [2:0] io_network_release_bits_header_src,
  input  [2:0] io_network_release_bits_header_dst,
  input  [2:0] io_network_release_bits_payload_addr_beat,
  input  [25:0] io_network_release_bits_payload_addr_block,
  input  [1:0] io_network_release_bits_payload_client_xact_id,
  input   io_network_release_bits_payload_voluntary,
  input  [2:0] io_network_release_bits_payload_r_type,
  input  [63:0] io_network_release_bits_payload_data
);
  wire  T_6829_ready;
  wire  T_6829_valid;
  wire [2:0] T_6829_bits_header_src;
  wire [2:0] T_6829_bits_header_dst;
  wire [2:0] T_6829_bits_payload_addr_beat;
  wire [1:0] T_6829_bits_payload_client_xact_id;
  wire [2:0] T_6829_bits_payload_manager_xact_id;
  wire  T_6829_bits_payload_is_builtin_type;
  wire [3:0] T_6829_bits_payload_g_type;
  wire [63:0] T_6829_bits_payload_data;
  wire [1:0] T_6829_bits_payload_client_id;
  wire  T_7459_ready;
  wire  T_7459_valid;
  wire [2:0] T_7459_bits_header_src;
  wire [2:0] T_7459_bits_header_dst;
  wire [25:0] T_7459_bits_payload_addr_block;
  wire [1:0] T_7459_bits_payload_p_type;
  wire [1:0] T_7459_bits_payload_client_id;
  wire  T_7774_ready;
  wire  T_7774_valid;
  wire [25:0] T_7774_bits_addr_block;
  wire [1:0] T_7774_bits_client_xact_id;
  wire [2:0] T_7774_bits_addr_beat;
  wire  T_7774_bits_is_builtin_type;
  wire [2:0] T_7774_bits_a_type;
  wire [11:0] T_7774_bits_union;
  wire [63:0] T_7774_bits_data;
  wire  T_7902_ready;
  wire  T_7902_valid;
  wire [2:0] T_7902_bits_addr_beat;
  wire [25:0] T_7902_bits_addr_block;
  wire [1:0] T_7902_bits_client_xact_id;
  wire  T_7902_bits_voluntary;
  wire [2:0] T_7902_bits_r_type;
  wire [63:0] T_7902_bits_data;
  wire  T_8018_ready;
  wire  T_8018_valid;
  wire [2:0] T_8018_bits_manager_xact_id;
  assign io_manager_acquire_valid = T_7774_valid;
  assign io_manager_acquire_bits_addr_block = T_7774_bits_addr_block;
  assign io_manager_acquire_bits_client_xact_id = T_7774_bits_client_xact_id;
  assign io_manager_acquire_bits_addr_beat = T_7774_bits_addr_beat;
  assign io_manager_acquire_bits_is_builtin_type = T_7774_bits_is_builtin_type;
  assign io_manager_acquire_bits_a_type = T_7774_bits_a_type;
  assign io_manager_acquire_bits_union = T_7774_bits_union;
  assign io_manager_acquire_bits_data = T_7774_bits_data;
  assign io_manager_acquire_bits_client_id = io_network_acquire_bits_header_src[1:0];
  assign io_manager_grant_ready = T_6829_ready;
  assign io_manager_finish_valid = T_8018_valid;
  assign io_manager_finish_bits_manager_xact_id = T_8018_bits_manager_xact_id;
  assign io_manager_probe_ready = T_7459_ready;
  assign io_manager_release_valid = T_7902_valid;
  assign io_manager_release_bits_addr_beat = T_7902_bits_addr_beat;
  assign io_manager_release_bits_addr_block = T_7902_bits_addr_block;
  assign io_manager_release_bits_client_xact_id = T_7902_bits_client_xact_id;
  assign io_manager_release_bits_voluntary = T_7902_bits_voluntary;
  assign io_manager_release_bits_r_type = T_7902_bits_r_type;
  assign io_manager_release_bits_data = T_7902_bits_data;
  assign io_manager_release_bits_client_id = io_network_release_bits_header_src[1:0];
  assign io_network_acquire_ready = T_7774_ready;
  assign io_network_grant_valid = T_6829_valid;
  assign io_network_grant_bits_header_src = T_6829_bits_header_src;
  assign io_network_grant_bits_header_dst = T_6829_bits_header_dst;
  assign io_network_grant_bits_payload_addr_beat = T_6829_bits_payload_addr_beat;
  assign io_network_grant_bits_payload_client_xact_id = T_6829_bits_payload_client_xact_id;
  assign io_network_grant_bits_payload_manager_xact_id = T_6829_bits_payload_manager_xact_id;
  assign io_network_grant_bits_payload_is_builtin_type = T_6829_bits_payload_is_builtin_type;
  assign io_network_grant_bits_payload_g_type = T_6829_bits_payload_g_type;
  assign io_network_grant_bits_payload_data = T_6829_bits_payload_data;
  assign io_network_finish_ready = T_8018_ready;
  assign io_network_probe_valid = T_7459_valid;
  assign io_network_probe_bits_header_src = T_7459_bits_header_src;
  assign io_network_probe_bits_header_dst = T_7459_bits_header_dst;
  assign io_network_probe_bits_payload_addr_block = T_7459_bits_payload_addr_block;
  assign io_network_probe_bits_payload_p_type = T_7459_bits_payload_p_type;
  assign io_network_release_ready = T_7902_ready;
  assign T_6829_ready = io_network_grant_ready;
  assign T_6829_valid = io_manager_grant_valid;
  assign T_6829_bits_header_src = {{2'd0}, 1'h1};
  assign T_6829_bits_header_dst = {{1'd0}, io_manager_grant_bits_client_id};
  assign T_6829_bits_payload_addr_beat = io_manager_grant_bits_addr_beat;
  assign T_6829_bits_payload_client_xact_id = io_manager_grant_bits_client_xact_id;
  assign T_6829_bits_payload_manager_xact_id = io_manager_grant_bits_manager_xact_id;
  assign T_6829_bits_payload_is_builtin_type = io_manager_grant_bits_is_builtin_type;
  assign T_6829_bits_payload_g_type = io_manager_grant_bits_g_type;
  assign T_6829_bits_payload_data = io_manager_grant_bits_data;
  assign T_6829_bits_payload_client_id = io_manager_grant_bits_client_id;
  assign T_7459_ready = io_network_probe_ready;
  assign T_7459_valid = io_manager_probe_valid;
  assign T_7459_bits_header_src = {{2'd0}, 1'h1};
  assign T_7459_bits_header_dst = {{1'd0}, io_manager_probe_bits_client_id};
  assign T_7459_bits_payload_addr_block = io_manager_probe_bits_addr_block;
  assign T_7459_bits_payload_p_type = io_manager_probe_bits_p_type;
  assign T_7459_bits_payload_client_id = io_manager_probe_bits_client_id;
  assign T_7774_ready = io_manager_acquire_ready;
  assign T_7774_valid = io_network_acquire_valid;
  assign T_7774_bits_addr_block = io_network_acquire_bits_payload_addr_block;
  assign T_7774_bits_client_xact_id = io_network_acquire_bits_payload_client_xact_id;
  assign T_7774_bits_addr_beat = io_network_acquire_bits_payload_addr_beat;
  assign T_7774_bits_is_builtin_type = io_network_acquire_bits_payload_is_builtin_type;
  assign T_7774_bits_a_type = io_network_acquire_bits_payload_a_type;
  assign T_7774_bits_union = io_network_acquire_bits_payload_union;
  assign T_7774_bits_data = io_network_acquire_bits_payload_data;
  assign T_7902_ready = io_manager_release_ready;
  assign T_7902_valid = io_network_release_valid;
  assign T_7902_bits_addr_beat = io_network_release_bits_payload_addr_beat;
  assign T_7902_bits_addr_block = io_network_release_bits_payload_addr_block;
  assign T_7902_bits_client_xact_id = io_network_release_bits_payload_client_xact_id;
  assign T_7902_bits_voluntary = io_network_release_bits_payload_voluntary;
  assign T_7902_bits_r_type = io_network_release_bits_payload_r_type;
  assign T_7902_bits_data = io_network_release_bits_payload_data;
  assign T_8018_ready = io_manager_finish_ready;
  assign T_8018_valid = io_network_finish_valid;
  assign T_8018_bits_manager_xact_id = io_network_finish_bits_payload_manager_xact_id;
endmodule
module LockingRRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input   io_in_4_bits_payload_is_builtin_type,
  input  [2:0] io_in_4_bits_payload_a_type,
  input  [11:0] io_in_4_bits_payload_union,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_header_src,
  output [2:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_addr_beat,
  output  io_out_bits_payload_is_builtin_type,
  output [2:0] io_out_bits_payload_a_type,
  output [11:0] io_out_bits_payload_union,
  output [63:0] io_out_bits_payload_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_62;
  wire  GEN_10;
  wire [2:0] GEN_63;
  wire  GEN_11;
  wire [2:0] GEN_64;
  wire  GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_1;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [2:0] GEN_16;
  wire [2:0] GEN_17;
  wire [2:0] GEN_2;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [25:0] GEN_3;
  wire [25:0] GEN_22;
  wire [25:0] GEN_23;
  wire [25:0] GEN_24;
  wire [25:0] GEN_25;
  wire [1:0] GEN_4;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [2:0] GEN_5;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [2:0] GEN_33;
  wire  GEN_6;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire [2:0] GEN_7;
  wire [2:0] GEN_38;
  wire [2:0] GEN_39;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [11:0] GEN_8;
  wire [11:0] GEN_42;
  wire [11:0] GEN_43;
  wire [11:0] GEN_44;
  wire [11:0] GEN_45;
  wire [63:0] GEN_9;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  reg [2:0] T_1380;
  reg [31:0] GEN_65;
  reg [2:0] T_1382;
  reg [31:0] GEN_66;
  wire [2:0] GEN_92;
  wire  T_1384;
  wire [2:0] T_1393_0;
  wire  T_1395;
  wire  T_1398;
  wire  T_1399;
  wire  T_1400;
  wire [3:0] T_1404;
  wire [2:0] T_1405;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  wire [2:0] GEN_52;
  reg [2:0] lastGrant;
  reg [31:0] GEN_67;
  wire [2:0] GEN_53;
  wire  T_1410;
  wire  T_1412;
  wire  T_1414;
  wire  T_1416;
  wire  T_1418;
  wire  T_1419;
  wire  T_1420;
  wire  T_1421;
  wire  T_1424;
  wire  T_1425;
  wire  T_1426;
  wire  T_1427;
  wire  T_1428;
  wire  T_1429;
  wire  T_1430;
  wire  T_1434;
  wire  T_1436;
  wire  T_1438;
  wire  T_1440;
  wire  T_1442;
  wire  T_1444;
  wire  T_1446;
  wire  T_1448;
  wire  T_1452;
  wire  T_1453;
  wire  T_1454;
  wire  T_1455;
  wire  T_1456;
  wire  T_1457;
  wire  T_1458;
  wire  T_1460;
  wire  T_1461;
  wire  T_1462;
  wire  T_1464;
  wire  T_1465;
  wire  T_1466;
  wire  T_1468;
  wire  T_1469;
  wire  T_1470;
  wire  T_1472;
  wire  T_1473;
  wire  T_1474;
  wire  T_1476;
  wire  T_1477;
  wire  T_1478;
  wire [2:0] GEN_54;
  wire [2:0] GEN_55;
  wire [2:0] GEN_56;
  wire [2:0] GEN_57;
  wire [2:0] GEN_58;
  wire [2:0] GEN_59;
  wire [2:0] GEN_60;
  wire [2:0] GEN_61;
  assign io_in_0_ready = T_1462;
  assign io_in_1_ready = T_1466;
  assign io_in_2_ready = T_1470;
  assign io_in_3_ready = T_1474;
  assign io_in_4_ready = T_1478;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_addr_beat = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_a_type = GEN_7;
  assign io_out_bits_payload_union = GEN_8;
  assign io_out_bits_payload_data = GEN_9;
  assign io_chosen = GEN_52;
  assign choice = GEN_61;
  assign GEN_0 = GEN_13;
  assign GEN_62 = {{2'd0}, 1'h1};
  assign GEN_10 = GEN_62 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_63 = {{1'd0}, 2'h2};
  assign GEN_11 = GEN_63 == io_chosen ? io_in_2_valid : GEN_10;
  assign GEN_64 = {{1'd0}, 2'h3};
  assign GEN_12 = GEN_64 == io_chosen ? io_in_3_valid : GEN_11;
  assign GEN_13 = 3'h4 == io_chosen ? io_in_4_valid : GEN_12;
  assign GEN_1 = GEN_17;
  assign GEN_14 = GEN_62 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_15 = GEN_63 == io_chosen ? io_in_2_bits_header_src : GEN_14;
  assign GEN_16 = GEN_64 == io_chosen ? io_in_3_bits_header_src : GEN_15;
  assign GEN_17 = 3'h4 == io_chosen ? io_in_4_bits_header_src : GEN_16;
  assign GEN_2 = GEN_21;
  assign GEN_18 = GEN_62 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_19 = GEN_63 == io_chosen ? io_in_2_bits_header_dst : GEN_18;
  assign GEN_20 = GEN_64 == io_chosen ? io_in_3_bits_header_dst : GEN_19;
  assign GEN_21 = 3'h4 == io_chosen ? io_in_4_bits_header_dst : GEN_20;
  assign GEN_3 = GEN_25;
  assign GEN_22 = GEN_62 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_23 = GEN_63 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_22;
  assign GEN_24 = GEN_64 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_23;
  assign GEN_25 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_block : GEN_24;
  assign GEN_4 = GEN_29;
  assign GEN_26 = GEN_62 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_27 = GEN_63 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_26;
  assign GEN_28 = GEN_64 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_27;
  assign GEN_29 = 3'h4 == io_chosen ? io_in_4_bits_payload_client_xact_id : GEN_28;
  assign GEN_5 = GEN_33;
  assign GEN_30 = GEN_62 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_31 = GEN_63 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_30;
  assign GEN_32 = GEN_64 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_31;
  assign GEN_33 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_beat : GEN_32;
  assign GEN_6 = GEN_37;
  assign GEN_34 = GEN_62 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_35 = GEN_63 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_34;
  assign GEN_36 = GEN_64 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_35;
  assign GEN_37 = 3'h4 == io_chosen ? io_in_4_bits_payload_is_builtin_type : GEN_36;
  assign GEN_7 = GEN_41;
  assign GEN_38 = GEN_62 == io_chosen ? io_in_1_bits_payload_a_type : io_in_0_bits_payload_a_type;
  assign GEN_39 = GEN_63 == io_chosen ? io_in_2_bits_payload_a_type : GEN_38;
  assign GEN_40 = GEN_64 == io_chosen ? io_in_3_bits_payload_a_type : GEN_39;
  assign GEN_41 = 3'h4 == io_chosen ? io_in_4_bits_payload_a_type : GEN_40;
  assign GEN_8 = GEN_45;
  assign GEN_42 = GEN_62 == io_chosen ? io_in_1_bits_payload_union : io_in_0_bits_payload_union;
  assign GEN_43 = GEN_63 == io_chosen ? io_in_2_bits_payload_union : GEN_42;
  assign GEN_44 = GEN_64 == io_chosen ? io_in_3_bits_payload_union : GEN_43;
  assign GEN_45 = 3'h4 == io_chosen ? io_in_4_bits_payload_union : GEN_44;
  assign GEN_9 = GEN_49;
  assign GEN_46 = GEN_62 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_47 = GEN_63 == io_chosen ? io_in_2_bits_payload_data : GEN_46;
  assign GEN_48 = GEN_64 == io_chosen ? io_in_3_bits_payload_data : GEN_47;
  assign GEN_49 = 3'h4 == io_chosen ? io_in_4_bits_payload_data : GEN_48;
  assign GEN_92 = {{2'd0}, 1'h0};
  assign T_1384 = T_1380 != GEN_92;
  assign T_1393_0 = 3'h3;
  assign T_1395 = T_1393_0 == io_out_bits_payload_a_type;
  assign T_1398 = io_out_bits_payload_is_builtin_type & T_1395;
  assign T_1399 = io_out_ready & io_out_valid;
  assign T_1400 = T_1399 & T_1398;
  assign T_1404 = T_1380 + GEN_62;
  assign T_1405 = T_1404[2:0];
  assign GEN_50 = T_1400 ? io_chosen : T_1382;
  assign GEN_51 = T_1400 ? T_1405 : T_1380;
  assign GEN_52 = T_1384 ? T_1382 : choice;
  assign GEN_53 = T_1399 ? io_chosen : lastGrant;
  assign T_1410 = GEN_62 > lastGrant;
  assign T_1412 = GEN_63 > lastGrant;
  assign T_1414 = GEN_64 > lastGrant;
  assign T_1416 = 3'h4 > lastGrant;
  assign T_1418 = io_in_1_valid & T_1410;
  assign T_1419 = io_in_2_valid & T_1412;
  assign T_1420 = io_in_3_valid & T_1414;
  assign T_1421 = io_in_4_valid & T_1416;
  assign T_1424 = T_1418 | T_1419;
  assign T_1425 = T_1424 | T_1420;
  assign T_1426 = T_1425 | T_1421;
  assign T_1427 = T_1426 | io_in_0_valid;
  assign T_1428 = T_1427 | io_in_1_valid;
  assign T_1429 = T_1428 | io_in_2_valid;
  assign T_1430 = T_1429 | io_in_3_valid;
  assign T_1434 = T_1418 == 1'h0;
  assign T_1436 = T_1424 == 1'h0;
  assign T_1438 = T_1425 == 1'h0;
  assign T_1440 = T_1426 == 1'h0;
  assign T_1442 = T_1427 == 1'h0;
  assign T_1444 = T_1428 == 1'h0;
  assign T_1446 = T_1429 == 1'h0;
  assign T_1448 = T_1430 == 1'h0;
  assign T_1452 = T_1410 | T_1442;
  assign T_1453 = T_1434 & T_1412;
  assign T_1454 = T_1453 | T_1444;
  assign T_1455 = T_1436 & T_1414;
  assign T_1456 = T_1455 | T_1446;
  assign T_1457 = T_1438 & T_1416;
  assign T_1458 = T_1457 | T_1448;
  assign T_1460 = T_1382 == GEN_92;
  assign T_1461 = T_1384 ? T_1460 : T_1440;
  assign T_1462 = T_1461 & io_out_ready;
  assign T_1464 = T_1382 == GEN_62;
  assign T_1465 = T_1384 ? T_1464 : T_1452;
  assign T_1466 = T_1465 & io_out_ready;
  assign T_1468 = T_1382 == GEN_63;
  assign T_1469 = T_1384 ? T_1468 : T_1454;
  assign T_1470 = T_1469 & io_out_ready;
  assign T_1472 = T_1382 == GEN_64;
  assign T_1473 = T_1384 ? T_1472 : T_1456;
  assign T_1474 = T_1473 & io_out_ready;
  assign T_1476 = T_1382 == 3'h4;
  assign T_1477 = T_1384 ? T_1476 : T_1458;
  assign T_1478 = T_1477 & io_out_ready;
  assign GEN_54 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_55 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_54;
  assign GEN_56 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_55;
  assign GEN_57 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_56;
  assign GEN_58 = T_1421 ? 3'h4 : GEN_57;
  assign GEN_59 = T_1420 ? {{1'd0}, 2'h3} : GEN_58;
  assign GEN_60 = T_1419 ? {{1'd0}, 2'h2} : GEN_59;
  assign GEN_61 = T_1418 ? {{2'd0}, 1'h1} : GEN_60;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_65 = {1{$random}};
  T_1380 = GEN_65[2:0];
  GEN_66 = {1{$random}};
  T_1382 = GEN_66[2:0];
  GEN_67 = {1{$random}};
  lastGrant = GEN_67[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1380 <= 3'h0;
    end else begin
      T_1380 <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      T_1382 <= GEN_50;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_53;
    end
  end
endmodule
module BasicBus(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [2:0] io_in_0_bits_payload_a_type,
  input  [11:0] io_in_0_bits_payload_union,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [2:0] io_in_1_bits_payload_a_type,
  input  [11:0] io_in_1_bits_payload_union,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [2:0] io_in_2_bits_payload_a_type,
  input  [11:0] io_in_2_bits_payload_union,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [2:0] io_in_3_bits_payload_a_type,
  input  [11:0] io_in_3_bits_payload_union,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input   io_in_4_bits_payload_is_builtin_type,
  input  [2:0] io_in_4_bits_payload_a_type,
  input  [11:0] io_in_4_bits_payload_union,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [2:0] io_out_0_bits_header_src,
  output [2:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output  io_out_0_bits_payload_is_builtin_type,
  output [2:0] io_out_0_bits_payload_a_type,
  output [11:0] io_out_0_bits_payload_union,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [2:0] io_out_1_bits_header_src,
  output [2:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output  io_out_1_bits_payload_is_builtin_type,
  output [2:0] io_out_1_bits_payload_a_type,
  output [11:0] io_out_1_bits_payload_union,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [2:0] io_out_2_bits_header_src,
  output [2:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output  io_out_2_bits_payload_is_builtin_type,
  output [2:0] io_out_2_bits_payload_a_type,
  output [11:0] io_out_2_bits_payload_union,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [2:0] io_out_3_bits_header_src,
  output [2:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output  io_out_3_bits_payload_is_builtin_type,
  output [2:0] io_out_3_bits_payload_a_type,
  output [11:0] io_out_3_bits_payload_union,
  output [63:0] io_out_3_bits_payload_data,
  input   io_out_4_ready,
  output  io_out_4_valid,
  output [2:0] io_out_4_bits_header_src,
  output [2:0] io_out_4_bits_header_dst,
  output [25:0] io_out_4_bits_payload_addr_block,
  output [1:0] io_out_4_bits_payload_client_xact_id,
  output [2:0] io_out_4_bits_payload_addr_beat,
  output  io_out_4_bits_payload_is_builtin_type,
  output [2:0] io_out_4_bits_payload_a_type,
  output [11:0] io_out_4_bits_payload_union,
  output [63:0] io_out_4_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [2:0] arb_io_in_0_bits_header_src;
  wire [2:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_0_bits_payload_a_type;
  wire [11:0] arb_io_in_0_bits_payload_union;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [2:0] arb_io_in_1_bits_header_src;
  wire [2:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_1_bits_payload_a_type;
  wire [11:0] arb_io_in_1_bits_payload_union;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [2:0] arb_io_in_2_bits_header_src;
  wire [2:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_2_bits_payload_a_type;
  wire [11:0] arb_io_in_2_bits_payload_union;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [2:0] arb_io_in_3_bits_header_src;
  wire [2:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_3_bits_payload_a_type;
  wire [11:0] arb_io_in_3_bits_payload_union;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_in_4_ready;
  wire  arb_io_in_4_valid;
  wire [2:0] arb_io_in_4_bits_header_src;
  wire [2:0] arb_io_in_4_bits_header_dst;
  wire [25:0] arb_io_in_4_bits_payload_addr_block;
  wire [1:0] arb_io_in_4_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_4_bits_payload_addr_beat;
  wire  arb_io_in_4_bits_payload_is_builtin_type;
  wire [2:0] arb_io_in_4_bits_payload_a_type;
  wire [11:0] arb_io_in_4_bits_payload_union;
  wire [63:0] arb_io_in_4_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [2:0] arb_io_out_bits_header_src;
  wire [2:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [2:0] arb_io_out_bits_payload_a_type;
  wire [11:0] arb_io_out_bits_payload_union;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [2:0] arb_io_chosen;
  wire  GEN_0;
  wire [2:0] GEN_5;
  wire  GEN_1;
  wire [2:0] GEN_6;
  wire  GEN_2;
  wire [2:0] GEN_7;
  wire  GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_8;
  wire  T_1883;
  wire  T_1884;
  wire  T_1886;
  wire  T_1887;
  wire  T_1889;
  wire  T_1890;
  wire  T_1892;
  wire  T_1893;
  wire  T_1895;
  wire  T_1896;
  LockingRRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(arb_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(arb_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(arb_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(arb_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(arb_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(arb_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(arb_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(arb_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_in_4_ready(arb_io_in_4_ready),
    .io_in_4_valid(arb_io_in_4_valid),
    .io_in_4_bits_header_src(arb_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(arb_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_block(arb_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_client_xact_id(arb_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_addr_beat(arb_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_is_builtin_type(arb_io_in_4_bits_payload_is_builtin_type),
    .io_in_4_bits_payload_a_type(arb_io_in_4_bits_payload_a_type),
    .io_in_4_bits_payload_union(arb_io_in_4_bits_payload_union),
    .io_in_4_bits_payload_data(arb_io_in_4_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_a_type(arb_io_out_bits_payload_a_type),
    .io_out_bits_payload_union(arb_io_out_bits_payload_union),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_in_4_ready = arb_io_in_4_ready;
  assign io_out_0_valid = T_1884;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_0_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1887;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_1_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1890;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_2_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1893;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_3_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_4_valid = T_1896;
  assign io_out_4_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_4_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_4_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_4_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_4_bits_payload_a_type = arb_io_out_bits_payload_a_type;
  assign io_out_4_bits_payload_union = arb_io_out_bits_payload_union;
  assign io_out_4_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_a_type = io_in_0_bits_payload_a_type;
  assign arb_io_in_0_bits_payload_union = io_in_0_bits_payload_union;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_a_type = io_in_1_bits_payload_a_type;
  assign arb_io_in_1_bits_payload_union = io_in_1_bits_payload_union;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_a_type = io_in_2_bits_payload_a_type;
  assign arb_io_in_2_bits_payload_union = io_in_2_bits_payload_union;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_a_type = io_in_3_bits_payload_a_type;
  assign arb_io_in_3_bits_payload_union = io_in_3_bits_payload_union;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_in_4_valid = io_in_4_valid;
  assign arb_io_in_4_bits_header_src = io_in_4_bits_header_src;
  assign arb_io_in_4_bits_header_dst = io_in_4_bits_header_dst;
  assign arb_io_in_4_bits_payload_addr_block = io_in_4_bits_payload_addr_block;
  assign arb_io_in_4_bits_payload_client_xact_id = io_in_4_bits_payload_client_xact_id;
  assign arb_io_in_4_bits_payload_addr_beat = io_in_4_bits_payload_addr_beat;
  assign arb_io_in_4_bits_payload_is_builtin_type = io_in_4_bits_payload_is_builtin_type;
  assign arb_io_in_4_bits_payload_a_type = io_in_4_bits_payload_a_type;
  assign arb_io_in_4_bits_payload_union = io_in_4_bits_payload_union;
  assign arb_io_in_4_bits_payload_data = io_in_4_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_4;
  assign GEN_5 = {{2'd0}, 1'h1};
  assign GEN_1 = GEN_5 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_6 = {{1'd0}, 2'h2};
  assign GEN_2 = GEN_6 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = {{1'd0}, 2'h3};
  assign GEN_3 = GEN_7 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_4 = 3'h4 == arb_io_out_bits_header_dst ? io_out_4_ready : GEN_3;
  assign GEN_8 = {{2'd0}, 1'h0};
  assign T_1883 = arb_io_out_bits_header_dst == GEN_8;
  assign T_1884 = arb_io_out_valid & T_1883;
  assign T_1886 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1887 = arb_io_out_valid & T_1886;
  assign T_1889 = arb_io_out_bits_header_dst == GEN_6;
  assign T_1890 = arb_io_out_valid & T_1889;
  assign T_1892 = arb_io_out_bits_header_dst == GEN_7;
  assign T_1893 = arb_io_out_valid & T_1892;
  assign T_1895 = arb_io_out_bits_header_dst == 3'h4;
  assign T_1896 = arb_io_out_valid & T_1895;
endmodule
module LockingRRArbiter_21(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input   io_in_4_bits_payload_voluntary,
  input  [2:0] io_in_4_bits_payload_r_type,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_header_src,
  output [2:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_client_xact_id,
  output  io_out_bits_payload_voluntary,
  output [2:0] io_out_bits_payload_r_type,
  output [63:0] io_out_bits_payload_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_57;
  wire  GEN_9;
  wire [2:0] GEN_58;
  wire  GEN_10;
  wire [2:0] GEN_59;
  wire  GEN_11;
  wire  GEN_12;
  wire [2:0] GEN_1;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [2:0] GEN_16;
  wire [2:0] GEN_2;
  wire [2:0] GEN_17;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_3;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire [2:0] GEN_24;
  wire [25:0] GEN_4;
  wire [25:0] GEN_25;
  wire [25:0] GEN_26;
  wire [25:0] GEN_27;
  wire [25:0] GEN_28;
  wire [1:0] GEN_5;
  wire [1:0] GEN_29;
  wire [1:0] GEN_30;
  wire [1:0] GEN_31;
  wire [1:0] GEN_32;
  wire  GEN_6;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [2:0] GEN_7;
  wire [2:0] GEN_37;
  wire [2:0] GEN_38;
  wire [2:0] GEN_39;
  wire [2:0] GEN_40;
  wire [63:0] GEN_8;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  reg [2:0] T_1342;
  reg [31:0] GEN_60;
  reg [2:0] T_1344;
  reg [31:0] GEN_61;
  wire [2:0] GEN_84;
  wire  T_1346;
  wire [2:0] T_1353_0;
  wire [2:0] T_1353_1;
  wire [2:0] T_1353_2;
  wire  T_1355;
  wire  T_1356;
  wire  T_1357;
  wire  T_1360;
  wire  T_1361;
  wire  T_1363;
  wire  T_1364;
  wire [3:0] T_1368;
  wire [2:0] T_1369;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  reg [2:0] lastGrant;
  reg [31:0] GEN_62;
  wire [2:0] GEN_48;
  wire  T_1374;
  wire  T_1376;
  wire  T_1378;
  wire  T_1380;
  wire  T_1382;
  wire  T_1383;
  wire  T_1384;
  wire  T_1385;
  wire  T_1388;
  wire  T_1389;
  wire  T_1390;
  wire  T_1391;
  wire  T_1392;
  wire  T_1393;
  wire  T_1394;
  wire  T_1398;
  wire  T_1400;
  wire  T_1402;
  wire  T_1404;
  wire  T_1406;
  wire  T_1408;
  wire  T_1410;
  wire  T_1412;
  wire  T_1416;
  wire  T_1417;
  wire  T_1418;
  wire  T_1419;
  wire  T_1420;
  wire  T_1421;
  wire  T_1422;
  wire  T_1424;
  wire  T_1425;
  wire  T_1426;
  wire  T_1428;
  wire  T_1429;
  wire  T_1430;
  wire  T_1432;
  wire  T_1433;
  wire  T_1434;
  wire  T_1436;
  wire  T_1437;
  wire  T_1438;
  wire  T_1440;
  wire  T_1441;
  wire  T_1442;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  wire [2:0] GEN_52;
  wire [2:0] GEN_53;
  wire [2:0] GEN_54;
  wire [2:0] GEN_55;
  wire [2:0] GEN_56;
  assign io_in_0_ready = T_1426;
  assign io_in_1_ready = T_1430;
  assign io_in_2_ready = T_1434;
  assign io_in_3_ready = T_1438;
  assign io_in_4_ready = T_1442;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_addr_block = GEN_4;
  assign io_out_bits_payload_client_xact_id = GEN_5;
  assign io_out_bits_payload_voluntary = GEN_6;
  assign io_out_bits_payload_r_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_47;
  assign choice = GEN_56;
  assign GEN_0 = GEN_12;
  assign GEN_57 = {{2'd0}, 1'h1};
  assign GEN_9 = GEN_57 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_58 = {{1'd0}, 2'h2};
  assign GEN_10 = GEN_58 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_59 = {{1'd0}, 2'h3};
  assign GEN_11 = GEN_59 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_12 = 3'h4 == io_chosen ? io_in_4_valid : GEN_11;
  assign GEN_1 = GEN_16;
  assign GEN_13 = GEN_57 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_14 = GEN_58 == io_chosen ? io_in_2_bits_header_src : GEN_13;
  assign GEN_15 = GEN_59 == io_chosen ? io_in_3_bits_header_src : GEN_14;
  assign GEN_16 = 3'h4 == io_chosen ? io_in_4_bits_header_src : GEN_15;
  assign GEN_2 = GEN_20;
  assign GEN_17 = GEN_57 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_18 = GEN_58 == io_chosen ? io_in_2_bits_header_dst : GEN_17;
  assign GEN_19 = GEN_59 == io_chosen ? io_in_3_bits_header_dst : GEN_18;
  assign GEN_20 = 3'h4 == io_chosen ? io_in_4_bits_header_dst : GEN_19;
  assign GEN_3 = GEN_24;
  assign GEN_21 = GEN_57 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_22 = GEN_58 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_21;
  assign GEN_23 = GEN_59 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_22;
  assign GEN_24 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_beat : GEN_23;
  assign GEN_4 = GEN_28;
  assign GEN_25 = GEN_57 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_26 = GEN_58 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_25;
  assign GEN_27 = GEN_59 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_26;
  assign GEN_28 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_block : GEN_27;
  assign GEN_5 = GEN_32;
  assign GEN_29 = GEN_57 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_30 = GEN_58 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_29;
  assign GEN_31 = GEN_59 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_30;
  assign GEN_32 = 3'h4 == io_chosen ? io_in_4_bits_payload_client_xact_id : GEN_31;
  assign GEN_6 = GEN_36;
  assign GEN_33 = GEN_57 == io_chosen ? io_in_1_bits_payload_voluntary : io_in_0_bits_payload_voluntary;
  assign GEN_34 = GEN_58 == io_chosen ? io_in_2_bits_payload_voluntary : GEN_33;
  assign GEN_35 = GEN_59 == io_chosen ? io_in_3_bits_payload_voluntary : GEN_34;
  assign GEN_36 = 3'h4 == io_chosen ? io_in_4_bits_payload_voluntary : GEN_35;
  assign GEN_7 = GEN_40;
  assign GEN_37 = GEN_57 == io_chosen ? io_in_1_bits_payload_r_type : io_in_0_bits_payload_r_type;
  assign GEN_38 = GEN_58 == io_chosen ? io_in_2_bits_payload_r_type : GEN_37;
  assign GEN_39 = GEN_59 == io_chosen ? io_in_3_bits_payload_r_type : GEN_38;
  assign GEN_40 = 3'h4 == io_chosen ? io_in_4_bits_payload_r_type : GEN_39;
  assign GEN_8 = GEN_44;
  assign GEN_41 = GEN_57 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_42 = GEN_58 == io_chosen ? io_in_2_bits_payload_data : GEN_41;
  assign GEN_43 = GEN_59 == io_chosen ? io_in_3_bits_payload_data : GEN_42;
  assign GEN_44 = 3'h4 == io_chosen ? io_in_4_bits_payload_data : GEN_43;
  assign GEN_84 = {{2'd0}, 1'h0};
  assign T_1346 = T_1342 != GEN_84;
  assign T_1353_0 = 3'h0;
  assign T_1353_1 = 3'h1;
  assign T_1353_2 = 3'h2;
  assign T_1355 = T_1353_0 == io_out_bits_payload_r_type;
  assign T_1356 = T_1353_1 == io_out_bits_payload_r_type;
  assign T_1357 = T_1353_2 == io_out_bits_payload_r_type;
  assign T_1360 = T_1355 | T_1356;
  assign T_1361 = T_1360 | T_1357;
  assign T_1363 = io_out_ready & io_out_valid;
  assign T_1364 = T_1363 & T_1361;
  assign T_1368 = T_1342 + GEN_57;
  assign T_1369 = T_1368[2:0];
  assign GEN_45 = T_1364 ? io_chosen : T_1344;
  assign GEN_46 = T_1364 ? T_1369 : T_1342;
  assign GEN_47 = T_1346 ? T_1344 : choice;
  assign GEN_48 = T_1363 ? io_chosen : lastGrant;
  assign T_1374 = GEN_57 > lastGrant;
  assign T_1376 = GEN_58 > lastGrant;
  assign T_1378 = GEN_59 > lastGrant;
  assign T_1380 = 3'h4 > lastGrant;
  assign T_1382 = io_in_1_valid & T_1374;
  assign T_1383 = io_in_2_valid & T_1376;
  assign T_1384 = io_in_3_valid & T_1378;
  assign T_1385 = io_in_4_valid & T_1380;
  assign T_1388 = T_1382 | T_1383;
  assign T_1389 = T_1388 | T_1384;
  assign T_1390 = T_1389 | T_1385;
  assign T_1391 = T_1390 | io_in_0_valid;
  assign T_1392 = T_1391 | io_in_1_valid;
  assign T_1393 = T_1392 | io_in_2_valid;
  assign T_1394 = T_1393 | io_in_3_valid;
  assign T_1398 = T_1382 == 1'h0;
  assign T_1400 = T_1388 == 1'h0;
  assign T_1402 = T_1389 == 1'h0;
  assign T_1404 = T_1390 == 1'h0;
  assign T_1406 = T_1391 == 1'h0;
  assign T_1408 = T_1392 == 1'h0;
  assign T_1410 = T_1393 == 1'h0;
  assign T_1412 = T_1394 == 1'h0;
  assign T_1416 = T_1374 | T_1406;
  assign T_1417 = T_1398 & T_1376;
  assign T_1418 = T_1417 | T_1408;
  assign T_1419 = T_1400 & T_1378;
  assign T_1420 = T_1419 | T_1410;
  assign T_1421 = T_1402 & T_1380;
  assign T_1422 = T_1421 | T_1412;
  assign T_1424 = T_1344 == GEN_84;
  assign T_1425 = T_1346 ? T_1424 : T_1404;
  assign T_1426 = T_1425 & io_out_ready;
  assign T_1428 = T_1344 == GEN_57;
  assign T_1429 = T_1346 ? T_1428 : T_1416;
  assign T_1430 = T_1429 & io_out_ready;
  assign T_1432 = T_1344 == GEN_58;
  assign T_1433 = T_1346 ? T_1432 : T_1418;
  assign T_1434 = T_1433 & io_out_ready;
  assign T_1436 = T_1344 == GEN_59;
  assign T_1437 = T_1346 ? T_1436 : T_1420;
  assign T_1438 = T_1437 & io_out_ready;
  assign T_1440 = T_1344 == 3'h4;
  assign T_1441 = T_1346 ? T_1440 : T_1422;
  assign T_1442 = T_1441 & io_out_ready;
  assign GEN_49 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_50 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_50;
  assign GEN_52 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_51;
  assign GEN_53 = T_1385 ? 3'h4 : GEN_52;
  assign GEN_54 = T_1384 ? {{1'd0}, 2'h3} : GEN_53;
  assign GEN_55 = T_1383 ? {{1'd0}, 2'h2} : GEN_54;
  assign GEN_56 = T_1382 ? {{2'd0}, 1'h1} : GEN_55;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_60 = {1{$random}};
  T_1342 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_1344 = GEN_61[2:0];
  GEN_62 = {1{$random}};
  lastGrant = GEN_62[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1342 <= 3'h0;
    end else begin
      T_1342 <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      T_1344 <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_48;
    end
  end
endmodule
module BasicBus_20(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input   io_in_0_bits_payload_voluntary,
  input  [2:0] io_in_0_bits_payload_r_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input   io_in_1_bits_payload_voluntary,
  input  [2:0] io_in_1_bits_payload_r_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input   io_in_2_bits_payload_voluntary,
  input  [2:0] io_in_2_bits_payload_r_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input   io_in_3_bits_payload_voluntary,
  input  [2:0] io_in_3_bits_payload_r_type,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input   io_in_4_bits_payload_voluntary,
  input  [2:0] io_in_4_bits_payload_r_type,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [2:0] io_out_0_bits_header_src,
  output [2:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output  io_out_0_bits_payload_voluntary,
  output [2:0] io_out_0_bits_payload_r_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [2:0] io_out_1_bits_header_src,
  output [2:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output  io_out_1_bits_payload_voluntary,
  output [2:0] io_out_1_bits_payload_r_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [2:0] io_out_2_bits_header_src,
  output [2:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output  io_out_2_bits_payload_voluntary,
  output [2:0] io_out_2_bits_payload_r_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [2:0] io_out_3_bits_header_src,
  output [2:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output  io_out_3_bits_payload_voluntary,
  output [2:0] io_out_3_bits_payload_r_type,
  output [63:0] io_out_3_bits_payload_data,
  input   io_out_4_ready,
  output  io_out_4_valid,
  output [2:0] io_out_4_bits_header_src,
  output [2:0] io_out_4_bits_header_dst,
  output [2:0] io_out_4_bits_payload_addr_beat,
  output [25:0] io_out_4_bits_payload_addr_block,
  output [1:0] io_out_4_bits_payload_client_xact_id,
  output  io_out_4_bits_payload_voluntary,
  output [2:0] io_out_4_bits_payload_r_type,
  output [63:0] io_out_4_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [2:0] arb_io_in_0_bits_header_src;
  wire [2:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire  arb_io_in_0_bits_payload_voluntary;
  wire [2:0] arb_io_in_0_bits_payload_r_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [2:0] arb_io_in_1_bits_header_src;
  wire [2:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire  arb_io_in_1_bits_payload_voluntary;
  wire [2:0] arb_io_in_1_bits_payload_r_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [2:0] arb_io_in_2_bits_header_src;
  wire [2:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire  arb_io_in_2_bits_payload_voluntary;
  wire [2:0] arb_io_in_2_bits_payload_r_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [2:0] arb_io_in_3_bits_header_src;
  wire [2:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire  arb_io_in_3_bits_payload_voluntary;
  wire [2:0] arb_io_in_3_bits_payload_r_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_in_4_ready;
  wire  arb_io_in_4_valid;
  wire [2:0] arb_io_in_4_bits_header_src;
  wire [2:0] arb_io_in_4_bits_header_dst;
  wire [2:0] arb_io_in_4_bits_payload_addr_beat;
  wire [25:0] arb_io_in_4_bits_payload_addr_block;
  wire [1:0] arb_io_in_4_bits_payload_client_xact_id;
  wire  arb_io_in_4_bits_payload_voluntary;
  wire [2:0] arb_io_in_4_bits_payload_r_type;
  wire [63:0] arb_io_in_4_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [2:0] arb_io_out_bits_header_src;
  wire [2:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire  arb_io_out_bits_payload_voluntary;
  wire [2:0] arb_io_out_bits_payload_r_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [2:0] arb_io_chosen;
  wire  GEN_0;
  wire [2:0] GEN_5;
  wire  GEN_1;
  wire [2:0] GEN_6;
  wire  GEN_2;
  wire [2:0] GEN_7;
  wire  GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_8;
  wire  T_1831;
  wire  T_1832;
  wire  T_1834;
  wire  T_1835;
  wire  T_1837;
  wire  T_1838;
  wire  T_1840;
  wire  T_1841;
  wire  T_1843;
  wire  T_1844;
  LockingRRArbiter_21 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(arb_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(arb_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(arb_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(arb_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(arb_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(arb_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(arb_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(arb_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_in_4_ready(arb_io_in_4_ready),
    .io_in_4_valid(arb_io_in_4_valid),
    .io_in_4_bits_header_src(arb_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(arb_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_beat(arb_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_addr_block(arb_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_client_xact_id(arb_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_voluntary(arb_io_in_4_bits_payload_voluntary),
    .io_in_4_bits_payload_r_type(arb_io_in_4_bits_payload_r_type),
    .io_in_4_bits_payload_data(arb_io_in_4_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_voluntary(arb_io_out_bits_payload_voluntary),
    .io_out_bits_payload_r_type(arb_io_out_bits_payload_r_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_in_4_ready = arb_io_in_4_ready;
  assign io_out_0_valid = T_1832;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_0_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1835;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_1_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1838;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_2_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1841;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_3_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_4_valid = T_1844;
  assign io_out_4_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_4_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_4_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_4_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_voluntary = arb_io_out_bits_payload_voluntary;
  assign io_out_4_bits_payload_r_type = arb_io_out_bits_payload_r_type;
  assign io_out_4_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_voluntary = io_in_0_bits_payload_voluntary;
  assign arb_io_in_0_bits_payload_r_type = io_in_0_bits_payload_r_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_voluntary = io_in_1_bits_payload_voluntary;
  assign arb_io_in_1_bits_payload_r_type = io_in_1_bits_payload_r_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_voluntary = io_in_2_bits_payload_voluntary;
  assign arb_io_in_2_bits_payload_r_type = io_in_2_bits_payload_r_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_voluntary = io_in_3_bits_payload_voluntary;
  assign arb_io_in_3_bits_payload_r_type = io_in_3_bits_payload_r_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_in_4_valid = io_in_4_valid;
  assign arb_io_in_4_bits_header_src = io_in_4_bits_header_src;
  assign arb_io_in_4_bits_header_dst = io_in_4_bits_header_dst;
  assign arb_io_in_4_bits_payload_addr_beat = io_in_4_bits_payload_addr_beat;
  assign arb_io_in_4_bits_payload_addr_block = io_in_4_bits_payload_addr_block;
  assign arb_io_in_4_bits_payload_client_xact_id = io_in_4_bits_payload_client_xact_id;
  assign arb_io_in_4_bits_payload_voluntary = io_in_4_bits_payload_voluntary;
  assign arb_io_in_4_bits_payload_r_type = io_in_4_bits_payload_r_type;
  assign arb_io_in_4_bits_payload_data = io_in_4_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_4;
  assign GEN_5 = {{2'd0}, 1'h1};
  assign GEN_1 = GEN_5 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_6 = {{1'd0}, 2'h2};
  assign GEN_2 = GEN_6 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = {{1'd0}, 2'h3};
  assign GEN_3 = GEN_7 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_4 = 3'h4 == arb_io_out_bits_header_dst ? io_out_4_ready : GEN_3;
  assign GEN_8 = {{2'd0}, 1'h0};
  assign T_1831 = arb_io_out_bits_header_dst == GEN_8;
  assign T_1832 = arb_io_out_valid & T_1831;
  assign T_1834 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1835 = arb_io_out_valid & T_1834;
  assign T_1837 = arb_io_out_bits_header_dst == GEN_6;
  assign T_1838 = arb_io_out_valid & T_1837;
  assign T_1840 = arb_io_out_bits_header_dst == GEN_7;
  assign T_1841 = arb_io_out_valid & T_1840;
  assign T_1843 = arb_io_out_bits_header_dst == 3'h4;
  assign T_1844 = arb_io_out_valid & T_1843;
endmodule
module LockingRRArbiter_23(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_p_type,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_header_src,
  output [2:0] io_out_bits_header_dst,
  output [25:0] io_out_bits_payload_addr_block,
  output [1:0] io_out_bits_payload_p_type,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_34;
  wire  GEN_5;
  wire [2:0] GEN_35;
  wire  GEN_6;
  wire [2:0] GEN_36;
  wire  GEN_7;
  wire  GEN_8;
  wire [2:0] GEN_1;
  wire [2:0] GEN_9;
  wire [2:0] GEN_10;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire [2:0] GEN_2;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [2:0] GEN_16;
  wire [25:0] GEN_3;
  wire [25:0] GEN_17;
  wire [25:0] GEN_18;
  wire [25:0] GEN_19;
  wire [25:0] GEN_20;
  wire [1:0] GEN_4;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_24;
  wire  T_1190;
  reg [2:0] lastGrant;
  reg [31:0] GEN_37;
  wire [2:0] GEN_25;
  wire  T_1193;
  wire  T_1195;
  wire  T_1197;
  wire  T_1199;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1204;
  wire  T_1207;
  wire  T_1208;
  wire  T_1209;
  wire  T_1210;
  wire  T_1211;
  wire  T_1212;
  wire  T_1213;
  wire  T_1217;
  wire  T_1219;
  wire  T_1221;
  wire  T_1223;
  wire  T_1225;
  wire  T_1227;
  wire  T_1229;
  wire  T_1231;
  wire  T_1235;
  wire  T_1236;
  wire  T_1237;
  wire  T_1238;
  wire  T_1239;
  wire  T_1240;
  wire  T_1241;
  wire  T_1242;
  wire  T_1243;
  wire  T_1244;
  wire  T_1245;
  wire  T_1246;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire [2:0] GEN_33;
  assign io_in_0_ready = T_1242;
  assign io_in_1_ready = T_1243;
  assign io_in_2_ready = T_1244;
  assign io_in_3_ready = T_1245;
  assign io_in_4_ready = T_1246;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_block = GEN_3;
  assign io_out_bits_payload_p_type = GEN_4;
  assign io_chosen = choice;
  assign choice = GEN_33;
  assign GEN_0 = GEN_8;
  assign GEN_34 = {{2'd0}, 1'h1};
  assign GEN_5 = GEN_34 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_35 = {{1'd0}, 2'h2};
  assign GEN_6 = GEN_35 == io_chosen ? io_in_2_valid : GEN_5;
  assign GEN_36 = {{1'd0}, 2'h3};
  assign GEN_7 = GEN_36 == io_chosen ? io_in_3_valid : GEN_6;
  assign GEN_8 = 3'h4 == io_chosen ? io_in_4_valid : GEN_7;
  assign GEN_1 = GEN_12;
  assign GEN_9 = GEN_34 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_10 = GEN_35 == io_chosen ? io_in_2_bits_header_src : GEN_9;
  assign GEN_11 = GEN_36 == io_chosen ? io_in_3_bits_header_src : GEN_10;
  assign GEN_12 = 3'h4 == io_chosen ? io_in_4_bits_header_src : GEN_11;
  assign GEN_2 = GEN_16;
  assign GEN_13 = GEN_34 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_14 = GEN_35 == io_chosen ? io_in_2_bits_header_dst : GEN_13;
  assign GEN_15 = GEN_36 == io_chosen ? io_in_3_bits_header_dst : GEN_14;
  assign GEN_16 = 3'h4 == io_chosen ? io_in_4_bits_header_dst : GEN_15;
  assign GEN_3 = GEN_20;
  assign GEN_17 = GEN_34 == io_chosen ? io_in_1_bits_payload_addr_block : io_in_0_bits_payload_addr_block;
  assign GEN_18 = GEN_35 == io_chosen ? io_in_2_bits_payload_addr_block : GEN_17;
  assign GEN_19 = GEN_36 == io_chosen ? io_in_3_bits_payload_addr_block : GEN_18;
  assign GEN_20 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_block : GEN_19;
  assign GEN_4 = GEN_24;
  assign GEN_21 = GEN_34 == io_chosen ? io_in_1_bits_payload_p_type : io_in_0_bits_payload_p_type;
  assign GEN_22 = GEN_35 == io_chosen ? io_in_2_bits_payload_p_type : GEN_21;
  assign GEN_23 = GEN_36 == io_chosen ? io_in_3_bits_payload_p_type : GEN_22;
  assign GEN_24 = 3'h4 == io_chosen ? io_in_4_bits_payload_p_type : GEN_23;
  assign T_1190 = io_out_ready & io_out_valid;
  assign GEN_25 = T_1190 ? io_chosen : lastGrant;
  assign T_1193 = GEN_34 > lastGrant;
  assign T_1195 = GEN_35 > lastGrant;
  assign T_1197 = GEN_36 > lastGrant;
  assign T_1199 = 3'h4 > lastGrant;
  assign T_1201 = io_in_1_valid & T_1193;
  assign T_1202 = io_in_2_valid & T_1195;
  assign T_1203 = io_in_3_valid & T_1197;
  assign T_1204 = io_in_4_valid & T_1199;
  assign T_1207 = T_1201 | T_1202;
  assign T_1208 = T_1207 | T_1203;
  assign T_1209 = T_1208 | T_1204;
  assign T_1210 = T_1209 | io_in_0_valid;
  assign T_1211 = T_1210 | io_in_1_valid;
  assign T_1212 = T_1211 | io_in_2_valid;
  assign T_1213 = T_1212 | io_in_3_valid;
  assign T_1217 = T_1201 == 1'h0;
  assign T_1219 = T_1207 == 1'h0;
  assign T_1221 = T_1208 == 1'h0;
  assign T_1223 = T_1209 == 1'h0;
  assign T_1225 = T_1210 == 1'h0;
  assign T_1227 = T_1211 == 1'h0;
  assign T_1229 = T_1212 == 1'h0;
  assign T_1231 = T_1213 == 1'h0;
  assign T_1235 = T_1193 | T_1225;
  assign T_1236 = T_1217 & T_1195;
  assign T_1237 = T_1236 | T_1227;
  assign T_1238 = T_1219 & T_1197;
  assign T_1239 = T_1238 | T_1229;
  assign T_1240 = T_1221 & T_1199;
  assign T_1241 = T_1240 | T_1231;
  assign T_1242 = T_1223 & io_out_ready;
  assign T_1243 = T_1235 & io_out_ready;
  assign T_1244 = T_1237 & io_out_ready;
  assign T_1245 = T_1239 & io_out_ready;
  assign T_1246 = T_1241 & io_out_ready;
  assign GEN_26 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_27 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_26;
  assign GEN_28 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_27;
  assign GEN_29 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_28;
  assign GEN_30 = T_1204 ? 3'h4 : GEN_29;
  assign GEN_31 = T_1203 ? {{1'd0}, 2'h3} : GEN_30;
  assign GEN_32 = T_1202 ? {{1'd0}, 2'h2} : GEN_31;
  assign GEN_33 = T_1201 ? {{2'd0}, 1'h1} : GEN_32;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_37 = {1{$random}};
  lastGrant = GEN_37[2:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_25;
    end
  end
endmodule
module BasicBus_22(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [25:0] io_in_0_bits_payload_addr_block,
  input  [1:0] io_in_0_bits_payload_p_type,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [25:0] io_in_1_bits_payload_addr_block,
  input  [1:0] io_in_1_bits_payload_p_type,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [25:0] io_in_2_bits_payload_addr_block,
  input  [1:0] io_in_2_bits_payload_p_type,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [25:0] io_in_3_bits_payload_addr_block,
  input  [1:0] io_in_3_bits_payload_p_type,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [25:0] io_in_4_bits_payload_addr_block,
  input  [1:0] io_in_4_bits_payload_p_type,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [2:0] io_out_0_bits_header_src,
  output [2:0] io_out_0_bits_header_dst,
  output [25:0] io_out_0_bits_payload_addr_block,
  output [1:0] io_out_0_bits_payload_p_type,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [2:0] io_out_1_bits_header_src,
  output [2:0] io_out_1_bits_header_dst,
  output [25:0] io_out_1_bits_payload_addr_block,
  output [1:0] io_out_1_bits_payload_p_type,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [2:0] io_out_2_bits_header_src,
  output [2:0] io_out_2_bits_header_dst,
  output [25:0] io_out_2_bits_payload_addr_block,
  output [1:0] io_out_2_bits_payload_p_type,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [2:0] io_out_3_bits_header_src,
  output [2:0] io_out_3_bits_header_dst,
  output [25:0] io_out_3_bits_payload_addr_block,
  output [1:0] io_out_3_bits_payload_p_type,
  input   io_out_4_ready,
  output  io_out_4_valid,
  output [2:0] io_out_4_bits_header_src,
  output [2:0] io_out_4_bits_header_dst,
  output [25:0] io_out_4_bits_payload_addr_block,
  output [1:0] io_out_4_bits_payload_p_type
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [2:0] arb_io_in_0_bits_header_src;
  wire [2:0] arb_io_in_0_bits_header_dst;
  wire [25:0] arb_io_in_0_bits_payload_addr_block;
  wire [1:0] arb_io_in_0_bits_payload_p_type;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [2:0] arb_io_in_1_bits_header_src;
  wire [2:0] arb_io_in_1_bits_header_dst;
  wire [25:0] arb_io_in_1_bits_payload_addr_block;
  wire [1:0] arb_io_in_1_bits_payload_p_type;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [2:0] arb_io_in_2_bits_header_src;
  wire [2:0] arb_io_in_2_bits_header_dst;
  wire [25:0] arb_io_in_2_bits_payload_addr_block;
  wire [1:0] arb_io_in_2_bits_payload_p_type;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [2:0] arb_io_in_3_bits_header_src;
  wire [2:0] arb_io_in_3_bits_header_dst;
  wire [25:0] arb_io_in_3_bits_payload_addr_block;
  wire [1:0] arb_io_in_3_bits_payload_p_type;
  wire  arb_io_in_4_ready;
  wire  arb_io_in_4_valid;
  wire [2:0] arb_io_in_4_bits_header_src;
  wire [2:0] arb_io_in_4_bits_header_dst;
  wire [25:0] arb_io_in_4_bits_payload_addr_block;
  wire [1:0] arb_io_in_4_bits_payload_p_type;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [2:0] arb_io_out_bits_header_src;
  wire [2:0] arb_io_out_bits_header_dst;
  wire [25:0] arb_io_out_bits_payload_addr_block;
  wire [1:0] arb_io_out_bits_payload_p_type;
  wire [2:0] arb_io_chosen;
  wire  GEN_0;
  wire [2:0] GEN_5;
  wire  GEN_1;
  wire [2:0] GEN_6;
  wire  GEN_2;
  wire [2:0] GEN_7;
  wire  GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_8;
  wire  T_1623;
  wire  T_1624;
  wire  T_1626;
  wire  T_1627;
  wire  T_1629;
  wire  T_1630;
  wire  T_1632;
  wire  T_1633;
  wire  T_1635;
  wire  T_1636;
  LockingRRArbiter_23 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(arb_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(arb_io_in_0_bits_payload_p_type),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(arb_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(arb_io_in_1_bits_payload_p_type),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(arb_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(arb_io_in_2_bits_payload_p_type),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(arb_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(arb_io_in_3_bits_payload_p_type),
    .io_in_4_ready(arb_io_in_4_ready),
    .io_in_4_valid(arb_io_in_4_valid),
    .io_in_4_bits_header_src(arb_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(arb_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_block(arb_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_p_type(arb_io_in_4_bits_payload_p_type),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_block(arb_io_out_bits_payload_addr_block),
    .io_out_bits_payload_p_type(arb_io_out_bits_payload_p_type),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_in_4_ready = arb_io_in_4_ready;
  assign io_out_0_valid = T_1624;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_0_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_1_valid = T_1627;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_1_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_2_valid = T_1630;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_2_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_3_valid = T_1633;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_3_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign io_out_4_valid = T_1636;
  assign io_out_4_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_4_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_4_bits_payload_addr_block = arb_io_out_bits_payload_addr_block;
  assign io_out_4_bits_payload_p_type = arb_io_out_bits_payload_p_type;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_block = io_in_0_bits_payload_addr_block;
  assign arb_io_in_0_bits_payload_p_type = io_in_0_bits_payload_p_type;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_block = io_in_1_bits_payload_addr_block;
  assign arb_io_in_1_bits_payload_p_type = io_in_1_bits_payload_p_type;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_block = io_in_2_bits_payload_addr_block;
  assign arb_io_in_2_bits_payload_p_type = io_in_2_bits_payload_p_type;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_block = io_in_3_bits_payload_addr_block;
  assign arb_io_in_3_bits_payload_p_type = io_in_3_bits_payload_p_type;
  assign arb_io_in_4_valid = io_in_4_valid;
  assign arb_io_in_4_bits_header_src = io_in_4_bits_header_src;
  assign arb_io_in_4_bits_header_dst = io_in_4_bits_header_dst;
  assign arb_io_in_4_bits_payload_addr_block = io_in_4_bits_payload_addr_block;
  assign arb_io_in_4_bits_payload_p_type = io_in_4_bits_payload_p_type;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_4;
  assign GEN_5 = {{2'd0}, 1'h1};
  assign GEN_1 = GEN_5 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_6 = {{1'd0}, 2'h2};
  assign GEN_2 = GEN_6 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = {{1'd0}, 2'h3};
  assign GEN_3 = GEN_7 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_4 = 3'h4 == arb_io_out_bits_header_dst ? io_out_4_ready : GEN_3;
  assign GEN_8 = {{2'd0}, 1'h0};
  assign T_1623 = arb_io_out_bits_header_dst == GEN_8;
  assign T_1624 = arb_io_out_valid & T_1623;
  assign T_1626 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1627 = arb_io_out_valid & T_1626;
  assign T_1629 = arb_io_out_bits_header_dst == GEN_6;
  assign T_1630 = arb_io_out_valid & T_1629;
  assign T_1632 = arb_io_out_bits_header_dst == GEN_7;
  assign T_1633 = arb_io_out_valid & T_1632;
  assign T_1635 = arb_io_out_bits_header_dst == 3'h4;
  assign T_1636 = arb_io_out_valid & T_1635;
endmodule
module LockingRRArbiter_25(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input  [2:0] io_in_4_bits_payload_manager_xact_id,
  input   io_in_4_bits_payload_is_builtin_type,
  input  [3:0] io_in_4_bits_payload_g_type,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_header_src,
  output [2:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_addr_beat,
  output [1:0] io_out_bits_payload_client_xact_id,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output  io_out_bits_payload_is_builtin_type,
  output [3:0] io_out_bits_payload_g_type,
  output [63:0] io_out_bits_payload_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_57;
  wire  GEN_9;
  wire [2:0] GEN_58;
  wire  GEN_10;
  wire [2:0] GEN_59;
  wire  GEN_11;
  wire  GEN_12;
  wire [2:0] GEN_1;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [2:0] GEN_16;
  wire [2:0] GEN_2;
  wire [2:0] GEN_17;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_20;
  wire [2:0] GEN_3;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire [2:0] GEN_24;
  wire [1:0] GEN_4;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  wire [2:0] GEN_5;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [2:0] GEN_32;
  wire  GEN_6;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [3:0] GEN_7;
  wire [3:0] GEN_37;
  wire [3:0] GEN_38;
  wire [3:0] GEN_39;
  wire [3:0] GEN_40;
  wire [63:0] GEN_8;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  reg [2:0] T_1342;
  reg [31:0] GEN_60;
  reg [2:0] T_1344;
  reg [31:0] GEN_61;
  wire [2:0] GEN_84;
  wire  T_1346;
  wire [2:0] T_1354_0;
  wire [3:0] GEN_85;
  wire  T_1356;
  wire [1:0] T_1364_0;
  wire [1:0] T_1364_1;
  wire [3:0] GEN_86;
  wire  T_1366;
  wire [3:0] GEN_87;
  wire  T_1367;
  wire  T_1370;
  wire  T_1371;
  wire  T_1373;
  wire  T_1374;
  wire [3:0] T_1378;
  wire [2:0] T_1379;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  reg [2:0] lastGrant;
  reg [31:0] GEN_62;
  wire [2:0] GEN_48;
  wire  T_1384;
  wire  T_1386;
  wire  T_1388;
  wire  T_1390;
  wire  T_1392;
  wire  T_1393;
  wire  T_1394;
  wire  T_1395;
  wire  T_1398;
  wire  T_1399;
  wire  T_1400;
  wire  T_1401;
  wire  T_1402;
  wire  T_1403;
  wire  T_1404;
  wire  T_1408;
  wire  T_1410;
  wire  T_1412;
  wire  T_1414;
  wire  T_1416;
  wire  T_1418;
  wire  T_1420;
  wire  T_1422;
  wire  T_1426;
  wire  T_1427;
  wire  T_1428;
  wire  T_1429;
  wire  T_1430;
  wire  T_1431;
  wire  T_1432;
  wire  T_1434;
  wire  T_1435;
  wire  T_1436;
  wire  T_1438;
  wire  T_1439;
  wire  T_1440;
  wire  T_1442;
  wire  T_1443;
  wire  T_1444;
  wire  T_1446;
  wire  T_1447;
  wire  T_1448;
  wire  T_1450;
  wire  T_1451;
  wire  T_1452;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  wire [2:0] GEN_52;
  wire [2:0] GEN_53;
  wire [2:0] GEN_54;
  wire [2:0] GEN_55;
  wire [2:0] GEN_56;
  assign io_in_0_ready = T_1436;
  assign io_in_1_ready = T_1440;
  assign io_in_2_ready = T_1444;
  assign io_in_3_ready = T_1448;
  assign io_in_4_ready = T_1452;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_addr_beat = GEN_3;
  assign io_out_bits_payload_client_xact_id = GEN_4;
  assign io_out_bits_payload_manager_xact_id = GEN_5;
  assign io_out_bits_payload_is_builtin_type = GEN_6;
  assign io_out_bits_payload_g_type = GEN_7;
  assign io_out_bits_payload_data = GEN_8;
  assign io_chosen = GEN_47;
  assign choice = GEN_56;
  assign GEN_0 = GEN_12;
  assign GEN_57 = {{2'd0}, 1'h1};
  assign GEN_9 = GEN_57 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_58 = {{1'd0}, 2'h2};
  assign GEN_10 = GEN_58 == io_chosen ? io_in_2_valid : GEN_9;
  assign GEN_59 = {{1'd0}, 2'h3};
  assign GEN_11 = GEN_59 == io_chosen ? io_in_3_valid : GEN_10;
  assign GEN_12 = 3'h4 == io_chosen ? io_in_4_valid : GEN_11;
  assign GEN_1 = GEN_16;
  assign GEN_13 = GEN_57 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_14 = GEN_58 == io_chosen ? io_in_2_bits_header_src : GEN_13;
  assign GEN_15 = GEN_59 == io_chosen ? io_in_3_bits_header_src : GEN_14;
  assign GEN_16 = 3'h4 == io_chosen ? io_in_4_bits_header_src : GEN_15;
  assign GEN_2 = GEN_20;
  assign GEN_17 = GEN_57 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_18 = GEN_58 == io_chosen ? io_in_2_bits_header_dst : GEN_17;
  assign GEN_19 = GEN_59 == io_chosen ? io_in_3_bits_header_dst : GEN_18;
  assign GEN_20 = 3'h4 == io_chosen ? io_in_4_bits_header_dst : GEN_19;
  assign GEN_3 = GEN_24;
  assign GEN_21 = GEN_57 == io_chosen ? io_in_1_bits_payload_addr_beat : io_in_0_bits_payload_addr_beat;
  assign GEN_22 = GEN_58 == io_chosen ? io_in_2_bits_payload_addr_beat : GEN_21;
  assign GEN_23 = GEN_59 == io_chosen ? io_in_3_bits_payload_addr_beat : GEN_22;
  assign GEN_24 = 3'h4 == io_chosen ? io_in_4_bits_payload_addr_beat : GEN_23;
  assign GEN_4 = GEN_28;
  assign GEN_25 = GEN_57 == io_chosen ? io_in_1_bits_payload_client_xact_id : io_in_0_bits_payload_client_xact_id;
  assign GEN_26 = GEN_58 == io_chosen ? io_in_2_bits_payload_client_xact_id : GEN_25;
  assign GEN_27 = GEN_59 == io_chosen ? io_in_3_bits_payload_client_xact_id : GEN_26;
  assign GEN_28 = 3'h4 == io_chosen ? io_in_4_bits_payload_client_xact_id : GEN_27;
  assign GEN_5 = GEN_32;
  assign GEN_29 = GEN_57 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_30 = GEN_58 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_29;
  assign GEN_31 = GEN_59 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_30;
  assign GEN_32 = 3'h4 == io_chosen ? io_in_4_bits_payload_manager_xact_id : GEN_31;
  assign GEN_6 = GEN_36;
  assign GEN_33 = GEN_57 == io_chosen ? io_in_1_bits_payload_is_builtin_type : io_in_0_bits_payload_is_builtin_type;
  assign GEN_34 = GEN_58 == io_chosen ? io_in_2_bits_payload_is_builtin_type : GEN_33;
  assign GEN_35 = GEN_59 == io_chosen ? io_in_3_bits_payload_is_builtin_type : GEN_34;
  assign GEN_36 = 3'h4 == io_chosen ? io_in_4_bits_payload_is_builtin_type : GEN_35;
  assign GEN_7 = GEN_40;
  assign GEN_37 = GEN_57 == io_chosen ? io_in_1_bits_payload_g_type : io_in_0_bits_payload_g_type;
  assign GEN_38 = GEN_58 == io_chosen ? io_in_2_bits_payload_g_type : GEN_37;
  assign GEN_39 = GEN_59 == io_chosen ? io_in_3_bits_payload_g_type : GEN_38;
  assign GEN_40 = 3'h4 == io_chosen ? io_in_4_bits_payload_g_type : GEN_39;
  assign GEN_8 = GEN_44;
  assign GEN_41 = GEN_57 == io_chosen ? io_in_1_bits_payload_data : io_in_0_bits_payload_data;
  assign GEN_42 = GEN_58 == io_chosen ? io_in_2_bits_payload_data : GEN_41;
  assign GEN_43 = GEN_59 == io_chosen ? io_in_3_bits_payload_data : GEN_42;
  assign GEN_44 = 3'h4 == io_chosen ? io_in_4_bits_payload_data : GEN_43;
  assign GEN_84 = {{2'd0}, 1'h0};
  assign T_1346 = T_1342 != GEN_84;
  assign T_1354_0 = 3'h5;
  assign GEN_85 = {{1'd0}, T_1354_0};
  assign T_1356 = GEN_85 == io_out_bits_payload_g_type;
  assign T_1364_0 = 2'h0;
  assign T_1364_1 = 2'h1;
  assign GEN_86 = {{2'd0}, T_1364_0};
  assign T_1366 = GEN_86 == io_out_bits_payload_g_type;
  assign GEN_87 = {{2'd0}, T_1364_1};
  assign T_1367 = GEN_87 == io_out_bits_payload_g_type;
  assign T_1370 = T_1366 | T_1367;
  assign T_1371 = io_out_bits_payload_is_builtin_type ? T_1356 : T_1370;
  assign T_1373 = io_out_ready & io_out_valid;
  assign T_1374 = T_1373 & T_1371;
  assign T_1378 = T_1342 + GEN_57;
  assign T_1379 = T_1378[2:0];
  assign GEN_45 = T_1374 ? io_chosen : T_1344;
  assign GEN_46 = T_1374 ? T_1379 : T_1342;
  assign GEN_47 = T_1346 ? T_1344 : choice;
  assign GEN_48 = T_1373 ? io_chosen : lastGrant;
  assign T_1384 = GEN_57 > lastGrant;
  assign T_1386 = GEN_58 > lastGrant;
  assign T_1388 = GEN_59 > lastGrant;
  assign T_1390 = 3'h4 > lastGrant;
  assign T_1392 = io_in_1_valid & T_1384;
  assign T_1393 = io_in_2_valid & T_1386;
  assign T_1394 = io_in_3_valid & T_1388;
  assign T_1395 = io_in_4_valid & T_1390;
  assign T_1398 = T_1392 | T_1393;
  assign T_1399 = T_1398 | T_1394;
  assign T_1400 = T_1399 | T_1395;
  assign T_1401 = T_1400 | io_in_0_valid;
  assign T_1402 = T_1401 | io_in_1_valid;
  assign T_1403 = T_1402 | io_in_2_valid;
  assign T_1404 = T_1403 | io_in_3_valid;
  assign T_1408 = T_1392 == 1'h0;
  assign T_1410 = T_1398 == 1'h0;
  assign T_1412 = T_1399 == 1'h0;
  assign T_1414 = T_1400 == 1'h0;
  assign T_1416 = T_1401 == 1'h0;
  assign T_1418 = T_1402 == 1'h0;
  assign T_1420 = T_1403 == 1'h0;
  assign T_1422 = T_1404 == 1'h0;
  assign T_1426 = T_1384 | T_1416;
  assign T_1427 = T_1408 & T_1386;
  assign T_1428 = T_1427 | T_1418;
  assign T_1429 = T_1410 & T_1388;
  assign T_1430 = T_1429 | T_1420;
  assign T_1431 = T_1412 & T_1390;
  assign T_1432 = T_1431 | T_1422;
  assign T_1434 = T_1344 == GEN_84;
  assign T_1435 = T_1346 ? T_1434 : T_1414;
  assign T_1436 = T_1435 & io_out_ready;
  assign T_1438 = T_1344 == GEN_57;
  assign T_1439 = T_1346 ? T_1438 : T_1426;
  assign T_1440 = T_1439 & io_out_ready;
  assign T_1442 = T_1344 == GEN_58;
  assign T_1443 = T_1346 ? T_1442 : T_1428;
  assign T_1444 = T_1443 & io_out_ready;
  assign T_1446 = T_1344 == GEN_59;
  assign T_1447 = T_1346 ? T_1446 : T_1430;
  assign T_1448 = T_1447 & io_out_ready;
  assign T_1450 = T_1344 == 3'h4;
  assign T_1451 = T_1346 ? T_1450 : T_1432;
  assign T_1452 = T_1451 & io_out_ready;
  assign GEN_49 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_50 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_50;
  assign GEN_52 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_51;
  assign GEN_53 = T_1395 ? 3'h4 : GEN_52;
  assign GEN_54 = T_1394 ? {{1'd0}, 2'h3} : GEN_53;
  assign GEN_55 = T_1393 ? {{1'd0}, 2'h2} : GEN_54;
  assign GEN_56 = T_1392 ? {{2'd0}, 1'h1} : GEN_55;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_60 = {1{$random}};
  T_1342 = GEN_60[2:0];
  GEN_61 = {1{$random}};
  T_1344 = GEN_61[2:0];
  GEN_62 = {1{$random}};
  lastGrant = GEN_62[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1342 <= 3'h0;
    end else begin
      T_1342 <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      T_1344 <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_48;
    end
  end
endmodule
module BasicBus_24(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_addr_beat,
  input  [1:0] io_in_0_bits_payload_client_xact_id,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  input   io_in_0_bits_payload_is_builtin_type,
  input  [3:0] io_in_0_bits_payload_g_type,
  input  [63:0] io_in_0_bits_payload_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_addr_beat,
  input  [1:0] io_in_1_bits_payload_client_xact_id,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  input   io_in_1_bits_payload_is_builtin_type,
  input  [3:0] io_in_1_bits_payload_g_type,
  input  [63:0] io_in_1_bits_payload_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_addr_beat,
  input  [1:0] io_in_2_bits_payload_client_xact_id,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  input   io_in_2_bits_payload_is_builtin_type,
  input  [3:0] io_in_2_bits_payload_g_type,
  input  [63:0] io_in_2_bits_payload_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_addr_beat,
  input  [1:0] io_in_3_bits_payload_client_xact_id,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  input   io_in_3_bits_payload_is_builtin_type,
  input  [3:0] io_in_3_bits_payload_g_type,
  input  [63:0] io_in_3_bits_payload_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_addr_beat,
  input  [1:0] io_in_4_bits_payload_client_xact_id,
  input  [2:0] io_in_4_bits_payload_manager_xact_id,
  input   io_in_4_bits_payload_is_builtin_type,
  input  [3:0] io_in_4_bits_payload_g_type,
  input  [63:0] io_in_4_bits_payload_data,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [2:0] io_out_0_bits_header_src,
  output [2:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_addr_beat,
  output [1:0] io_out_0_bits_payload_client_xact_id,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  output  io_out_0_bits_payload_is_builtin_type,
  output [3:0] io_out_0_bits_payload_g_type,
  output [63:0] io_out_0_bits_payload_data,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [2:0] io_out_1_bits_header_src,
  output [2:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_addr_beat,
  output [1:0] io_out_1_bits_payload_client_xact_id,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  output  io_out_1_bits_payload_is_builtin_type,
  output [3:0] io_out_1_bits_payload_g_type,
  output [63:0] io_out_1_bits_payload_data,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [2:0] io_out_2_bits_header_src,
  output [2:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_addr_beat,
  output [1:0] io_out_2_bits_payload_client_xact_id,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  output  io_out_2_bits_payload_is_builtin_type,
  output [3:0] io_out_2_bits_payload_g_type,
  output [63:0] io_out_2_bits_payload_data,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [2:0] io_out_3_bits_header_src,
  output [2:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_addr_beat,
  output [1:0] io_out_3_bits_payload_client_xact_id,
  output [2:0] io_out_3_bits_payload_manager_xact_id,
  output  io_out_3_bits_payload_is_builtin_type,
  output [3:0] io_out_3_bits_payload_g_type,
  output [63:0] io_out_3_bits_payload_data,
  input   io_out_4_ready,
  output  io_out_4_valid,
  output [2:0] io_out_4_bits_header_src,
  output [2:0] io_out_4_bits_header_dst,
  output [2:0] io_out_4_bits_payload_addr_beat,
  output [1:0] io_out_4_bits_payload_client_xact_id,
  output [2:0] io_out_4_bits_payload_manager_xact_id,
  output  io_out_4_bits_payload_is_builtin_type,
  output [3:0] io_out_4_bits_payload_g_type,
  output [63:0] io_out_4_bits_payload_data
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [2:0] arb_io_in_0_bits_header_src;
  wire [2:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_addr_beat;
  wire [1:0] arb_io_in_0_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_0_bits_payload_g_type;
  wire [63:0] arb_io_in_0_bits_payload_data;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [2:0] arb_io_in_1_bits_header_src;
  wire [2:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_addr_beat;
  wire [1:0] arb_io_in_1_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_1_bits_payload_g_type;
  wire [63:0] arb_io_in_1_bits_payload_data;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [2:0] arb_io_in_2_bits_header_src;
  wire [2:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_addr_beat;
  wire [1:0] arb_io_in_2_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_2_bits_payload_g_type;
  wire [63:0] arb_io_in_2_bits_payload_data;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [2:0] arb_io_in_3_bits_header_src;
  wire [2:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_addr_beat;
  wire [1:0] arb_io_in_3_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_3_bits_payload_g_type;
  wire [63:0] arb_io_in_3_bits_payload_data;
  wire  arb_io_in_4_ready;
  wire  arb_io_in_4_valid;
  wire [2:0] arb_io_in_4_bits_header_src;
  wire [2:0] arb_io_in_4_bits_header_dst;
  wire [2:0] arb_io_in_4_bits_payload_addr_beat;
  wire [1:0] arb_io_in_4_bits_payload_client_xact_id;
  wire [2:0] arb_io_in_4_bits_payload_manager_xact_id;
  wire  arb_io_in_4_bits_payload_is_builtin_type;
  wire [3:0] arb_io_in_4_bits_payload_g_type;
  wire [63:0] arb_io_in_4_bits_payload_data;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [2:0] arb_io_out_bits_header_src;
  wire [2:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_addr_beat;
  wire [1:0] arb_io_out_bits_payload_client_xact_id;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire  arb_io_out_bits_payload_is_builtin_type;
  wire [3:0] arb_io_out_bits_payload_g_type;
  wire [63:0] arb_io_out_bits_payload_data;
  wire [2:0] arb_io_chosen;
  wire  GEN_0;
  wire [2:0] GEN_5;
  wire  GEN_1;
  wire [2:0] GEN_6;
  wire  GEN_2;
  wire [2:0] GEN_7;
  wire  GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_8;
  wire  T_1831;
  wire  T_1832;
  wire  T_1834;
  wire  T_1835;
  wire  T_1837;
  wire  T_1838;
  wire  T_1840;
  wire  T_1841;
  wire  T_1843;
  wire  T_1844;
  LockingRRArbiter_25 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(arb_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(arb_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(arb_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(arb_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(arb_io_in_0_bits_payload_data),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(arb_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(arb_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(arb_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(arb_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(arb_io_in_1_bits_payload_data),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(arb_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(arb_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(arb_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(arb_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(arb_io_in_2_bits_payload_data),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(arb_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(arb_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(arb_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(arb_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(arb_io_in_3_bits_payload_data),
    .io_in_4_ready(arb_io_in_4_ready),
    .io_in_4_valid(arb_io_in_4_valid),
    .io_in_4_bits_header_src(arb_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(arb_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_beat(arb_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_client_xact_id(arb_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_manager_xact_id(arb_io_in_4_bits_payload_manager_xact_id),
    .io_in_4_bits_payload_is_builtin_type(arb_io_in_4_bits_payload_is_builtin_type),
    .io_in_4_bits_payload_g_type(arb_io_in_4_bits_payload_g_type),
    .io_in_4_bits_payload_data(arb_io_in_4_bits_payload_data),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_addr_beat(arb_io_out_bits_payload_addr_beat),
    .io_out_bits_payload_client_xact_id(arb_io_out_bits_payload_client_xact_id),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_out_bits_payload_is_builtin_type(arb_io_out_bits_payload_is_builtin_type),
    .io_out_bits_payload_g_type(arb_io_out_bits_payload_g_type),
    .io_out_bits_payload_data(arb_io_out_bits_payload_data),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_in_4_ready = arb_io_in_4_ready;
  assign io_out_0_valid = T_1832;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_0_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_0_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_0_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_0_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_1_valid = T_1835;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_1_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_1_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_1_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_2_valid = T_1838;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_2_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_2_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_2_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_3_valid = T_1841;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_3_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_3_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_3_bits_payload_data = arb_io_out_bits_payload_data;
  assign io_out_4_valid = T_1844;
  assign io_out_4_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_4_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_4_bits_payload_addr_beat = arb_io_out_bits_payload_addr_beat;
  assign io_out_4_bits_payload_client_xact_id = arb_io_out_bits_payload_client_xact_id;
  assign io_out_4_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_4_bits_payload_is_builtin_type = arb_io_out_bits_payload_is_builtin_type;
  assign io_out_4_bits_payload_g_type = arb_io_out_bits_payload_g_type;
  assign io_out_4_bits_payload_data = arb_io_out_bits_payload_data;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_addr_beat = io_in_0_bits_payload_addr_beat;
  assign arb_io_in_0_bits_payload_client_xact_id = io_in_0_bits_payload_client_xact_id;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_0_bits_payload_is_builtin_type = io_in_0_bits_payload_is_builtin_type;
  assign arb_io_in_0_bits_payload_g_type = io_in_0_bits_payload_g_type;
  assign arb_io_in_0_bits_payload_data = io_in_0_bits_payload_data;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_addr_beat = io_in_1_bits_payload_addr_beat;
  assign arb_io_in_1_bits_payload_client_xact_id = io_in_1_bits_payload_client_xact_id;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_1_bits_payload_is_builtin_type = io_in_1_bits_payload_is_builtin_type;
  assign arb_io_in_1_bits_payload_g_type = io_in_1_bits_payload_g_type;
  assign arb_io_in_1_bits_payload_data = io_in_1_bits_payload_data;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_addr_beat = io_in_2_bits_payload_addr_beat;
  assign arb_io_in_2_bits_payload_client_xact_id = io_in_2_bits_payload_client_xact_id;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_2_bits_payload_is_builtin_type = io_in_2_bits_payload_is_builtin_type;
  assign arb_io_in_2_bits_payload_g_type = io_in_2_bits_payload_g_type;
  assign arb_io_in_2_bits_payload_data = io_in_2_bits_payload_data;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_addr_beat = io_in_3_bits_payload_addr_beat;
  assign arb_io_in_3_bits_payload_client_xact_id = io_in_3_bits_payload_client_xact_id;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_3_bits_payload_is_builtin_type = io_in_3_bits_payload_is_builtin_type;
  assign arb_io_in_3_bits_payload_g_type = io_in_3_bits_payload_g_type;
  assign arb_io_in_3_bits_payload_data = io_in_3_bits_payload_data;
  assign arb_io_in_4_valid = io_in_4_valid;
  assign arb_io_in_4_bits_header_src = io_in_4_bits_header_src;
  assign arb_io_in_4_bits_header_dst = io_in_4_bits_header_dst;
  assign arb_io_in_4_bits_payload_addr_beat = io_in_4_bits_payload_addr_beat;
  assign arb_io_in_4_bits_payload_client_xact_id = io_in_4_bits_payload_client_xact_id;
  assign arb_io_in_4_bits_payload_manager_xact_id = io_in_4_bits_payload_manager_xact_id;
  assign arb_io_in_4_bits_payload_is_builtin_type = io_in_4_bits_payload_is_builtin_type;
  assign arb_io_in_4_bits_payload_g_type = io_in_4_bits_payload_g_type;
  assign arb_io_in_4_bits_payload_data = io_in_4_bits_payload_data;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_4;
  assign GEN_5 = {{2'd0}, 1'h1};
  assign GEN_1 = GEN_5 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_6 = {{1'd0}, 2'h2};
  assign GEN_2 = GEN_6 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = {{1'd0}, 2'h3};
  assign GEN_3 = GEN_7 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_4 = 3'h4 == arb_io_out_bits_header_dst ? io_out_4_ready : GEN_3;
  assign GEN_8 = {{2'd0}, 1'h0};
  assign T_1831 = arb_io_out_bits_header_dst == GEN_8;
  assign T_1832 = arb_io_out_valid & T_1831;
  assign T_1834 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1835 = arb_io_out_valid & T_1834;
  assign T_1837 = arb_io_out_bits_header_dst == GEN_6;
  assign T_1838 = arb_io_out_valid & T_1837;
  assign T_1840 = arb_io_out_bits_header_dst == GEN_7;
  assign T_1841 = arb_io_out_valid & T_1840;
  assign T_1843 = arb_io_out_bits_header_dst == 3'h4;
  assign T_1844 = arb_io_out_valid & T_1843;
endmodule
module LockingRRArbiter_27(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_manager_xact_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_header_src,
  output [2:0] io_out_bits_header_dst,
  output [2:0] io_out_bits_payload_manager_xact_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_29;
  wire  GEN_4;
  wire [2:0] GEN_30;
  wire  GEN_5;
  wire [2:0] GEN_31;
  wire  GEN_6;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [2:0] GEN_9;
  wire [2:0] GEN_10;
  wire [2:0] GEN_11;
  wire [2:0] GEN_2;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [2:0] GEN_3;
  wire [2:0] GEN_16;
  wire [2:0] GEN_17;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire  T_1152;
  reg [2:0] lastGrant;
  reg [31:0] GEN_32;
  wire [2:0] GEN_20;
  wire  T_1155;
  wire  T_1157;
  wire  T_1159;
  wire  T_1161;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1166;
  wire  T_1169;
  wire  T_1170;
  wire  T_1171;
  wire  T_1172;
  wire  T_1173;
  wire  T_1174;
  wire  T_1175;
  wire  T_1179;
  wire  T_1181;
  wire  T_1183;
  wire  T_1185;
  wire  T_1187;
  wire  T_1189;
  wire  T_1191;
  wire  T_1193;
  wire  T_1197;
  wire  T_1198;
  wire  T_1199;
  wire  T_1200;
  wire  T_1201;
  wire  T_1202;
  wire  T_1203;
  wire  T_1204;
  wire  T_1205;
  wire  T_1206;
  wire  T_1207;
  wire  T_1208;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire [2:0] GEN_28;
  assign io_in_0_ready = T_1204;
  assign io_in_1_ready = T_1205;
  assign io_in_2_ready = T_1206;
  assign io_in_3_ready = T_1207;
  assign io_in_4_ready = T_1208;
  assign io_out_valid = GEN_0;
  assign io_out_bits_header_src = GEN_1;
  assign io_out_bits_header_dst = GEN_2;
  assign io_out_bits_payload_manager_xact_id = GEN_3;
  assign io_chosen = choice;
  assign choice = GEN_28;
  assign GEN_0 = GEN_7;
  assign GEN_29 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_29 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_30 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_30 == io_chosen ? io_in_2_valid : GEN_4;
  assign GEN_31 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_31 == io_chosen ? io_in_3_valid : GEN_5;
  assign GEN_7 = 3'h4 == io_chosen ? io_in_4_valid : GEN_6;
  assign GEN_1 = GEN_11;
  assign GEN_8 = GEN_29 == io_chosen ? io_in_1_bits_header_src : io_in_0_bits_header_src;
  assign GEN_9 = GEN_30 == io_chosen ? io_in_2_bits_header_src : GEN_8;
  assign GEN_10 = GEN_31 == io_chosen ? io_in_3_bits_header_src : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_bits_header_src : GEN_10;
  assign GEN_2 = GEN_15;
  assign GEN_12 = GEN_29 == io_chosen ? io_in_1_bits_header_dst : io_in_0_bits_header_dst;
  assign GEN_13 = GEN_30 == io_chosen ? io_in_2_bits_header_dst : GEN_12;
  assign GEN_14 = GEN_31 == io_chosen ? io_in_3_bits_header_dst : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_header_dst : GEN_14;
  assign GEN_3 = GEN_19;
  assign GEN_16 = GEN_29 == io_chosen ? io_in_1_bits_payload_manager_xact_id : io_in_0_bits_payload_manager_xact_id;
  assign GEN_17 = GEN_30 == io_chosen ? io_in_2_bits_payload_manager_xact_id : GEN_16;
  assign GEN_18 = GEN_31 == io_chosen ? io_in_3_bits_payload_manager_xact_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_payload_manager_xact_id : GEN_18;
  assign T_1152 = io_out_ready & io_out_valid;
  assign GEN_20 = T_1152 ? io_chosen : lastGrant;
  assign T_1155 = GEN_29 > lastGrant;
  assign T_1157 = GEN_30 > lastGrant;
  assign T_1159 = GEN_31 > lastGrant;
  assign T_1161 = 3'h4 > lastGrant;
  assign T_1163 = io_in_1_valid & T_1155;
  assign T_1164 = io_in_2_valid & T_1157;
  assign T_1165 = io_in_3_valid & T_1159;
  assign T_1166 = io_in_4_valid & T_1161;
  assign T_1169 = T_1163 | T_1164;
  assign T_1170 = T_1169 | T_1165;
  assign T_1171 = T_1170 | T_1166;
  assign T_1172 = T_1171 | io_in_0_valid;
  assign T_1173 = T_1172 | io_in_1_valid;
  assign T_1174 = T_1173 | io_in_2_valid;
  assign T_1175 = T_1174 | io_in_3_valid;
  assign T_1179 = T_1163 == 1'h0;
  assign T_1181 = T_1169 == 1'h0;
  assign T_1183 = T_1170 == 1'h0;
  assign T_1185 = T_1171 == 1'h0;
  assign T_1187 = T_1172 == 1'h0;
  assign T_1189 = T_1173 == 1'h0;
  assign T_1191 = T_1174 == 1'h0;
  assign T_1193 = T_1175 == 1'h0;
  assign T_1197 = T_1155 | T_1187;
  assign T_1198 = T_1179 & T_1157;
  assign T_1199 = T_1198 | T_1189;
  assign T_1200 = T_1181 & T_1159;
  assign T_1201 = T_1200 | T_1191;
  assign T_1202 = T_1183 & T_1161;
  assign T_1203 = T_1202 | T_1193;
  assign T_1204 = T_1185 & io_out_ready;
  assign T_1205 = T_1197 & io_out_ready;
  assign T_1206 = T_1199 & io_out_ready;
  assign T_1207 = T_1201 & io_out_ready;
  assign T_1208 = T_1203 & io_out_ready;
  assign GEN_21 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_22 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_21;
  assign GEN_23 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_22;
  assign GEN_24 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_23;
  assign GEN_25 = T_1166 ? 3'h4 : GEN_24;
  assign GEN_26 = T_1165 ? {{1'd0}, 2'h3} : GEN_25;
  assign GEN_27 = T_1164 ? {{1'd0}, 2'h2} : GEN_26;
  assign GEN_28 = T_1163 ? {{2'd0}, 1'h1} : GEN_27;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_32 = {1{$random}};
  lastGrant = GEN_32[2:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_20;
    end
  end
endmodule
module BasicBus_26(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_header_src,
  input  [2:0] io_in_0_bits_header_dst,
  input  [2:0] io_in_0_bits_payload_manager_xact_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_header_src,
  input  [2:0] io_in_1_bits_header_dst,
  input  [2:0] io_in_1_bits_payload_manager_xact_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_header_src,
  input  [2:0] io_in_2_bits_header_dst,
  input  [2:0] io_in_2_bits_payload_manager_xact_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_header_src,
  input  [2:0] io_in_3_bits_header_dst,
  input  [2:0] io_in_3_bits_payload_manager_xact_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_header_src,
  input  [2:0] io_in_4_bits_header_dst,
  input  [2:0] io_in_4_bits_payload_manager_xact_id,
  input   io_out_0_ready,
  output  io_out_0_valid,
  output [2:0] io_out_0_bits_header_src,
  output [2:0] io_out_0_bits_header_dst,
  output [2:0] io_out_0_bits_payload_manager_xact_id,
  input   io_out_1_ready,
  output  io_out_1_valid,
  output [2:0] io_out_1_bits_header_src,
  output [2:0] io_out_1_bits_header_dst,
  output [2:0] io_out_1_bits_payload_manager_xact_id,
  input   io_out_2_ready,
  output  io_out_2_valid,
  output [2:0] io_out_2_bits_header_src,
  output [2:0] io_out_2_bits_header_dst,
  output [2:0] io_out_2_bits_payload_manager_xact_id,
  input   io_out_3_ready,
  output  io_out_3_valid,
  output [2:0] io_out_3_bits_header_src,
  output [2:0] io_out_3_bits_header_dst,
  output [2:0] io_out_3_bits_payload_manager_xact_id,
  input   io_out_4_ready,
  output  io_out_4_valid,
  output [2:0] io_out_4_bits_header_src,
  output [2:0] io_out_4_bits_header_dst,
  output [2:0] io_out_4_bits_payload_manager_xact_id
);
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [2:0] arb_io_in_0_bits_header_src;
  wire [2:0] arb_io_in_0_bits_header_dst;
  wire [2:0] arb_io_in_0_bits_payload_manager_xact_id;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [2:0] arb_io_in_1_bits_header_src;
  wire [2:0] arb_io_in_1_bits_header_dst;
  wire [2:0] arb_io_in_1_bits_payload_manager_xact_id;
  wire  arb_io_in_2_ready;
  wire  arb_io_in_2_valid;
  wire [2:0] arb_io_in_2_bits_header_src;
  wire [2:0] arb_io_in_2_bits_header_dst;
  wire [2:0] arb_io_in_2_bits_payload_manager_xact_id;
  wire  arb_io_in_3_ready;
  wire  arb_io_in_3_valid;
  wire [2:0] arb_io_in_3_bits_header_src;
  wire [2:0] arb_io_in_3_bits_header_dst;
  wire [2:0] arb_io_in_3_bits_payload_manager_xact_id;
  wire  arb_io_in_4_ready;
  wire  arb_io_in_4_valid;
  wire [2:0] arb_io_in_4_bits_header_src;
  wire [2:0] arb_io_in_4_bits_header_dst;
  wire [2:0] arb_io_in_4_bits_payload_manager_xact_id;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [2:0] arb_io_out_bits_header_src;
  wire [2:0] arb_io_out_bits_header_dst;
  wire [2:0] arb_io_out_bits_payload_manager_xact_id;
  wire [2:0] arb_io_chosen;
  wire  GEN_0;
  wire [2:0] GEN_5;
  wire  GEN_1;
  wire [2:0] GEN_6;
  wire  GEN_2;
  wire [2:0] GEN_7;
  wire  GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_8;
  wire  T_1571;
  wire  T_1572;
  wire  T_1574;
  wire  T_1575;
  wire  T_1577;
  wire  T_1578;
  wire  T_1580;
  wire  T_1581;
  wire  T_1583;
  wire  T_1584;
  LockingRRArbiter_27 arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_header_src(arb_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(arb_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(arb_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_header_src(arb_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(arb_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(arb_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(arb_io_in_2_ready),
    .io_in_2_valid(arb_io_in_2_valid),
    .io_in_2_bits_header_src(arb_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(arb_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(arb_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(arb_io_in_3_ready),
    .io_in_3_valid(arb_io_in_3_valid),
    .io_in_3_bits_header_src(arb_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(arb_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(arb_io_in_3_bits_payload_manager_xact_id),
    .io_in_4_ready(arb_io_in_4_ready),
    .io_in_4_valid(arb_io_in_4_valid),
    .io_in_4_bits_header_src(arb_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(arb_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_manager_xact_id(arb_io_in_4_bits_payload_manager_xact_id),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_header_src(arb_io_out_bits_header_src),
    .io_out_bits_header_dst(arb_io_out_bits_header_dst),
    .io_out_bits_payload_manager_xact_id(arb_io_out_bits_payload_manager_xact_id),
    .io_chosen(arb_io_chosen)
  );
  assign io_in_0_ready = arb_io_in_0_ready;
  assign io_in_1_ready = arb_io_in_1_ready;
  assign io_in_2_ready = arb_io_in_2_ready;
  assign io_in_3_ready = arb_io_in_3_ready;
  assign io_in_4_ready = arb_io_in_4_ready;
  assign io_out_0_valid = T_1572;
  assign io_out_0_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_0_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_0_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_1_valid = T_1575;
  assign io_out_1_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_1_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_1_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_2_valid = T_1578;
  assign io_out_2_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_2_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_2_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_3_valid = T_1581;
  assign io_out_3_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_3_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_3_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign io_out_4_valid = T_1584;
  assign io_out_4_bits_header_src = arb_io_out_bits_header_src;
  assign io_out_4_bits_header_dst = arb_io_out_bits_header_dst;
  assign io_out_4_bits_payload_manager_xact_id = arb_io_out_bits_payload_manager_xact_id;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_in_0_valid;
  assign arb_io_in_0_bits_header_src = io_in_0_bits_header_src;
  assign arb_io_in_0_bits_header_dst = io_in_0_bits_header_dst;
  assign arb_io_in_0_bits_payload_manager_xact_id = io_in_0_bits_payload_manager_xact_id;
  assign arb_io_in_1_valid = io_in_1_valid;
  assign arb_io_in_1_bits_header_src = io_in_1_bits_header_src;
  assign arb_io_in_1_bits_header_dst = io_in_1_bits_header_dst;
  assign arb_io_in_1_bits_payload_manager_xact_id = io_in_1_bits_payload_manager_xact_id;
  assign arb_io_in_2_valid = io_in_2_valid;
  assign arb_io_in_2_bits_header_src = io_in_2_bits_header_src;
  assign arb_io_in_2_bits_header_dst = io_in_2_bits_header_dst;
  assign arb_io_in_2_bits_payload_manager_xact_id = io_in_2_bits_payload_manager_xact_id;
  assign arb_io_in_3_valid = io_in_3_valid;
  assign arb_io_in_3_bits_header_src = io_in_3_bits_header_src;
  assign arb_io_in_3_bits_header_dst = io_in_3_bits_header_dst;
  assign arb_io_in_3_bits_payload_manager_xact_id = io_in_3_bits_payload_manager_xact_id;
  assign arb_io_in_4_valid = io_in_4_valid;
  assign arb_io_in_4_bits_header_src = io_in_4_bits_header_src;
  assign arb_io_in_4_bits_header_dst = io_in_4_bits_header_dst;
  assign arb_io_in_4_bits_payload_manager_xact_id = io_in_4_bits_payload_manager_xact_id;
  assign arb_io_out_ready = GEN_0;
  assign GEN_0 = GEN_4;
  assign GEN_5 = {{2'd0}, 1'h1};
  assign GEN_1 = GEN_5 == arb_io_out_bits_header_dst ? io_out_1_ready : io_out_0_ready;
  assign GEN_6 = {{1'd0}, 2'h2};
  assign GEN_2 = GEN_6 == arb_io_out_bits_header_dst ? io_out_2_ready : GEN_1;
  assign GEN_7 = {{1'd0}, 2'h3};
  assign GEN_3 = GEN_7 == arb_io_out_bits_header_dst ? io_out_3_ready : GEN_2;
  assign GEN_4 = 3'h4 == arb_io_out_bits_header_dst ? io_out_4_ready : GEN_3;
  assign GEN_8 = {{2'd0}, 1'h0};
  assign T_1571 = arb_io_out_bits_header_dst == GEN_8;
  assign T_1572 = arb_io_out_valid & T_1571;
  assign T_1574 = arb_io_out_bits_header_dst == GEN_5;
  assign T_1575 = arb_io_out_valid & T_1574;
  assign T_1577 = arb_io_out_bits_header_dst == GEN_6;
  assign T_1578 = arb_io_out_valid & T_1577;
  assign T_1580 = arb_io_out_bits_header_dst == GEN_7;
  assign T_1581 = arb_io_out_valid & T_1580;
  assign T_1583 = arb_io_out_bits_header_dst == 3'h4;
  assign T_1584 = arb_io_out_valid & T_1583;
endmodule
module PortedTileLinkCrossbar(
  input   clk,
  input   reset,
  output  io_clients_cached_0_acquire_ready,
  input   io_clients_cached_0_acquire_valid,
  input  [25:0] io_clients_cached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_cached_0_acquire_bits_addr_beat,
  input   io_clients_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_cached_0_acquire_bits_a_type,
  input  [11:0] io_clients_cached_0_acquire_bits_union,
  input  [63:0] io_clients_cached_0_acquire_bits_data,
  input   io_clients_cached_0_probe_ready,
  output  io_clients_cached_0_probe_valid,
  output [25:0] io_clients_cached_0_probe_bits_addr_block,
  output [1:0] io_clients_cached_0_probe_bits_p_type,
  output  io_clients_cached_0_release_ready,
  input   io_clients_cached_0_release_valid,
  input  [2:0] io_clients_cached_0_release_bits_addr_beat,
  input  [25:0] io_clients_cached_0_release_bits_addr_block,
  input  [1:0] io_clients_cached_0_release_bits_client_xact_id,
  input   io_clients_cached_0_release_bits_voluntary,
  input  [2:0] io_clients_cached_0_release_bits_r_type,
  input  [63:0] io_clients_cached_0_release_bits_data,
  input   io_clients_cached_0_grant_ready,
  output  io_clients_cached_0_grant_valid,
  output [2:0] io_clients_cached_0_grant_bits_addr_beat,
  output [1:0] io_clients_cached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_cached_0_grant_bits_manager_xact_id,
  output  io_clients_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_cached_0_grant_bits_g_type,
  output [63:0] io_clients_cached_0_grant_bits_data,
  output  io_clients_cached_0_grant_bits_manager_id,
  output  io_clients_cached_0_finish_ready,
  input   io_clients_cached_0_finish_valid,
  input  [2:0] io_clients_cached_0_finish_bits_manager_xact_id,
  input   io_clients_cached_0_finish_bits_manager_id,
  output  io_clients_uncached_0_acquire_ready,
  input   io_clients_uncached_0_acquire_valid,
  input  [25:0] io_clients_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_clients_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_0_acquire_bits_addr_beat,
  input   io_clients_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_0_acquire_bits_a_type,
  input  [11:0] io_clients_uncached_0_acquire_bits_union,
  input  [63:0] io_clients_uncached_0_acquire_bits_data,
  input   io_clients_uncached_0_grant_ready,
  output  io_clients_uncached_0_grant_valid,
  output [2:0] io_clients_uncached_0_grant_bits_addr_beat,
  output [1:0] io_clients_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_clients_uncached_0_grant_bits_manager_xact_id,
  output  io_clients_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_0_grant_bits_g_type,
  output [63:0] io_clients_uncached_0_grant_bits_data,
  output  io_clients_uncached_1_acquire_ready,
  input   io_clients_uncached_1_acquire_valid,
  input  [25:0] io_clients_uncached_1_acquire_bits_addr_block,
  input  [1:0] io_clients_uncached_1_acquire_bits_client_xact_id,
  input  [2:0] io_clients_uncached_1_acquire_bits_addr_beat,
  input   io_clients_uncached_1_acquire_bits_is_builtin_type,
  input  [2:0] io_clients_uncached_1_acquire_bits_a_type,
  input  [11:0] io_clients_uncached_1_acquire_bits_union,
  input  [63:0] io_clients_uncached_1_acquire_bits_data,
  input   io_clients_uncached_1_grant_ready,
  output  io_clients_uncached_1_grant_valid,
  output [2:0] io_clients_uncached_1_grant_bits_addr_beat,
  output [1:0] io_clients_uncached_1_grant_bits_client_xact_id,
  output [2:0] io_clients_uncached_1_grant_bits_manager_xact_id,
  output  io_clients_uncached_1_grant_bits_is_builtin_type,
  output [3:0] io_clients_uncached_1_grant_bits_g_type,
  output [63:0] io_clients_uncached_1_grant_bits_data,
  input   io_managers_0_acquire_ready,
  output  io_managers_0_acquire_valid,
  output [25:0] io_managers_0_acquire_bits_addr_block,
  output [1:0] io_managers_0_acquire_bits_client_xact_id,
  output [2:0] io_managers_0_acquire_bits_addr_beat,
  output  io_managers_0_acquire_bits_is_builtin_type,
  output [2:0] io_managers_0_acquire_bits_a_type,
  output [11:0] io_managers_0_acquire_bits_union,
  output [63:0] io_managers_0_acquire_bits_data,
  output [1:0] io_managers_0_acquire_bits_client_id,
  output  io_managers_0_grant_ready,
  input   io_managers_0_grant_valid,
  input  [2:0] io_managers_0_grant_bits_addr_beat,
  input  [1:0] io_managers_0_grant_bits_client_xact_id,
  input  [2:0] io_managers_0_grant_bits_manager_xact_id,
  input   io_managers_0_grant_bits_is_builtin_type,
  input  [3:0] io_managers_0_grant_bits_g_type,
  input  [63:0] io_managers_0_grant_bits_data,
  input  [1:0] io_managers_0_grant_bits_client_id,
  input   io_managers_0_finish_ready,
  output  io_managers_0_finish_valid,
  output [2:0] io_managers_0_finish_bits_manager_xact_id,
  output  io_managers_0_probe_ready,
  input   io_managers_0_probe_valid,
  input  [25:0] io_managers_0_probe_bits_addr_block,
  input  [1:0] io_managers_0_probe_bits_p_type,
  input  [1:0] io_managers_0_probe_bits_client_id,
  input   io_managers_0_release_ready,
  output  io_managers_0_release_valid,
  output [2:0] io_managers_0_release_bits_addr_beat,
  output [25:0] io_managers_0_release_bits_addr_block,
  output [1:0] io_managers_0_release_bits_client_xact_id,
  output  io_managers_0_release_bits_voluntary,
  output [2:0] io_managers_0_release_bits_r_type,
  output [63:0] io_managers_0_release_bits_data,
  output [1:0] io_managers_0_release_bits_client_id,
  input   io_managers_1_acquire_ready,
  output  io_managers_1_acquire_valid,
  output [25:0] io_managers_1_acquire_bits_addr_block,
  output [1:0] io_managers_1_acquire_bits_client_xact_id,
  output [2:0] io_managers_1_acquire_bits_addr_beat,
  output  io_managers_1_acquire_bits_is_builtin_type,
  output [2:0] io_managers_1_acquire_bits_a_type,
  output [11:0] io_managers_1_acquire_bits_union,
  output [63:0] io_managers_1_acquire_bits_data,
  output [1:0] io_managers_1_acquire_bits_client_id,
  output  io_managers_1_grant_ready,
  input   io_managers_1_grant_valid,
  input  [2:0] io_managers_1_grant_bits_addr_beat,
  input  [1:0] io_managers_1_grant_bits_client_xact_id,
  input  [2:0] io_managers_1_grant_bits_manager_xact_id,
  input   io_managers_1_grant_bits_is_builtin_type,
  input  [3:0] io_managers_1_grant_bits_g_type,
  input  [63:0] io_managers_1_grant_bits_data,
  input  [1:0] io_managers_1_grant_bits_client_id,
  input   io_managers_1_finish_ready,
  output  io_managers_1_finish_valid,
  output [2:0] io_managers_1_finish_bits_manager_xact_id,
  output  io_managers_1_probe_ready,
  input   io_managers_1_probe_valid,
  input  [25:0] io_managers_1_probe_bits_addr_block,
  input  [1:0] io_managers_1_probe_bits_p_type,
  input  [1:0] io_managers_1_probe_bits_client_id,
  input   io_managers_1_release_ready,
  output  io_managers_1_release_valid,
  output [2:0] io_managers_1_release_bits_addr_beat,
  output [25:0] io_managers_1_release_bits_addr_block,
  output [1:0] io_managers_1_release_bits_client_xact_id,
  output  io_managers_1_release_bits_voluntary,
  output [2:0] io_managers_1_release_bits_r_type,
  output [63:0] io_managers_1_release_bits_data,
  output [1:0] io_managers_1_release_bits_client_id
);
  wire  TileLinkEnqueuer_14127_clk;
  wire  TileLinkEnqueuer_14127_reset;
  wire  TileLinkEnqueuer_14127_io_client_acquire_ready;
  wire  TileLinkEnqueuer_14127_io_client_acquire_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_client_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_14127_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_14127_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_14127_io_client_grant_ready;
  wire  TileLinkEnqueuer_14127_io_client_grant_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_client_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_14127_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_14127_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_14127_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_14127_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_14127_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_14127_io_client_finish_ready;
  wire  TileLinkEnqueuer_14127_io_client_finish_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_client_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_14127_io_client_probe_ready;
  wire  TileLinkEnqueuer_14127_io_client_probe_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_client_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_14127_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_14127_io_client_release_ready;
  wire  TileLinkEnqueuer_14127_io_client_release_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_client_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_14127_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_14127_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_14127_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_14127_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_14127_io_manager_acquire_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_14127_io_manager_grant_ready;
  wire  TileLinkEnqueuer_14127_io_manager_grant_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_14127_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_14127_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_14127_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_14127_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_14127_io_manager_finish_ready;
  wire  TileLinkEnqueuer_14127_io_manager_finish_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_14127_io_manager_probe_ready;
  wire  TileLinkEnqueuer_14127_io_manager_probe_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_14127_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_14127_io_manager_release_ready;
  wire  TileLinkEnqueuer_14127_io_manager_release_valid;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_14127_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_14127_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_14127_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_14127_io_manager_release_bits_payload_data;
  wire  ClientTileLinkNetworkPort_14128_clk;
  wire  ClientTileLinkNetworkPort_14128_reset;
  wire  ClientTileLinkNetworkPort_14128_io_client_acquire_ready;
  wire  ClientTileLinkNetworkPort_14128_io_client_acquire_valid;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_beat;
  wire  ClientTileLinkNetworkPort_14128_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_a_type;
  wire [11:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_union;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_client_acquire_bits_data;
  wire  ClientTileLinkNetworkPort_14128_io_client_probe_ready;
  wire  ClientTileLinkNetworkPort_14128_io_client_probe_valid;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_client_probe_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_client_probe_bits_p_type;
  wire  ClientTileLinkNetworkPort_14128_io_client_release_ready;
  wire  ClientTileLinkNetworkPort_14128_io_client_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_client_release_bits_client_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_client_release_bits_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_release_bits_r_type;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_client_release_bits_data;
  wire  ClientTileLinkNetworkPort_14128_io_client_grant_ready;
  wire  ClientTileLinkNetworkPort_14128_io_client_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_grant_bits_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_14128_io_client_grant_bits_g_type;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_client_grant_bits_data;
  wire  ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_id;
  wire  ClientTileLinkNetworkPort_14128_io_client_finish_ready;
  wire  ClientTileLinkNetworkPort_14128_io_client_finish_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_id;
  wire  ClientTileLinkNetworkPort_14128_io_network_acquire_ready;
  wire  ClientTileLinkNetworkPort_14128_io_network_acquire_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_src;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_beat;
  wire  ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_union;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_data;
  wire  ClientTileLinkNetworkPort_14128_io_network_grant_ready;
  wire  ClientTileLinkNetworkPort_14128_io_network_grant_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_src;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_data;
  wire  ClientTileLinkNetworkPort_14128_io_network_finish_ready;
  wire  ClientTileLinkNetworkPort_14128_io_network_finish_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_src;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_network_probe_ready;
  wire  ClientTileLinkNetworkPort_14128_io_network_probe_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_src;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_dst;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_p_type;
  wire  ClientTileLinkNetworkPort_14128_io_network_release_ready;
  wire  ClientTileLinkNetworkPort_14128_io_network_release_valid;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_header_src;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_header_dst;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_client_xact_id;
  wire  ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_r_type;
  wire [63:0] ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_clk;
  wire  TileLinkEnqueuer_4_14129_reset;
  wire  TileLinkEnqueuer_4_14129_io_client_acquire_ready;
  wire  TileLinkEnqueuer_4_14129_io_client_acquire_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_io_client_grant_ready;
  wire  TileLinkEnqueuer_4_14129_io_client_grant_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_io_client_finish_ready;
  wire  TileLinkEnqueuer_4_14129_io_client_finish_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_client_probe_ready;
  wire  TileLinkEnqueuer_4_14129_io_client_probe_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_14129_io_client_release_ready;
  wire  TileLinkEnqueuer_4_14129_io_client_release_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_14129_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_14129_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_4_14129_io_manager_acquire_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_io_manager_grant_ready;
  wire  TileLinkEnqueuer_4_14129_io_manager_grant_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_4_14129_io_manager_finish_ready;
  wire  TileLinkEnqueuer_4_14129_io_manager_finish_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_manager_probe_ready;
  wire  TileLinkEnqueuer_4_14129_io_manager_probe_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_4_14129_io_manager_release_ready;
  wire  TileLinkEnqueuer_4_14129_io_manager_release_valid;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14130_clk;
  wire  ClientUncachedTileLinkNetworkPort_14130_reset;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_finish_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_probe_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_release_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_clk;
  wire  TileLinkEnqueuer_9_14131_reset;
  wire  TileLinkEnqueuer_9_14131_io_client_acquire_ready;
  wire  TileLinkEnqueuer_9_14131_io_client_acquire_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_io_client_grant_ready;
  wire  TileLinkEnqueuer_9_14131_io_client_grant_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_io_client_finish_ready;
  wire  TileLinkEnqueuer_9_14131_io_client_finish_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_client_probe_ready;
  wire  TileLinkEnqueuer_9_14131_io_client_probe_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_9_14131_io_client_release_ready;
  wire  TileLinkEnqueuer_9_14131_io_client_release_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_9_14131_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_9_14131_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_9_14131_io_manager_acquire_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_io_manager_grant_ready;
  wire  TileLinkEnqueuer_9_14131_io_manager_grant_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_9_14131_io_manager_finish_ready;
  wire  TileLinkEnqueuer_9_14131_io_manager_finish_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_manager_probe_ready;
  wire  TileLinkEnqueuer_9_14131_io_manager_probe_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_9_14131_io_manager_release_ready;
  wire  TileLinkEnqueuer_9_14131_io_manager_release_valid;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_clk;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_reset;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_valid;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_data;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_beat;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_a_type;
  wire [11:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_union;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_g_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_data;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_payload_manager_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_dst;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_p_type;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_ready;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_valid;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_src;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_dst;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_beat;
  wire [25:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_block;
  wire [1:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_client_xact_id;
  wire  ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_voluntary;
  wire [2:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_r_type;
  wire [63:0] ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_14133_clk;
  wire  ManagerTileLinkNetworkPort_14133_reset;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_p_type;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_14133_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_network_acquire_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_14133_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_network_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_14133_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_network_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_network_probe_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_14133_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_14133_io_network_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_clk;
  wire  TileLinkEnqueuer_17_14134_reset;
  wire  TileLinkEnqueuer_17_14134_io_client_acquire_ready;
  wire  TileLinkEnqueuer_17_14134_io_client_acquire_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_io_client_grant_ready;
  wire  TileLinkEnqueuer_17_14134_io_client_grant_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_io_client_finish_ready;
  wire  TileLinkEnqueuer_17_14134_io_client_finish_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_client_probe_ready;
  wire  TileLinkEnqueuer_17_14134_io_client_probe_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_17_14134_io_client_release_ready;
  wire  TileLinkEnqueuer_17_14134_io_client_release_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_17_14134_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_17_14134_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_17_14134_io_manager_acquire_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_io_manager_grant_ready;
  wire  TileLinkEnqueuer_17_14134_io_manager_grant_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_17_14134_io_manager_finish_ready;
  wire  TileLinkEnqueuer_17_14134_io_manager_finish_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_manager_probe_ready;
  wire  TileLinkEnqueuer_17_14134_io_manager_probe_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_17_14134_io_manager_release_ready;
  wire  TileLinkEnqueuer_17_14134_io_manager_release_valid;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_18_14135_clk;
  wire  ManagerTileLinkNetworkPort_18_14135_reset;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_valid;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_beat;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_union;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_grant_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_finish_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_finish_bits_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_probe_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_probe_valid;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_p_type;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_client_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_release_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_data;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_acquire_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_acquire_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_beat;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_is_builtin_type;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_a_type;
  wire [11:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_union;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_grant_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_grant_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_addr_beat;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_client_xact_id;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_is_builtin_type;
  wire [3:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_g_type;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_data;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_finish_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_finish_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_payload_manager_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_probe_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_probe_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_dst;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_p_type;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_release_ready;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_release_valid;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_src;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_dst;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_beat;
  wire [25:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_block;
  wire [1:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_client_xact_id;
  wire  ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_voluntary;
  wire [2:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_r_type;
  wire [63:0] ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_clk;
  wire  TileLinkEnqueuer_19_14136_reset;
  wire  TileLinkEnqueuer_19_14136_io_client_acquire_ready;
  wire  TileLinkEnqueuer_19_14136_io_client_acquire_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_io_client_grant_ready;
  wire  TileLinkEnqueuer_19_14136_io_client_grant_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_io_client_finish_ready;
  wire  TileLinkEnqueuer_19_14136_io_client_finish_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_client_probe_ready;
  wire  TileLinkEnqueuer_19_14136_io_client_probe_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_19_14136_io_client_release_ready;
  wire  TileLinkEnqueuer_19_14136_io_client_release_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_client_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_client_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_19_14136_io_client_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_19_14136_io_client_release_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_io_manager_acquire_ready;
  wire  TileLinkEnqueuer_19_14136_io_manager_acquire_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_beat;
  wire  TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_is_builtin_type;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_a_type;
  wire [11:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_union;
  wire [63:0] TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_io_manager_grant_ready;
  wire  TileLinkEnqueuer_19_14136_io_manager_grant_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_addr_beat;
  wire [1:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_client_xact_id;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_is_builtin_type;
  wire [3:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_g_type;
  wire [63:0] TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_data;
  wire  TileLinkEnqueuer_19_14136_io_manager_finish_ready;
  wire  TileLinkEnqueuer_19_14136_io_manager_finish_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_finish_bits_payload_manager_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_manager_probe_ready;
  wire  TileLinkEnqueuer_19_14136_io_manager_probe_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_dst;
  wire [25:0] TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_p_type;
  wire  TileLinkEnqueuer_19_14136_io_manager_release_ready;
  wire  TileLinkEnqueuer_19_14136_io_manager_release_valid;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_header_src;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_header_dst;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_beat;
  wire [25:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_block;
  wire [1:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_client_xact_id;
  wire  TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_voluntary;
  wire [2:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_r_type;
  wire [63:0] TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_data;
  wire  acqNet_clk;
  wire  acqNet_reset;
  wire  acqNet_io_in_0_ready;
  wire  acqNet_io_in_0_valid;
  wire [2:0] acqNet_io_in_0_bits_header_src;
  wire [2:0] acqNet_io_in_0_bits_header_dst;
  wire [25:0] acqNet_io_in_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_0_bits_payload_addr_beat;
  wire  acqNet_io_in_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_0_bits_payload_a_type;
  wire [11:0] acqNet_io_in_0_bits_payload_union;
  wire [63:0] acqNet_io_in_0_bits_payload_data;
  wire  acqNet_io_in_1_ready;
  wire  acqNet_io_in_1_valid;
  wire [2:0] acqNet_io_in_1_bits_header_src;
  wire [2:0] acqNet_io_in_1_bits_header_dst;
  wire [25:0] acqNet_io_in_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_1_bits_payload_addr_beat;
  wire  acqNet_io_in_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_1_bits_payload_a_type;
  wire [11:0] acqNet_io_in_1_bits_payload_union;
  wire [63:0] acqNet_io_in_1_bits_payload_data;
  wire  acqNet_io_in_2_ready;
  wire  acqNet_io_in_2_valid;
  wire [2:0] acqNet_io_in_2_bits_header_src;
  wire [2:0] acqNet_io_in_2_bits_header_dst;
  wire [25:0] acqNet_io_in_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_2_bits_payload_addr_beat;
  wire  acqNet_io_in_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_2_bits_payload_a_type;
  wire [11:0] acqNet_io_in_2_bits_payload_union;
  wire [63:0] acqNet_io_in_2_bits_payload_data;
  wire  acqNet_io_in_3_ready;
  wire  acqNet_io_in_3_valid;
  wire [2:0] acqNet_io_in_3_bits_header_src;
  wire [2:0] acqNet_io_in_3_bits_header_dst;
  wire [25:0] acqNet_io_in_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_3_bits_payload_addr_beat;
  wire  acqNet_io_in_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_3_bits_payload_a_type;
  wire [11:0] acqNet_io_in_3_bits_payload_union;
  wire [63:0] acqNet_io_in_3_bits_payload_data;
  wire  acqNet_io_in_4_ready;
  wire  acqNet_io_in_4_valid;
  wire [2:0] acqNet_io_in_4_bits_header_src;
  wire [2:0] acqNet_io_in_4_bits_header_dst;
  wire [25:0] acqNet_io_in_4_bits_payload_addr_block;
  wire [1:0] acqNet_io_in_4_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_in_4_bits_payload_addr_beat;
  wire  acqNet_io_in_4_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_in_4_bits_payload_a_type;
  wire [11:0] acqNet_io_in_4_bits_payload_union;
  wire [63:0] acqNet_io_in_4_bits_payload_data;
  wire  acqNet_io_out_0_ready;
  wire  acqNet_io_out_0_valid;
  wire [2:0] acqNet_io_out_0_bits_header_src;
  wire [2:0] acqNet_io_out_0_bits_header_dst;
  wire [25:0] acqNet_io_out_0_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_0_bits_payload_addr_beat;
  wire  acqNet_io_out_0_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_0_bits_payload_a_type;
  wire [11:0] acqNet_io_out_0_bits_payload_union;
  wire [63:0] acqNet_io_out_0_bits_payload_data;
  wire  acqNet_io_out_1_ready;
  wire  acqNet_io_out_1_valid;
  wire [2:0] acqNet_io_out_1_bits_header_src;
  wire [2:0] acqNet_io_out_1_bits_header_dst;
  wire [25:0] acqNet_io_out_1_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_1_bits_payload_addr_beat;
  wire  acqNet_io_out_1_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_1_bits_payload_a_type;
  wire [11:0] acqNet_io_out_1_bits_payload_union;
  wire [63:0] acqNet_io_out_1_bits_payload_data;
  wire  acqNet_io_out_2_ready;
  wire  acqNet_io_out_2_valid;
  wire [2:0] acqNet_io_out_2_bits_header_src;
  wire [2:0] acqNet_io_out_2_bits_header_dst;
  wire [25:0] acqNet_io_out_2_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_2_bits_payload_addr_beat;
  wire  acqNet_io_out_2_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_2_bits_payload_a_type;
  wire [11:0] acqNet_io_out_2_bits_payload_union;
  wire [63:0] acqNet_io_out_2_bits_payload_data;
  wire  acqNet_io_out_3_ready;
  wire  acqNet_io_out_3_valid;
  wire [2:0] acqNet_io_out_3_bits_header_src;
  wire [2:0] acqNet_io_out_3_bits_header_dst;
  wire [25:0] acqNet_io_out_3_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_3_bits_payload_addr_beat;
  wire  acqNet_io_out_3_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_3_bits_payload_a_type;
  wire [11:0] acqNet_io_out_3_bits_payload_union;
  wire [63:0] acqNet_io_out_3_bits_payload_data;
  wire  acqNet_io_out_4_ready;
  wire  acqNet_io_out_4_valid;
  wire [2:0] acqNet_io_out_4_bits_header_src;
  wire [2:0] acqNet_io_out_4_bits_header_dst;
  wire [25:0] acqNet_io_out_4_bits_payload_addr_block;
  wire [1:0] acqNet_io_out_4_bits_payload_client_xact_id;
  wire [2:0] acqNet_io_out_4_bits_payload_addr_beat;
  wire  acqNet_io_out_4_bits_payload_is_builtin_type;
  wire [2:0] acqNet_io_out_4_bits_payload_a_type;
  wire [11:0] acqNet_io_out_4_bits_payload_union;
  wire [63:0] acqNet_io_out_4_bits_payload_data;
  wire  relNet_clk;
  wire  relNet_reset;
  wire  relNet_io_in_0_ready;
  wire  relNet_io_in_0_valid;
  wire [2:0] relNet_io_in_0_bits_header_src;
  wire [2:0] relNet_io_in_0_bits_header_dst;
  wire [2:0] relNet_io_in_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_0_bits_payload_addr_block;
  wire [1:0] relNet_io_in_0_bits_payload_client_xact_id;
  wire  relNet_io_in_0_bits_payload_voluntary;
  wire [2:0] relNet_io_in_0_bits_payload_r_type;
  wire [63:0] relNet_io_in_0_bits_payload_data;
  wire  relNet_io_in_1_ready;
  wire  relNet_io_in_1_valid;
  wire [2:0] relNet_io_in_1_bits_header_src;
  wire [2:0] relNet_io_in_1_bits_header_dst;
  wire [2:0] relNet_io_in_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_1_bits_payload_addr_block;
  wire [1:0] relNet_io_in_1_bits_payload_client_xact_id;
  wire  relNet_io_in_1_bits_payload_voluntary;
  wire [2:0] relNet_io_in_1_bits_payload_r_type;
  wire [63:0] relNet_io_in_1_bits_payload_data;
  wire  relNet_io_in_2_ready;
  wire  relNet_io_in_2_valid;
  wire [2:0] relNet_io_in_2_bits_header_src;
  wire [2:0] relNet_io_in_2_bits_header_dst;
  wire [2:0] relNet_io_in_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_2_bits_payload_addr_block;
  wire [1:0] relNet_io_in_2_bits_payload_client_xact_id;
  wire  relNet_io_in_2_bits_payload_voluntary;
  wire [2:0] relNet_io_in_2_bits_payload_r_type;
  wire [63:0] relNet_io_in_2_bits_payload_data;
  wire  relNet_io_in_3_ready;
  wire  relNet_io_in_3_valid;
  wire [2:0] relNet_io_in_3_bits_header_src;
  wire [2:0] relNet_io_in_3_bits_header_dst;
  wire [2:0] relNet_io_in_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_3_bits_payload_addr_block;
  wire [1:0] relNet_io_in_3_bits_payload_client_xact_id;
  wire  relNet_io_in_3_bits_payload_voluntary;
  wire [2:0] relNet_io_in_3_bits_payload_r_type;
  wire [63:0] relNet_io_in_3_bits_payload_data;
  wire  relNet_io_in_4_ready;
  wire  relNet_io_in_4_valid;
  wire [2:0] relNet_io_in_4_bits_header_src;
  wire [2:0] relNet_io_in_4_bits_header_dst;
  wire [2:0] relNet_io_in_4_bits_payload_addr_beat;
  wire [25:0] relNet_io_in_4_bits_payload_addr_block;
  wire [1:0] relNet_io_in_4_bits_payload_client_xact_id;
  wire  relNet_io_in_4_bits_payload_voluntary;
  wire [2:0] relNet_io_in_4_bits_payload_r_type;
  wire [63:0] relNet_io_in_4_bits_payload_data;
  wire  relNet_io_out_0_ready;
  wire  relNet_io_out_0_valid;
  wire [2:0] relNet_io_out_0_bits_header_src;
  wire [2:0] relNet_io_out_0_bits_header_dst;
  wire [2:0] relNet_io_out_0_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_0_bits_payload_addr_block;
  wire [1:0] relNet_io_out_0_bits_payload_client_xact_id;
  wire  relNet_io_out_0_bits_payload_voluntary;
  wire [2:0] relNet_io_out_0_bits_payload_r_type;
  wire [63:0] relNet_io_out_0_bits_payload_data;
  wire  relNet_io_out_1_ready;
  wire  relNet_io_out_1_valid;
  wire [2:0] relNet_io_out_1_bits_header_src;
  wire [2:0] relNet_io_out_1_bits_header_dst;
  wire [2:0] relNet_io_out_1_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_1_bits_payload_addr_block;
  wire [1:0] relNet_io_out_1_bits_payload_client_xact_id;
  wire  relNet_io_out_1_bits_payload_voluntary;
  wire [2:0] relNet_io_out_1_bits_payload_r_type;
  wire [63:0] relNet_io_out_1_bits_payload_data;
  wire  relNet_io_out_2_ready;
  wire  relNet_io_out_2_valid;
  wire [2:0] relNet_io_out_2_bits_header_src;
  wire [2:0] relNet_io_out_2_bits_header_dst;
  wire [2:0] relNet_io_out_2_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_2_bits_payload_addr_block;
  wire [1:0] relNet_io_out_2_bits_payload_client_xact_id;
  wire  relNet_io_out_2_bits_payload_voluntary;
  wire [2:0] relNet_io_out_2_bits_payload_r_type;
  wire [63:0] relNet_io_out_2_bits_payload_data;
  wire  relNet_io_out_3_ready;
  wire  relNet_io_out_3_valid;
  wire [2:0] relNet_io_out_3_bits_header_src;
  wire [2:0] relNet_io_out_3_bits_header_dst;
  wire [2:0] relNet_io_out_3_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_3_bits_payload_addr_block;
  wire [1:0] relNet_io_out_3_bits_payload_client_xact_id;
  wire  relNet_io_out_3_bits_payload_voluntary;
  wire [2:0] relNet_io_out_3_bits_payload_r_type;
  wire [63:0] relNet_io_out_3_bits_payload_data;
  wire  relNet_io_out_4_ready;
  wire  relNet_io_out_4_valid;
  wire [2:0] relNet_io_out_4_bits_header_src;
  wire [2:0] relNet_io_out_4_bits_header_dst;
  wire [2:0] relNet_io_out_4_bits_payload_addr_beat;
  wire [25:0] relNet_io_out_4_bits_payload_addr_block;
  wire [1:0] relNet_io_out_4_bits_payload_client_xact_id;
  wire  relNet_io_out_4_bits_payload_voluntary;
  wire [2:0] relNet_io_out_4_bits_payload_r_type;
  wire [63:0] relNet_io_out_4_bits_payload_data;
  wire  prbNet_clk;
  wire  prbNet_reset;
  wire  prbNet_io_in_0_ready;
  wire  prbNet_io_in_0_valid;
  wire [2:0] prbNet_io_in_0_bits_header_src;
  wire [2:0] prbNet_io_in_0_bits_header_dst;
  wire [25:0] prbNet_io_in_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_0_bits_payload_p_type;
  wire  prbNet_io_in_1_ready;
  wire  prbNet_io_in_1_valid;
  wire [2:0] prbNet_io_in_1_bits_header_src;
  wire [2:0] prbNet_io_in_1_bits_header_dst;
  wire [25:0] prbNet_io_in_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_1_bits_payload_p_type;
  wire  prbNet_io_in_2_ready;
  wire  prbNet_io_in_2_valid;
  wire [2:0] prbNet_io_in_2_bits_header_src;
  wire [2:0] prbNet_io_in_2_bits_header_dst;
  wire [25:0] prbNet_io_in_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_2_bits_payload_p_type;
  wire  prbNet_io_in_3_ready;
  wire  prbNet_io_in_3_valid;
  wire [2:0] prbNet_io_in_3_bits_header_src;
  wire [2:0] prbNet_io_in_3_bits_header_dst;
  wire [25:0] prbNet_io_in_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_3_bits_payload_p_type;
  wire  prbNet_io_in_4_ready;
  wire  prbNet_io_in_4_valid;
  wire [2:0] prbNet_io_in_4_bits_header_src;
  wire [2:0] prbNet_io_in_4_bits_header_dst;
  wire [25:0] prbNet_io_in_4_bits_payload_addr_block;
  wire [1:0] prbNet_io_in_4_bits_payload_p_type;
  wire  prbNet_io_out_0_ready;
  wire  prbNet_io_out_0_valid;
  wire [2:0] prbNet_io_out_0_bits_header_src;
  wire [2:0] prbNet_io_out_0_bits_header_dst;
  wire [25:0] prbNet_io_out_0_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_0_bits_payload_p_type;
  wire  prbNet_io_out_1_ready;
  wire  prbNet_io_out_1_valid;
  wire [2:0] prbNet_io_out_1_bits_header_src;
  wire [2:0] prbNet_io_out_1_bits_header_dst;
  wire [25:0] prbNet_io_out_1_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_1_bits_payload_p_type;
  wire  prbNet_io_out_2_ready;
  wire  prbNet_io_out_2_valid;
  wire [2:0] prbNet_io_out_2_bits_header_src;
  wire [2:0] prbNet_io_out_2_bits_header_dst;
  wire [25:0] prbNet_io_out_2_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_2_bits_payload_p_type;
  wire  prbNet_io_out_3_ready;
  wire  prbNet_io_out_3_valid;
  wire [2:0] prbNet_io_out_3_bits_header_src;
  wire [2:0] prbNet_io_out_3_bits_header_dst;
  wire [25:0] prbNet_io_out_3_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_3_bits_payload_p_type;
  wire  prbNet_io_out_4_ready;
  wire  prbNet_io_out_4_valid;
  wire [2:0] prbNet_io_out_4_bits_header_src;
  wire [2:0] prbNet_io_out_4_bits_header_dst;
  wire [25:0] prbNet_io_out_4_bits_payload_addr_block;
  wire [1:0] prbNet_io_out_4_bits_payload_p_type;
  wire  gntNet_clk;
  wire  gntNet_reset;
  wire  gntNet_io_in_0_ready;
  wire  gntNet_io_in_0_valid;
  wire [2:0] gntNet_io_in_0_bits_header_src;
  wire [2:0] gntNet_io_in_0_bits_header_dst;
  wire [2:0] gntNet_io_in_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_0_bits_payload_manager_xact_id;
  wire  gntNet_io_in_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_0_bits_payload_g_type;
  wire [63:0] gntNet_io_in_0_bits_payload_data;
  wire  gntNet_io_in_1_ready;
  wire  gntNet_io_in_1_valid;
  wire [2:0] gntNet_io_in_1_bits_header_src;
  wire [2:0] gntNet_io_in_1_bits_header_dst;
  wire [2:0] gntNet_io_in_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_1_bits_payload_manager_xact_id;
  wire  gntNet_io_in_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_1_bits_payload_g_type;
  wire [63:0] gntNet_io_in_1_bits_payload_data;
  wire  gntNet_io_in_2_ready;
  wire  gntNet_io_in_2_valid;
  wire [2:0] gntNet_io_in_2_bits_header_src;
  wire [2:0] gntNet_io_in_2_bits_header_dst;
  wire [2:0] gntNet_io_in_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_2_bits_payload_manager_xact_id;
  wire  gntNet_io_in_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_2_bits_payload_g_type;
  wire [63:0] gntNet_io_in_2_bits_payload_data;
  wire  gntNet_io_in_3_ready;
  wire  gntNet_io_in_3_valid;
  wire [2:0] gntNet_io_in_3_bits_header_src;
  wire [2:0] gntNet_io_in_3_bits_header_dst;
  wire [2:0] gntNet_io_in_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_3_bits_payload_manager_xact_id;
  wire  gntNet_io_in_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_3_bits_payload_g_type;
  wire [63:0] gntNet_io_in_3_bits_payload_data;
  wire  gntNet_io_in_4_ready;
  wire  gntNet_io_in_4_valid;
  wire [2:0] gntNet_io_in_4_bits_header_src;
  wire [2:0] gntNet_io_in_4_bits_header_dst;
  wire [2:0] gntNet_io_in_4_bits_payload_addr_beat;
  wire [1:0] gntNet_io_in_4_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_in_4_bits_payload_manager_xact_id;
  wire  gntNet_io_in_4_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_in_4_bits_payload_g_type;
  wire [63:0] gntNet_io_in_4_bits_payload_data;
  wire  gntNet_io_out_0_ready;
  wire  gntNet_io_out_0_valid;
  wire [2:0] gntNet_io_out_0_bits_header_src;
  wire [2:0] gntNet_io_out_0_bits_header_dst;
  wire [2:0] gntNet_io_out_0_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_0_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_0_bits_payload_manager_xact_id;
  wire  gntNet_io_out_0_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_0_bits_payload_g_type;
  wire [63:0] gntNet_io_out_0_bits_payload_data;
  wire  gntNet_io_out_1_ready;
  wire  gntNet_io_out_1_valid;
  wire [2:0] gntNet_io_out_1_bits_header_src;
  wire [2:0] gntNet_io_out_1_bits_header_dst;
  wire [2:0] gntNet_io_out_1_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_1_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_1_bits_payload_manager_xact_id;
  wire  gntNet_io_out_1_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_1_bits_payload_g_type;
  wire [63:0] gntNet_io_out_1_bits_payload_data;
  wire  gntNet_io_out_2_ready;
  wire  gntNet_io_out_2_valid;
  wire [2:0] gntNet_io_out_2_bits_header_src;
  wire [2:0] gntNet_io_out_2_bits_header_dst;
  wire [2:0] gntNet_io_out_2_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_2_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_2_bits_payload_manager_xact_id;
  wire  gntNet_io_out_2_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_2_bits_payload_g_type;
  wire [63:0] gntNet_io_out_2_bits_payload_data;
  wire  gntNet_io_out_3_ready;
  wire  gntNet_io_out_3_valid;
  wire [2:0] gntNet_io_out_3_bits_header_src;
  wire [2:0] gntNet_io_out_3_bits_header_dst;
  wire [2:0] gntNet_io_out_3_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_3_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_3_bits_payload_manager_xact_id;
  wire  gntNet_io_out_3_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_3_bits_payload_g_type;
  wire [63:0] gntNet_io_out_3_bits_payload_data;
  wire  gntNet_io_out_4_ready;
  wire  gntNet_io_out_4_valid;
  wire [2:0] gntNet_io_out_4_bits_header_src;
  wire [2:0] gntNet_io_out_4_bits_header_dst;
  wire [2:0] gntNet_io_out_4_bits_payload_addr_beat;
  wire [1:0] gntNet_io_out_4_bits_payload_client_xact_id;
  wire [2:0] gntNet_io_out_4_bits_payload_manager_xact_id;
  wire  gntNet_io_out_4_bits_payload_is_builtin_type;
  wire [3:0] gntNet_io_out_4_bits_payload_g_type;
  wire [63:0] gntNet_io_out_4_bits_payload_data;
  wire  ackNet_clk;
  wire  ackNet_reset;
  wire  ackNet_io_in_0_ready;
  wire  ackNet_io_in_0_valid;
  wire [2:0] ackNet_io_in_0_bits_header_src;
  wire [2:0] ackNet_io_in_0_bits_header_dst;
  wire [2:0] ackNet_io_in_0_bits_payload_manager_xact_id;
  wire  ackNet_io_in_1_ready;
  wire  ackNet_io_in_1_valid;
  wire [2:0] ackNet_io_in_1_bits_header_src;
  wire [2:0] ackNet_io_in_1_bits_header_dst;
  wire [2:0] ackNet_io_in_1_bits_payload_manager_xact_id;
  wire  ackNet_io_in_2_ready;
  wire  ackNet_io_in_2_valid;
  wire [2:0] ackNet_io_in_2_bits_header_src;
  wire [2:0] ackNet_io_in_2_bits_header_dst;
  wire [2:0] ackNet_io_in_2_bits_payload_manager_xact_id;
  wire  ackNet_io_in_3_ready;
  wire  ackNet_io_in_3_valid;
  wire [2:0] ackNet_io_in_3_bits_header_src;
  wire [2:0] ackNet_io_in_3_bits_header_dst;
  wire [2:0] ackNet_io_in_3_bits_payload_manager_xact_id;
  wire  ackNet_io_in_4_ready;
  wire  ackNet_io_in_4_valid;
  wire [2:0] ackNet_io_in_4_bits_header_src;
  wire [2:0] ackNet_io_in_4_bits_header_dst;
  wire [2:0] ackNet_io_in_4_bits_payload_manager_xact_id;
  wire  ackNet_io_out_0_ready;
  wire  ackNet_io_out_0_valid;
  wire [2:0] ackNet_io_out_0_bits_header_src;
  wire [2:0] ackNet_io_out_0_bits_header_dst;
  wire [2:0] ackNet_io_out_0_bits_payload_manager_xact_id;
  wire  ackNet_io_out_1_ready;
  wire  ackNet_io_out_1_valid;
  wire [2:0] ackNet_io_out_1_bits_header_src;
  wire [2:0] ackNet_io_out_1_bits_header_dst;
  wire [2:0] ackNet_io_out_1_bits_payload_manager_xact_id;
  wire  ackNet_io_out_2_ready;
  wire  ackNet_io_out_2_valid;
  wire [2:0] ackNet_io_out_2_bits_header_src;
  wire [2:0] ackNet_io_out_2_bits_header_dst;
  wire [2:0] ackNet_io_out_2_bits_payload_manager_xact_id;
  wire  ackNet_io_out_3_ready;
  wire  ackNet_io_out_3_valid;
  wire [2:0] ackNet_io_out_3_bits_header_src;
  wire [2:0] ackNet_io_out_3_bits_header_dst;
  wire [2:0] ackNet_io_out_3_bits_payload_manager_xact_id;
  wire  ackNet_io_out_4_ready;
  wire  ackNet_io_out_4_valid;
  wire [2:0] ackNet_io_out_4_bits_header_src;
  wire [2:0] ackNet_io_out_4_bits_header_dst;
  wire [2:0] ackNet_io_out_4_bits_payload_manager_xact_id;
  wire  T_14709_ready;
  wire  T_14709_valid;
  wire [2:0] T_14709_bits_header_src;
  wire [2:0] T_14709_bits_header_dst;
  wire [25:0] T_14709_bits_payload_addr_block;
  wire [1:0] T_14709_bits_payload_client_xact_id;
  wire [2:0] T_14709_bits_payload_addr_beat;
  wire  T_14709_bits_payload_is_builtin_type;
  wire [2:0] T_14709_bits_payload_a_type;
  wire [11:0] T_14709_bits_payload_union;
  wire [63:0] T_14709_bits_payload_data;
  wire [2:0] GEN_0;
  wire [3:0] T_14967;
  wire [2:0] T_14968;
  wire  T_15354_ready;
  wire  T_15354_valid;
  wire [2:0] T_15354_bits_header_src;
  wire [2:0] T_15354_bits_header_dst;
  wire [25:0] T_15354_bits_payload_addr_block;
  wire [1:0] T_15354_bits_payload_client_xact_id;
  wire [2:0] T_15354_bits_payload_addr_beat;
  wire  T_15354_bits_payload_is_builtin_type;
  wire [2:0] T_15354_bits_payload_a_type;
  wire [11:0] T_15354_bits_payload_union;
  wire [63:0] T_15354_bits_payload_data;
  wire [3:0] T_15612;
  wire [2:0] T_15613;
  wire  T_15723_ready;
  wire  T_15723_valid;
  wire [2:0] T_15723_bits_header_src;
  wire [2:0] T_15723_bits_header_dst;
  wire [25:0] T_15723_bits_payload_addr_block;
  wire [1:0] T_15723_bits_payload_client_xact_id;
  wire [2:0] T_15723_bits_payload_addr_beat;
  wire  T_15723_bits_payload_is_builtin_type;
  wire [2:0] T_15723_bits_payload_a_type;
  wire [11:0] T_15723_bits_payload_union;
  wire [63:0] T_15723_bits_payload_data;
  wire [3:0] T_15797;
  wire [2:0] T_15798;
  wire  T_15908_ready;
  wire  T_15908_valid;
  wire [2:0] T_15908_bits_header_src;
  wire [2:0] T_15908_bits_header_dst;
  wire [25:0] T_15908_bits_payload_addr_block;
  wire [1:0] T_15908_bits_payload_client_xact_id;
  wire [2:0] T_15908_bits_payload_addr_beat;
  wire  T_15908_bits_payload_is_builtin_type;
  wire [2:0] T_15908_bits_payload_a_type;
  wire [11:0] T_15908_bits_payload_union;
  wire [63:0] T_15908_bits_payload_data;
  wire [3:0] T_15982;
  wire [2:0] T_15983;
  wire  T_16093_ready;
  wire  T_16093_valid;
  wire [2:0] T_16093_bits_header_src;
  wire [2:0] T_16093_bits_header_dst;
  wire [25:0] T_16093_bits_payload_addr_block;
  wire [1:0] T_16093_bits_payload_client_xact_id;
  wire [2:0] T_16093_bits_payload_addr_beat;
  wire  T_16093_bits_payload_is_builtin_type;
  wire [2:0] T_16093_bits_payload_a_type;
  wire [11:0] T_16093_bits_payload_union;
  wire [63:0] T_16093_bits_payload_data;
  wire [3:0] T_16167;
  wire [2:0] T_16168;
  wire  T_16551_ready;
  wire  T_16551_valid;
  wire [2:0] T_16551_bits_header_src;
  wire [2:0] T_16551_bits_header_dst;
  wire [2:0] T_16551_bits_payload_addr_beat;
  wire [25:0] T_16551_bits_payload_addr_block;
  wire [1:0] T_16551_bits_payload_client_xact_id;
  wire  T_16551_bits_payload_voluntary;
  wire [2:0] T_16551_bits_payload_r_type;
  wire [63:0] T_16551_bits_payload_data;
  wire [3:0] T_16807;
  wire [2:0] T_16808;
  wire  T_17191_ready;
  wire  T_17191_valid;
  wire [2:0] T_17191_bits_header_src;
  wire [2:0] T_17191_bits_header_dst;
  wire [2:0] T_17191_bits_payload_addr_beat;
  wire [25:0] T_17191_bits_payload_addr_block;
  wire [1:0] T_17191_bits_payload_client_xact_id;
  wire  T_17191_bits_payload_voluntary;
  wire [2:0] T_17191_bits_payload_r_type;
  wire [63:0] T_17191_bits_payload_data;
  wire [3:0] T_17447;
  wire [2:0] T_17448;
  wire  T_17555_ready;
  wire  T_17555_valid;
  wire [2:0] T_17555_bits_header_src;
  wire [2:0] T_17555_bits_header_dst;
  wire [2:0] T_17555_bits_payload_addr_beat;
  wire [25:0] T_17555_bits_payload_addr_block;
  wire [1:0] T_17555_bits_payload_client_xact_id;
  wire  T_17555_bits_payload_voluntary;
  wire [2:0] T_17555_bits_payload_r_type;
  wire [63:0] T_17555_bits_payload_data;
  wire [3:0] T_17627;
  wire [2:0] T_17628;
  wire  T_17735_ready;
  wire  T_17735_valid;
  wire [2:0] T_17735_bits_header_src;
  wire [2:0] T_17735_bits_header_dst;
  wire [2:0] T_17735_bits_payload_addr_beat;
  wire [25:0] T_17735_bits_payload_addr_block;
  wire [1:0] T_17735_bits_payload_client_xact_id;
  wire  T_17735_bits_payload_voluntary;
  wire [2:0] T_17735_bits_payload_r_type;
  wire [63:0] T_17735_bits_payload_data;
  wire [3:0] T_17807;
  wire [2:0] T_17808;
  wire  T_17915_ready;
  wire  T_17915_valid;
  wire [2:0] T_17915_bits_header_src;
  wire [2:0] T_17915_bits_header_dst;
  wire [2:0] T_17915_bits_payload_addr_beat;
  wire [25:0] T_17915_bits_payload_addr_block;
  wire [1:0] T_17915_bits_payload_client_xact_id;
  wire  T_17915_bits_payload_voluntary;
  wire [2:0] T_17915_bits_payload_r_type;
  wire [63:0] T_17915_bits_payload_data;
  wire [3:0] T_17987;
  wire [2:0] T_17988;
  wire  T_18083_ready;
  wire  T_18083_valid;
  wire [2:0] T_18083_bits_header_src;
  wire [2:0] T_18083_bits_header_dst;
  wire [25:0] T_18083_bits_payload_addr_block;
  wire [1:0] T_18083_bits_payload_p_type;
  wire [3:0] T_18147;
  wire [2:0] T_18148;
  wire  T_18243_ready;
  wire  T_18243_valid;
  wire [2:0] T_18243_bits_header_src;
  wire [2:0] T_18243_bits_header_dst;
  wire [25:0] T_18243_bits_payload_addr_block;
  wire [1:0] T_18243_bits_payload_p_type;
  wire [3:0] T_18307;
  wire [2:0] T_18308;
  wire  T_18679_ready;
  wire  T_18679_valid;
  wire [2:0] T_18679_bits_header_src;
  wire [2:0] T_18679_bits_header_dst;
  wire [25:0] T_18679_bits_payload_addr_block;
  wire [1:0] T_18679_bits_payload_p_type;
  wire [3:0] T_18927;
  wire [2:0] T_18928;
  wire  T_19299_ready;
  wire  T_19299_valid;
  wire [2:0] T_19299_bits_header_src;
  wire [2:0] T_19299_bits_header_dst;
  wire [25:0] T_19299_bits_payload_addr_block;
  wire [1:0] T_19299_bits_payload_p_type;
  wire [3:0] T_19547;
  wire [2:0] T_19548;
  wire  T_19919_ready;
  wire  T_19919_valid;
  wire [2:0] T_19919_bits_header_src;
  wire [2:0] T_19919_bits_header_dst;
  wire [25:0] T_19919_bits_payload_addr_block;
  wire [1:0] T_19919_bits_payload_p_type;
  wire [3:0] T_20167;
  wire [2:0] T_20168;
  wire  T_20275_ready;
  wire  T_20275_valid;
  wire [2:0] T_20275_bits_header_src;
  wire [2:0] T_20275_bits_header_dst;
  wire [2:0] T_20275_bits_payload_addr_beat;
  wire [1:0] T_20275_bits_payload_client_xact_id;
  wire [2:0] T_20275_bits_payload_manager_xact_id;
  wire  T_20275_bits_payload_is_builtin_type;
  wire [3:0] T_20275_bits_payload_g_type;
  wire [63:0] T_20275_bits_payload_data;
  wire [3:0] T_20347;
  wire [2:0] T_20348;
  wire  T_20455_ready;
  wire  T_20455_valid;
  wire [2:0] T_20455_bits_header_src;
  wire [2:0] T_20455_bits_header_dst;
  wire [2:0] T_20455_bits_payload_addr_beat;
  wire [1:0] T_20455_bits_payload_client_xact_id;
  wire [2:0] T_20455_bits_payload_manager_xact_id;
  wire  T_20455_bits_payload_is_builtin_type;
  wire [3:0] T_20455_bits_payload_g_type;
  wire [63:0] T_20455_bits_payload_data;
  wire [3:0] T_20527;
  wire [2:0] T_20528;
  wire  T_20911_ready;
  wire  T_20911_valid;
  wire [2:0] T_20911_bits_header_src;
  wire [2:0] T_20911_bits_header_dst;
  wire [2:0] T_20911_bits_payload_addr_beat;
  wire [1:0] T_20911_bits_payload_client_xact_id;
  wire [2:0] T_20911_bits_payload_manager_xact_id;
  wire  T_20911_bits_payload_is_builtin_type;
  wire [3:0] T_20911_bits_payload_g_type;
  wire [63:0] T_20911_bits_payload_data;
  wire [3:0] T_21167;
  wire [2:0] T_21168;
  wire  T_21551_ready;
  wire  T_21551_valid;
  wire [2:0] T_21551_bits_header_src;
  wire [2:0] T_21551_bits_header_dst;
  wire [2:0] T_21551_bits_payload_addr_beat;
  wire [1:0] T_21551_bits_payload_client_xact_id;
  wire [2:0] T_21551_bits_payload_manager_xact_id;
  wire  T_21551_bits_payload_is_builtin_type;
  wire [3:0] T_21551_bits_payload_g_type;
  wire [63:0] T_21551_bits_payload_data;
  wire [3:0] T_21807;
  wire [2:0] T_21808;
  wire  T_22191_ready;
  wire  T_22191_valid;
  wire [2:0] T_22191_bits_header_src;
  wire [2:0] T_22191_bits_header_dst;
  wire [2:0] T_22191_bits_payload_addr_beat;
  wire [1:0] T_22191_bits_payload_client_xact_id;
  wire [2:0] T_22191_bits_payload_manager_xact_id;
  wire  T_22191_bits_payload_is_builtin_type;
  wire [3:0] T_22191_bits_payload_g_type;
  wire [63:0] T_22191_bits_payload_data;
  wire [3:0] T_22447;
  wire [2:0] T_22448;
  wire  T_22816_ready;
  wire  T_22816_valid;
  wire [2:0] T_22816_bits_header_src;
  wire [2:0] T_22816_bits_header_dst;
  wire [2:0] T_22816_bits_payload_manager_xact_id;
  wire [3:0] T_23062;
  wire [2:0] T_23063;
  wire  T_23431_ready;
  wire  T_23431_valid;
  wire [2:0] T_23431_bits_header_src;
  wire [2:0] T_23431_bits_header_dst;
  wire [2:0] T_23431_bits_payload_manager_xact_id;
  wire [3:0] T_23677;
  wire [2:0] T_23678;
  wire  T_23770_ready;
  wire  T_23770_valid;
  wire [2:0] T_23770_bits_header_src;
  wire [2:0] T_23770_bits_header_dst;
  wire [2:0] T_23770_bits_payload_manager_xact_id;
  wire [3:0] T_23832;
  wire [2:0] T_23833;
  wire  T_23925_ready;
  wire  T_23925_valid;
  wire [2:0] T_23925_bits_header_src;
  wire [2:0] T_23925_bits_header_dst;
  wire [2:0] T_23925_bits_payload_manager_xact_id;
  wire [3:0] T_23987;
  wire [2:0] T_23988;
  wire  T_24080_ready;
  wire  T_24080_valid;
  wire [2:0] T_24080_bits_header_src;
  wire [2:0] T_24080_bits_header_dst;
  wire [2:0] T_24080_bits_payload_manager_xact_id;
  wire [3:0] T_24142;
  wire [2:0] T_24143;
  reg [2:0] GEN_1;
  reg [31:0] GEN_77;
  reg [2:0] GEN_2;
  reg [31:0] GEN_78;
  reg [25:0] GEN_3;
  reg [31:0] GEN_79;
  reg [1:0] GEN_4;
  reg [31:0] GEN_80;
  reg [2:0] GEN_5;
  reg [31:0] GEN_81;
  reg  GEN_6;
  reg [31:0] GEN_82;
  reg [2:0] GEN_7;
  reg [31:0] GEN_83;
  reg [11:0] GEN_8;
  reg [31:0] GEN_84;
  reg [63:0] GEN_9;
  reg [63:0] GEN_85;
  reg [2:0] GEN_10;
  reg [31:0] GEN_86;
  reg [2:0] GEN_11;
  reg [31:0] GEN_87;
  reg [25:0] GEN_12;
  reg [31:0] GEN_88;
  reg [1:0] GEN_13;
  reg [31:0] GEN_89;
  reg [2:0] GEN_14;
  reg [31:0] GEN_90;
  reg  GEN_15;
  reg [31:0] GEN_91;
  reg [2:0] GEN_16;
  reg [31:0] GEN_92;
  reg [11:0] GEN_17;
  reg [31:0] GEN_93;
  reg [63:0] GEN_18;
  reg [63:0] GEN_94;
  reg [2:0] GEN_19;
  reg [31:0] GEN_95;
  reg [2:0] GEN_20;
  reg [31:0] GEN_96;
  reg [2:0] GEN_21;
  reg [31:0] GEN_97;
  reg [25:0] GEN_22;
  reg [31:0] GEN_98;
  reg [1:0] GEN_23;
  reg [31:0] GEN_99;
  reg  GEN_24;
  reg [31:0] GEN_100;
  reg [2:0] GEN_25;
  reg [31:0] GEN_101;
  reg [63:0] GEN_26;
  reg [63:0] GEN_102;
  reg [2:0] GEN_27;
  reg [31:0] GEN_103;
  reg [2:0] GEN_28;
  reg [31:0] GEN_104;
  reg [2:0] GEN_29;
  reg [31:0] GEN_105;
  reg [25:0] GEN_30;
  reg [31:0] GEN_106;
  reg [1:0] GEN_31;
  reg [31:0] GEN_107;
  reg  GEN_32;
  reg [31:0] GEN_108;
  reg [2:0] GEN_33;
  reg [31:0] GEN_109;
  reg [63:0] GEN_34;
  reg [63:0] GEN_110;
  reg [2:0] GEN_35;
  reg [31:0] GEN_111;
  reg [2:0] GEN_36;
  reg [31:0] GEN_112;
  reg [25:0] GEN_37;
  reg [31:0] GEN_113;
  reg [1:0] GEN_38;
  reg [31:0] GEN_114;
  reg [2:0] GEN_39;
  reg [31:0] GEN_115;
  reg [2:0] GEN_40;
  reg [31:0] GEN_116;
  reg [25:0] GEN_41;
  reg [31:0] GEN_117;
  reg [1:0] GEN_42;
  reg [31:0] GEN_118;
  reg [2:0] GEN_43;
  reg [31:0] GEN_119;
  reg [2:0] GEN_44;
  reg [31:0] GEN_120;
  reg [25:0] GEN_45;
  reg [31:0] GEN_121;
  reg [1:0] GEN_46;
  reg [31:0] GEN_122;
  reg [2:0] GEN_47;
  reg [31:0] GEN_123;
  reg [2:0] GEN_48;
  reg [31:0] GEN_124;
  reg [2:0] GEN_49;
  reg [31:0] GEN_125;
  reg [1:0] GEN_50;
  reg [31:0] GEN_126;
  reg [2:0] GEN_51;
  reg [31:0] GEN_127;
  reg  GEN_52;
  reg [31:0] GEN_128;
  reg [3:0] GEN_53;
  reg [31:0] GEN_129;
  reg [63:0] GEN_54;
  reg [63:0] GEN_130;
  reg [2:0] GEN_55;
  reg [31:0] GEN_131;
  reg [2:0] GEN_56;
  reg [31:0] GEN_132;
  reg [2:0] GEN_57;
  reg [31:0] GEN_133;
  reg [1:0] GEN_58;
  reg [31:0] GEN_134;
  reg [2:0] GEN_59;
  reg [31:0] GEN_135;
  reg  GEN_60;
  reg [31:0] GEN_136;
  reg [3:0] GEN_61;
  reg [31:0] GEN_137;
  reg [63:0] GEN_62;
  reg [63:0] GEN_138;
  reg [2:0] GEN_63;
  reg [31:0] GEN_139;
  reg [2:0] GEN_64;
  reg [31:0] GEN_140;
  reg [2:0] GEN_65;
  reg [31:0] GEN_141;
  reg [1:0] GEN_66;
  reg [31:0] GEN_142;
  reg [2:0] GEN_67;
  reg [31:0] GEN_143;
  reg  GEN_68;
  reg [31:0] GEN_144;
  reg [3:0] GEN_69;
  reg [31:0] GEN_145;
  reg [63:0] GEN_70;
  reg [63:0] GEN_146;
  reg [2:0] GEN_71;
  reg [31:0] GEN_147;
  reg [2:0] GEN_72;
  reg [31:0] GEN_148;
  reg [2:0] GEN_73;
  reg [31:0] GEN_149;
  reg [2:0] GEN_74;
  reg [31:0] GEN_150;
  reg [2:0] GEN_75;
  reg [31:0] GEN_151;
  reg [2:0] GEN_76;
  reg [31:0] GEN_152;
  TileLinkEnqueuer TileLinkEnqueuer_14127 (
    .clk(TileLinkEnqueuer_14127_clk),
    .reset(TileLinkEnqueuer_14127_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_14127_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_14127_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_14127_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_14127_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_14127_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_14127_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_14127_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_14127_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_14127_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_14127_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_14127_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_14127_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_14127_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_14127_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_14127_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_14127_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_14127_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_14127_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_14127_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_14127_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_14127_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_14127_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_14127_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_14127_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_14127_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_14127_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_14127_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_14127_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_14127_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_14127_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_14127_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_14127_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_14127_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_14127_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_14127_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_14127_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_14127_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_14127_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_14127_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_14127_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_14127_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_14127_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_14127_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_14127_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_14127_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_14127_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_14127_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_14127_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_14127_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_14127_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_14127_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_14127_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_14127_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_14127_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_14127_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_14127_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_14127_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_14127_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_14127_io_manager_release_bits_payload_data)
  );
  ClientTileLinkNetworkPort ClientTileLinkNetworkPort_14128 (
    .clk(ClientTileLinkNetworkPort_14128_clk),
    .reset(ClientTileLinkNetworkPort_14128_reset),
    .io_client_acquire_ready(ClientTileLinkNetworkPort_14128_io_client_acquire_ready),
    .io_client_acquire_valid(ClientTileLinkNetworkPort_14128_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientTileLinkNetworkPort_14128_io_client_acquire_bits_data),
    .io_client_probe_ready(ClientTileLinkNetworkPort_14128_io_client_probe_ready),
    .io_client_probe_valid(ClientTileLinkNetworkPort_14128_io_client_probe_valid),
    .io_client_probe_bits_addr_block(ClientTileLinkNetworkPort_14128_io_client_probe_bits_addr_block),
    .io_client_probe_bits_p_type(ClientTileLinkNetworkPort_14128_io_client_probe_bits_p_type),
    .io_client_release_ready(ClientTileLinkNetworkPort_14128_io_client_release_ready),
    .io_client_release_valid(ClientTileLinkNetworkPort_14128_io_client_release_valid),
    .io_client_release_bits_addr_beat(ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_beat),
    .io_client_release_bits_addr_block(ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_block),
    .io_client_release_bits_client_xact_id(ClientTileLinkNetworkPort_14128_io_client_release_bits_client_xact_id),
    .io_client_release_bits_voluntary(ClientTileLinkNetworkPort_14128_io_client_release_bits_voluntary),
    .io_client_release_bits_r_type(ClientTileLinkNetworkPort_14128_io_client_release_bits_r_type),
    .io_client_release_bits_data(ClientTileLinkNetworkPort_14128_io_client_release_bits_data),
    .io_client_grant_ready(ClientTileLinkNetworkPort_14128_io_client_grant_ready),
    .io_client_grant_valid(ClientTileLinkNetworkPort_14128_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientTileLinkNetworkPort_14128_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientTileLinkNetworkPort_14128_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientTileLinkNetworkPort_14128_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientTileLinkNetworkPort_14128_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientTileLinkNetworkPort_14128_io_client_grant_bits_data),
    .io_client_grant_bits_manager_id(ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_id),
    .io_client_finish_ready(ClientTileLinkNetworkPort_14128_io_client_finish_ready),
    .io_client_finish_valid(ClientTileLinkNetworkPort_14128_io_client_finish_valid),
    .io_client_finish_bits_manager_xact_id(ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_xact_id),
    .io_client_finish_bits_manager_id(ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_id),
    .io_network_acquire_ready(ClientTileLinkNetworkPort_14128_io_network_acquire_ready),
    .io_network_acquire_valid(ClientTileLinkNetworkPort_14128_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientTileLinkNetworkPort_14128_io_network_grant_ready),
    .io_network_grant_valid(ClientTileLinkNetworkPort_14128_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientTileLinkNetworkPort_14128_io_network_finish_ready),
    .io_network_finish_valid(ClientTileLinkNetworkPort_14128_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientTileLinkNetworkPort_14128_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientTileLinkNetworkPort_14128_io_network_probe_ready),
    .io_network_probe_valid(ClientTileLinkNetworkPort_14128_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientTileLinkNetworkPort_14128_io_network_release_ready),
    .io_network_release_valid(ClientTileLinkNetworkPort_14128_io_network_release_valid),
    .io_network_release_bits_header_src(ClientTileLinkNetworkPort_14128_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientTileLinkNetworkPort_14128_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_4 TileLinkEnqueuer_4_14129 (
    .clk(TileLinkEnqueuer_4_14129_clk),
    .reset(TileLinkEnqueuer_4_14129_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_4_14129_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_4_14129_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_4_14129_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_4_14129_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_4_14129_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_4_14129_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_4_14129_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_4_14129_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_4_14129_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_4_14129_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_14129_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_4_14129_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_4_14129_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_4_14129_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_4_14129_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_4_14129_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_4_14129_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_4_14129_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_4_14129_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_4_14129_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_4_14129_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_4_14129_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_4_14129_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_4_14129_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_4_14129_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_4_14129_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_4_14129_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_4_14129_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_4_14129_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_4_14129_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_4_14129_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_4_14129_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_4_14129_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort ClientUncachedTileLinkNetworkPort_14130 (
    .clk(ClientUncachedTileLinkNetworkPort_14130_clk),
    .reset(ClientUncachedTileLinkNetworkPort_14130_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_14130_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_14130_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_14130_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_14130_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_9 TileLinkEnqueuer_9_14131 (
    .clk(TileLinkEnqueuer_9_14131_clk),
    .reset(TileLinkEnqueuer_9_14131_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_9_14131_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_9_14131_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_9_14131_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_9_14131_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_9_14131_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_9_14131_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_9_14131_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_9_14131_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_9_14131_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_9_14131_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_9_14131_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_9_14131_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_9_14131_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_9_14131_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_9_14131_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_9_14131_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_9_14131_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_9_14131_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_9_14131_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_9_14131_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_9_14131_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_9_14131_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_9_14131_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_9_14131_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_9_14131_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_9_14131_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_9_14131_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_9_14131_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_9_14131_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_9_14131_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_9_14131_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_9_14131_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_9_14131_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_data)
  );
  ClientUncachedTileLinkNetworkPort_14 ClientUncachedTileLinkNetworkPort_14_14132 (
    .clk(ClientUncachedTileLinkNetworkPort_14_14132_clk),
    .reset(ClientUncachedTileLinkNetworkPort_14_14132_reset),
    .io_client_acquire_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_ready),
    .io_client_acquire_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_valid),
    .io_client_acquire_bits_addr_block(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_block),
    .io_client_acquire_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_client_xact_id),
    .io_client_acquire_bits_addr_beat(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_beat),
    .io_client_acquire_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_is_builtin_type),
    .io_client_acquire_bits_a_type(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_a_type),
    .io_client_acquire_bits_union(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_union),
    .io_client_acquire_bits_data(ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_data),
    .io_client_grant_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_ready),
    .io_client_grant_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_valid),
    .io_client_grant_bits_addr_beat(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_addr_beat),
    .io_client_grant_bits_client_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_client_xact_id),
    .io_client_grant_bits_manager_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_manager_xact_id),
    .io_client_grant_bits_is_builtin_type(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_is_builtin_type),
    .io_client_grant_bits_g_type(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_g_type),
    .io_client_grant_bits_data(ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_data),
    .io_network_acquire_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_ready),
    .io_network_acquire_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_ready),
    .io_network_grant_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_valid),
    .io_network_grant_bits_header_src(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_ready),
    .io_network_finish_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_valid),
    .io_network_finish_bits_header_src(ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_ready),
    .io_network_probe_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_valid),
    .io_network_probe_bits_header_src(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_ready),
    .io_network_release_valid(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_valid),
    .io_network_release_bits_header_src(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort ManagerTileLinkNetworkPort_14133 (
    .clk(ManagerTileLinkNetworkPort_14133_clk),
    .reset(ManagerTileLinkNetworkPort_14133_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_14133_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_14133_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_14133_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_14133_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_14133_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_14133_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_14133_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_14133_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_14133_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_14133_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_14133_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_14133_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_14133_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_14133_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_14133_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_14133_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_14133_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_14133_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_14133_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_14133_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_14133_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_14133_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_17 TileLinkEnqueuer_17_14134 (
    .clk(TileLinkEnqueuer_17_14134_clk),
    .reset(TileLinkEnqueuer_17_14134_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_17_14134_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_17_14134_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_17_14134_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_17_14134_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_17_14134_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_17_14134_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_17_14134_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_17_14134_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_17_14134_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_17_14134_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_17_14134_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_17_14134_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_17_14134_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_17_14134_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_17_14134_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_17_14134_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_17_14134_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_17_14134_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_17_14134_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_17_14134_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_17_14134_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_17_14134_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_17_14134_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_17_14134_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_17_14134_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_17_14134_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_17_14134_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_17_14134_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_17_14134_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_17_14134_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_17_14134_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_17_14134_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_17_14134_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_data)
  );
  ManagerTileLinkNetworkPort_18 ManagerTileLinkNetworkPort_18_14135 (
    .clk(ManagerTileLinkNetworkPort_18_14135_clk),
    .reset(ManagerTileLinkNetworkPort_18_14135_reset),
    .io_manager_acquire_ready(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_ready),
    .io_manager_acquire_valid(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_valid),
    .io_manager_acquire_bits_addr_block(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_block),
    .io_manager_acquire_bits_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_xact_id),
    .io_manager_acquire_bits_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_beat),
    .io_manager_acquire_bits_is_builtin_type(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_is_builtin_type),
    .io_manager_acquire_bits_a_type(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_a_type),
    .io_manager_acquire_bits_union(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_union),
    .io_manager_acquire_bits_data(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_data),
    .io_manager_acquire_bits_client_id(ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_id),
    .io_manager_grant_ready(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_ready),
    .io_manager_grant_valid(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_valid),
    .io_manager_grant_bits_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_addr_beat),
    .io_manager_grant_bits_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_xact_id),
    .io_manager_grant_bits_manager_xact_id(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_manager_xact_id),
    .io_manager_grant_bits_is_builtin_type(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_is_builtin_type),
    .io_manager_grant_bits_g_type(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_g_type),
    .io_manager_grant_bits_data(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_data),
    .io_manager_grant_bits_client_id(ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_id),
    .io_manager_finish_ready(ManagerTileLinkNetworkPort_18_14135_io_manager_finish_ready),
    .io_manager_finish_valid(ManagerTileLinkNetworkPort_18_14135_io_manager_finish_valid),
    .io_manager_finish_bits_manager_xact_id(ManagerTileLinkNetworkPort_18_14135_io_manager_finish_bits_manager_xact_id),
    .io_manager_probe_ready(ManagerTileLinkNetworkPort_18_14135_io_manager_probe_ready),
    .io_manager_probe_valid(ManagerTileLinkNetworkPort_18_14135_io_manager_probe_valid),
    .io_manager_probe_bits_addr_block(ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_addr_block),
    .io_manager_probe_bits_p_type(ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_p_type),
    .io_manager_probe_bits_client_id(ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_client_id),
    .io_manager_release_ready(ManagerTileLinkNetworkPort_18_14135_io_manager_release_ready),
    .io_manager_release_valid(ManagerTileLinkNetworkPort_18_14135_io_manager_release_valid),
    .io_manager_release_bits_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_beat),
    .io_manager_release_bits_addr_block(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_block),
    .io_manager_release_bits_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_xact_id),
    .io_manager_release_bits_voluntary(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_voluntary),
    .io_manager_release_bits_r_type(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_r_type),
    .io_manager_release_bits_data(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_data),
    .io_manager_release_bits_client_id(ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_id),
    .io_network_acquire_ready(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_ready),
    .io_network_acquire_valid(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_valid),
    .io_network_acquire_bits_header_src(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_src),
    .io_network_acquire_bits_header_dst(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_dst),
    .io_network_acquire_bits_payload_addr_block(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_block),
    .io_network_acquire_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_client_xact_id),
    .io_network_acquire_bits_payload_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_beat),
    .io_network_acquire_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_is_builtin_type),
    .io_network_acquire_bits_payload_a_type(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_a_type),
    .io_network_acquire_bits_payload_union(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_union),
    .io_network_acquire_bits_payload_data(ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_data),
    .io_network_grant_ready(ManagerTileLinkNetworkPort_18_14135_io_network_grant_ready),
    .io_network_grant_valid(ManagerTileLinkNetworkPort_18_14135_io_network_grant_valid),
    .io_network_grant_bits_header_src(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_src),
    .io_network_grant_bits_header_dst(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_dst),
    .io_network_grant_bits_payload_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_addr_beat),
    .io_network_grant_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_client_xact_id),
    .io_network_grant_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_manager_xact_id),
    .io_network_grant_bits_payload_is_builtin_type(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_is_builtin_type),
    .io_network_grant_bits_payload_g_type(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_g_type),
    .io_network_grant_bits_payload_data(ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_data),
    .io_network_finish_ready(ManagerTileLinkNetworkPort_18_14135_io_network_finish_ready),
    .io_network_finish_valid(ManagerTileLinkNetworkPort_18_14135_io_network_finish_valid),
    .io_network_finish_bits_header_src(ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_src),
    .io_network_finish_bits_header_dst(ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_dst),
    .io_network_finish_bits_payload_manager_xact_id(ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_payload_manager_xact_id),
    .io_network_probe_ready(ManagerTileLinkNetworkPort_18_14135_io_network_probe_ready),
    .io_network_probe_valid(ManagerTileLinkNetworkPort_18_14135_io_network_probe_valid),
    .io_network_probe_bits_header_src(ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_src),
    .io_network_probe_bits_header_dst(ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_dst),
    .io_network_probe_bits_payload_addr_block(ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_addr_block),
    .io_network_probe_bits_payload_p_type(ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_p_type),
    .io_network_release_ready(ManagerTileLinkNetworkPort_18_14135_io_network_release_ready),
    .io_network_release_valid(ManagerTileLinkNetworkPort_18_14135_io_network_release_valid),
    .io_network_release_bits_header_src(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_src),
    .io_network_release_bits_header_dst(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_dst),
    .io_network_release_bits_payload_addr_beat(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_beat),
    .io_network_release_bits_payload_addr_block(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_block),
    .io_network_release_bits_payload_client_xact_id(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_client_xact_id),
    .io_network_release_bits_payload_voluntary(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_voluntary),
    .io_network_release_bits_payload_r_type(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_r_type),
    .io_network_release_bits_payload_data(ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_data)
  );
  TileLinkEnqueuer_17 TileLinkEnqueuer_19_14136 (
    .clk(TileLinkEnqueuer_19_14136_clk),
    .reset(TileLinkEnqueuer_19_14136_reset),
    .io_client_acquire_ready(TileLinkEnqueuer_19_14136_io_client_acquire_ready),
    .io_client_acquire_valid(TileLinkEnqueuer_19_14136_io_client_acquire_valid),
    .io_client_acquire_bits_header_src(TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_src),
    .io_client_acquire_bits_header_dst(TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_dst),
    .io_client_acquire_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_block),
    .io_client_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_client_xact_id),
    .io_client_acquire_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_beat),
    .io_client_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_is_builtin_type),
    .io_client_acquire_bits_payload_a_type(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_a_type),
    .io_client_acquire_bits_payload_union(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_union),
    .io_client_acquire_bits_payload_data(TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_data),
    .io_client_grant_ready(TileLinkEnqueuer_19_14136_io_client_grant_ready),
    .io_client_grant_valid(TileLinkEnqueuer_19_14136_io_client_grant_valid),
    .io_client_grant_bits_header_src(TileLinkEnqueuer_19_14136_io_client_grant_bits_header_src),
    .io_client_grant_bits_header_dst(TileLinkEnqueuer_19_14136_io_client_grant_bits_header_dst),
    .io_client_grant_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_addr_beat),
    .io_client_grant_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_client_xact_id),
    .io_client_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_manager_xact_id),
    .io_client_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_is_builtin_type),
    .io_client_grant_bits_payload_g_type(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_g_type),
    .io_client_grant_bits_payload_data(TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_data),
    .io_client_finish_ready(TileLinkEnqueuer_19_14136_io_client_finish_ready),
    .io_client_finish_valid(TileLinkEnqueuer_19_14136_io_client_finish_valid),
    .io_client_finish_bits_header_src(TileLinkEnqueuer_19_14136_io_client_finish_bits_header_src),
    .io_client_finish_bits_header_dst(TileLinkEnqueuer_19_14136_io_client_finish_bits_header_dst),
    .io_client_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_19_14136_io_client_finish_bits_payload_manager_xact_id),
    .io_client_probe_ready(TileLinkEnqueuer_19_14136_io_client_probe_ready),
    .io_client_probe_valid(TileLinkEnqueuer_19_14136_io_client_probe_valid),
    .io_client_probe_bits_header_src(TileLinkEnqueuer_19_14136_io_client_probe_bits_header_src),
    .io_client_probe_bits_header_dst(TileLinkEnqueuer_19_14136_io_client_probe_bits_header_dst),
    .io_client_probe_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_addr_block),
    .io_client_probe_bits_payload_p_type(TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_p_type),
    .io_client_release_ready(TileLinkEnqueuer_19_14136_io_client_release_ready),
    .io_client_release_valid(TileLinkEnqueuer_19_14136_io_client_release_valid),
    .io_client_release_bits_header_src(TileLinkEnqueuer_19_14136_io_client_release_bits_header_src),
    .io_client_release_bits_header_dst(TileLinkEnqueuer_19_14136_io_client_release_bits_header_dst),
    .io_client_release_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_beat),
    .io_client_release_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_block),
    .io_client_release_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_client_xact_id),
    .io_client_release_bits_payload_voluntary(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_voluntary),
    .io_client_release_bits_payload_r_type(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_r_type),
    .io_client_release_bits_payload_data(TileLinkEnqueuer_19_14136_io_client_release_bits_payload_data),
    .io_manager_acquire_ready(TileLinkEnqueuer_19_14136_io_manager_acquire_ready),
    .io_manager_acquire_valid(TileLinkEnqueuer_19_14136_io_manager_acquire_valid),
    .io_manager_acquire_bits_header_src(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_src),
    .io_manager_acquire_bits_header_dst(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_dst),
    .io_manager_acquire_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_block),
    .io_manager_acquire_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_client_xact_id),
    .io_manager_acquire_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_beat),
    .io_manager_acquire_bits_payload_is_builtin_type(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_is_builtin_type),
    .io_manager_acquire_bits_payload_a_type(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_a_type),
    .io_manager_acquire_bits_payload_union(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_union),
    .io_manager_acquire_bits_payload_data(TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_data),
    .io_manager_grant_ready(TileLinkEnqueuer_19_14136_io_manager_grant_ready),
    .io_manager_grant_valid(TileLinkEnqueuer_19_14136_io_manager_grant_valid),
    .io_manager_grant_bits_header_src(TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_src),
    .io_manager_grant_bits_header_dst(TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_dst),
    .io_manager_grant_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_addr_beat),
    .io_manager_grant_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_client_xact_id),
    .io_manager_grant_bits_payload_manager_xact_id(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_manager_xact_id),
    .io_manager_grant_bits_payload_is_builtin_type(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_is_builtin_type),
    .io_manager_grant_bits_payload_g_type(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_g_type),
    .io_manager_grant_bits_payload_data(TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_data),
    .io_manager_finish_ready(TileLinkEnqueuer_19_14136_io_manager_finish_ready),
    .io_manager_finish_valid(TileLinkEnqueuer_19_14136_io_manager_finish_valid),
    .io_manager_finish_bits_header_src(TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_src),
    .io_manager_finish_bits_header_dst(TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_dst),
    .io_manager_finish_bits_payload_manager_xact_id(TileLinkEnqueuer_19_14136_io_manager_finish_bits_payload_manager_xact_id),
    .io_manager_probe_ready(TileLinkEnqueuer_19_14136_io_manager_probe_ready),
    .io_manager_probe_valid(TileLinkEnqueuer_19_14136_io_manager_probe_valid),
    .io_manager_probe_bits_header_src(TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_src),
    .io_manager_probe_bits_header_dst(TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_dst),
    .io_manager_probe_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_addr_block),
    .io_manager_probe_bits_payload_p_type(TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_p_type),
    .io_manager_release_ready(TileLinkEnqueuer_19_14136_io_manager_release_ready),
    .io_manager_release_valid(TileLinkEnqueuer_19_14136_io_manager_release_valid),
    .io_manager_release_bits_header_src(TileLinkEnqueuer_19_14136_io_manager_release_bits_header_src),
    .io_manager_release_bits_header_dst(TileLinkEnqueuer_19_14136_io_manager_release_bits_header_dst),
    .io_manager_release_bits_payload_addr_beat(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_beat),
    .io_manager_release_bits_payload_addr_block(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_block),
    .io_manager_release_bits_payload_client_xact_id(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_client_xact_id),
    .io_manager_release_bits_payload_voluntary(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_voluntary),
    .io_manager_release_bits_payload_r_type(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_r_type),
    .io_manager_release_bits_payload_data(TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_data)
  );
  BasicBus acqNet (
    .clk(acqNet_clk),
    .reset(acqNet_reset),
    .io_in_0_ready(acqNet_io_in_0_ready),
    .io_in_0_valid(acqNet_io_in_0_valid),
    .io_in_0_bits_header_src(acqNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(acqNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(acqNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(acqNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_addr_beat(acqNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_is_builtin_type(acqNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_a_type(acqNet_io_in_0_bits_payload_a_type),
    .io_in_0_bits_payload_union(acqNet_io_in_0_bits_payload_union),
    .io_in_0_bits_payload_data(acqNet_io_in_0_bits_payload_data),
    .io_in_1_ready(acqNet_io_in_1_ready),
    .io_in_1_valid(acqNet_io_in_1_valid),
    .io_in_1_bits_header_src(acqNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(acqNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(acqNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(acqNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_addr_beat(acqNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_is_builtin_type(acqNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_a_type(acqNet_io_in_1_bits_payload_a_type),
    .io_in_1_bits_payload_union(acqNet_io_in_1_bits_payload_union),
    .io_in_1_bits_payload_data(acqNet_io_in_1_bits_payload_data),
    .io_in_2_ready(acqNet_io_in_2_ready),
    .io_in_2_valid(acqNet_io_in_2_valid),
    .io_in_2_bits_header_src(acqNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(acqNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(acqNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(acqNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_addr_beat(acqNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_is_builtin_type(acqNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_a_type(acqNet_io_in_2_bits_payload_a_type),
    .io_in_2_bits_payload_union(acqNet_io_in_2_bits_payload_union),
    .io_in_2_bits_payload_data(acqNet_io_in_2_bits_payload_data),
    .io_in_3_ready(acqNet_io_in_3_ready),
    .io_in_3_valid(acqNet_io_in_3_valid),
    .io_in_3_bits_header_src(acqNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(acqNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(acqNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(acqNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_addr_beat(acqNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_is_builtin_type(acqNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_a_type(acqNet_io_in_3_bits_payload_a_type),
    .io_in_3_bits_payload_union(acqNet_io_in_3_bits_payload_union),
    .io_in_3_bits_payload_data(acqNet_io_in_3_bits_payload_data),
    .io_in_4_ready(acqNet_io_in_4_ready),
    .io_in_4_valid(acqNet_io_in_4_valid),
    .io_in_4_bits_header_src(acqNet_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(acqNet_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_block(acqNet_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_client_xact_id(acqNet_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_addr_beat(acqNet_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_is_builtin_type(acqNet_io_in_4_bits_payload_is_builtin_type),
    .io_in_4_bits_payload_a_type(acqNet_io_in_4_bits_payload_a_type),
    .io_in_4_bits_payload_union(acqNet_io_in_4_bits_payload_union),
    .io_in_4_bits_payload_data(acqNet_io_in_4_bits_payload_data),
    .io_out_0_ready(acqNet_io_out_0_ready),
    .io_out_0_valid(acqNet_io_out_0_valid),
    .io_out_0_bits_header_src(acqNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(acqNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(acqNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(acqNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_addr_beat(acqNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_is_builtin_type(acqNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_a_type(acqNet_io_out_0_bits_payload_a_type),
    .io_out_0_bits_payload_union(acqNet_io_out_0_bits_payload_union),
    .io_out_0_bits_payload_data(acqNet_io_out_0_bits_payload_data),
    .io_out_1_ready(acqNet_io_out_1_ready),
    .io_out_1_valid(acqNet_io_out_1_valid),
    .io_out_1_bits_header_src(acqNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(acqNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(acqNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(acqNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_addr_beat(acqNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_is_builtin_type(acqNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_a_type(acqNet_io_out_1_bits_payload_a_type),
    .io_out_1_bits_payload_union(acqNet_io_out_1_bits_payload_union),
    .io_out_1_bits_payload_data(acqNet_io_out_1_bits_payload_data),
    .io_out_2_ready(acqNet_io_out_2_ready),
    .io_out_2_valid(acqNet_io_out_2_valid),
    .io_out_2_bits_header_src(acqNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(acqNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(acqNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(acqNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_addr_beat(acqNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_is_builtin_type(acqNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_a_type(acqNet_io_out_2_bits_payload_a_type),
    .io_out_2_bits_payload_union(acqNet_io_out_2_bits_payload_union),
    .io_out_2_bits_payload_data(acqNet_io_out_2_bits_payload_data),
    .io_out_3_ready(acqNet_io_out_3_ready),
    .io_out_3_valid(acqNet_io_out_3_valid),
    .io_out_3_bits_header_src(acqNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(acqNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(acqNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(acqNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_addr_beat(acqNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_is_builtin_type(acqNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_a_type(acqNet_io_out_3_bits_payload_a_type),
    .io_out_3_bits_payload_union(acqNet_io_out_3_bits_payload_union),
    .io_out_3_bits_payload_data(acqNet_io_out_3_bits_payload_data),
    .io_out_4_ready(acqNet_io_out_4_ready),
    .io_out_4_valid(acqNet_io_out_4_valid),
    .io_out_4_bits_header_src(acqNet_io_out_4_bits_header_src),
    .io_out_4_bits_header_dst(acqNet_io_out_4_bits_header_dst),
    .io_out_4_bits_payload_addr_block(acqNet_io_out_4_bits_payload_addr_block),
    .io_out_4_bits_payload_client_xact_id(acqNet_io_out_4_bits_payload_client_xact_id),
    .io_out_4_bits_payload_addr_beat(acqNet_io_out_4_bits_payload_addr_beat),
    .io_out_4_bits_payload_is_builtin_type(acqNet_io_out_4_bits_payload_is_builtin_type),
    .io_out_4_bits_payload_a_type(acqNet_io_out_4_bits_payload_a_type),
    .io_out_4_bits_payload_union(acqNet_io_out_4_bits_payload_union),
    .io_out_4_bits_payload_data(acqNet_io_out_4_bits_payload_data)
  );
  BasicBus_20 relNet (
    .clk(relNet_clk),
    .reset(relNet_reset),
    .io_in_0_ready(relNet_io_in_0_ready),
    .io_in_0_valid(relNet_io_in_0_valid),
    .io_in_0_bits_header_src(relNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(relNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(relNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_addr_block(relNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_client_xact_id(relNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_voluntary(relNet_io_in_0_bits_payload_voluntary),
    .io_in_0_bits_payload_r_type(relNet_io_in_0_bits_payload_r_type),
    .io_in_0_bits_payload_data(relNet_io_in_0_bits_payload_data),
    .io_in_1_ready(relNet_io_in_1_ready),
    .io_in_1_valid(relNet_io_in_1_valid),
    .io_in_1_bits_header_src(relNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(relNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(relNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_addr_block(relNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_client_xact_id(relNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_voluntary(relNet_io_in_1_bits_payload_voluntary),
    .io_in_1_bits_payload_r_type(relNet_io_in_1_bits_payload_r_type),
    .io_in_1_bits_payload_data(relNet_io_in_1_bits_payload_data),
    .io_in_2_ready(relNet_io_in_2_ready),
    .io_in_2_valid(relNet_io_in_2_valid),
    .io_in_2_bits_header_src(relNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(relNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(relNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_addr_block(relNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_client_xact_id(relNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_voluntary(relNet_io_in_2_bits_payload_voluntary),
    .io_in_2_bits_payload_r_type(relNet_io_in_2_bits_payload_r_type),
    .io_in_2_bits_payload_data(relNet_io_in_2_bits_payload_data),
    .io_in_3_ready(relNet_io_in_3_ready),
    .io_in_3_valid(relNet_io_in_3_valid),
    .io_in_3_bits_header_src(relNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(relNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(relNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_addr_block(relNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_client_xact_id(relNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_voluntary(relNet_io_in_3_bits_payload_voluntary),
    .io_in_3_bits_payload_r_type(relNet_io_in_3_bits_payload_r_type),
    .io_in_3_bits_payload_data(relNet_io_in_3_bits_payload_data),
    .io_in_4_ready(relNet_io_in_4_ready),
    .io_in_4_valid(relNet_io_in_4_valid),
    .io_in_4_bits_header_src(relNet_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(relNet_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_beat(relNet_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_addr_block(relNet_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_client_xact_id(relNet_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_voluntary(relNet_io_in_4_bits_payload_voluntary),
    .io_in_4_bits_payload_r_type(relNet_io_in_4_bits_payload_r_type),
    .io_in_4_bits_payload_data(relNet_io_in_4_bits_payload_data),
    .io_out_0_ready(relNet_io_out_0_ready),
    .io_out_0_valid(relNet_io_out_0_valid),
    .io_out_0_bits_header_src(relNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(relNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(relNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_addr_block(relNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_client_xact_id(relNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_voluntary(relNet_io_out_0_bits_payload_voluntary),
    .io_out_0_bits_payload_r_type(relNet_io_out_0_bits_payload_r_type),
    .io_out_0_bits_payload_data(relNet_io_out_0_bits_payload_data),
    .io_out_1_ready(relNet_io_out_1_ready),
    .io_out_1_valid(relNet_io_out_1_valid),
    .io_out_1_bits_header_src(relNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(relNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(relNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_addr_block(relNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_client_xact_id(relNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_voluntary(relNet_io_out_1_bits_payload_voluntary),
    .io_out_1_bits_payload_r_type(relNet_io_out_1_bits_payload_r_type),
    .io_out_1_bits_payload_data(relNet_io_out_1_bits_payload_data),
    .io_out_2_ready(relNet_io_out_2_ready),
    .io_out_2_valid(relNet_io_out_2_valid),
    .io_out_2_bits_header_src(relNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(relNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(relNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_addr_block(relNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_client_xact_id(relNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_voluntary(relNet_io_out_2_bits_payload_voluntary),
    .io_out_2_bits_payload_r_type(relNet_io_out_2_bits_payload_r_type),
    .io_out_2_bits_payload_data(relNet_io_out_2_bits_payload_data),
    .io_out_3_ready(relNet_io_out_3_ready),
    .io_out_3_valid(relNet_io_out_3_valid),
    .io_out_3_bits_header_src(relNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(relNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(relNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_addr_block(relNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_client_xact_id(relNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_voluntary(relNet_io_out_3_bits_payload_voluntary),
    .io_out_3_bits_payload_r_type(relNet_io_out_3_bits_payload_r_type),
    .io_out_3_bits_payload_data(relNet_io_out_3_bits_payload_data),
    .io_out_4_ready(relNet_io_out_4_ready),
    .io_out_4_valid(relNet_io_out_4_valid),
    .io_out_4_bits_header_src(relNet_io_out_4_bits_header_src),
    .io_out_4_bits_header_dst(relNet_io_out_4_bits_header_dst),
    .io_out_4_bits_payload_addr_beat(relNet_io_out_4_bits_payload_addr_beat),
    .io_out_4_bits_payload_addr_block(relNet_io_out_4_bits_payload_addr_block),
    .io_out_4_bits_payload_client_xact_id(relNet_io_out_4_bits_payload_client_xact_id),
    .io_out_4_bits_payload_voluntary(relNet_io_out_4_bits_payload_voluntary),
    .io_out_4_bits_payload_r_type(relNet_io_out_4_bits_payload_r_type),
    .io_out_4_bits_payload_data(relNet_io_out_4_bits_payload_data)
  );
  BasicBus_22 prbNet (
    .clk(prbNet_clk),
    .reset(prbNet_reset),
    .io_in_0_ready(prbNet_io_in_0_ready),
    .io_in_0_valid(prbNet_io_in_0_valid),
    .io_in_0_bits_header_src(prbNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(prbNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_block(prbNet_io_in_0_bits_payload_addr_block),
    .io_in_0_bits_payload_p_type(prbNet_io_in_0_bits_payload_p_type),
    .io_in_1_ready(prbNet_io_in_1_ready),
    .io_in_1_valid(prbNet_io_in_1_valid),
    .io_in_1_bits_header_src(prbNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(prbNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_block(prbNet_io_in_1_bits_payload_addr_block),
    .io_in_1_bits_payload_p_type(prbNet_io_in_1_bits_payload_p_type),
    .io_in_2_ready(prbNet_io_in_2_ready),
    .io_in_2_valid(prbNet_io_in_2_valid),
    .io_in_2_bits_header_src(prbNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(prbNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_block(prbNet_io_in_2_bits_payload_addr_block),
    .io_in_2_bits_payload_p_type(prbNet_io_in_2_bits_payload_p_type),
    .io_in_3_ready(prbNet_io_in_3_ready),
    .io_in_3_valid(prbNet_io_in_3_valid),
    .io_in_3_bits_header_src(prbNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(prbNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_block(prbNet_io_in_3_bits_payload_addr_block),
    .io_in_3_bits_payload_p_type(prbNet_io_in_3_bits_payload_p_type),
    .io_in_4_ready(prbNet_io_in_4_ready),
    .io_in_4_valid(prbNet_io_in_4_valid),
    .io_in_4_bits_header_src(prbNet_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(prbNet_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_block(prbNet_io_in_4_bits_payload_addr_block),
    .io_in_4_bits_payload_p_type(prbNet_io_in_4_bits_payload_p_type),
    .io_out_0_ready(prbNet_io_out_0_ready),
    .io_out_0_valid(prbNet_io_out_0_valid),
    .io_out_0_bits_header_src(prbNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(prbNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_block(prbNet_io_out_0_bits_payload_addr_block),
    .io_out_0_bits_payload_p_type(prbNet_io_out_0_bits_payload_p_type),
    .io_out_1_ready(prbNet_io_out_1_ready),
    .io_out_1_valid(prbNet_io_out_1_valid),
    .io_out_1_bits_header_src(prbNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(prbNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_block(prbNet_io_out_1_bits_payload_addr_block),
    .io_out_1_bits_payload_p_type(prbNet_io_out_1_bits_payload_p_type),
    .io_out_2_ready(prbNet_io_out_2_ready),
    .io_out_2_valid(prbNet_io_out_2_valid),
    .io_out_2_bits_header_src(prbNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(prbNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_block(prbNet_io_out_2_bits_payload_addr_block),
    .io_out_2_bits_payload_p_type(prbNet_io_out_2_bits_payload_p_type),
    .io_out_3_ready(prbNet_io_out_3_ready),
    .io_out_3_valid(prbNet_io_out_3_valid),
    .io_out_3_bits_header_src(prbNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(prbNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_block(prbNet_io_out_3_bits_payload_addr_block),
    .io_out_3_bits_payload_p_type(prbNet_io_out_3_bits_payload_p_type),
    .io_out_4_ready(prbNet_io_out_4_ready),
    .io_out_4_valid(prbNet_io_out_4_valid),
    .io_out_4_bits_header_src(prbNet_io_out_4_bits_header_src),
    .io_out_4_bits_header_dst(prbNet_io_out_4_bits_header_dst),
    .io_out_4_bits_payload_addr_block(prbNet_io_out_4_bits_payload_addr_block),
    .io_out_4_bits_payload_p_type(prbNet_io_out_4_bits_payload_p_type)
  );
  BasicBus_24 gntNet (
    .clk(gntNet_clk),
    .reset(gntNet_reset),
    .io_in_0_ready(gntNet_io_in_0_ready),
    .io_in_0_valid(gntNet_io_in_0_valid),
    .io_in_0_bits_header_src(gntNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(gntNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_addr_beat(gntNet_io_in_0_bits_payload_addr_beat),
    .io_in_0_bits_payload_client_xact_id(gntNet_io_in_0_bits_payload_client_xact_id),
    .io_in_0_bits_payload_manager_xact_id(gntNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_0_bits_payload_is_builtin_type(gntNet_io_in_0_bits_payload_is_builtin_type),
    .io_in_0_bits_payload_g_type(gntNet_io_in_0_bits_payload_g_type),
    .io_in_0_bits_payload_data(gntNet_io_in_0_bits_payload_data),
    .io_in_1_ready(gntNet_io_in_1_ready),
    .io_in_1_valid(gntNet_io_in_1_valid),
    .io_in_1_bits_header_src(gntNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(gntNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_addr_beat(gntNet_io_in_1_bits_payload_addr_beat),
    .io_in_1_bits_payload_client_xact_id(gntNet_io_in_1_bits_payload_client_xact_id),
    .io_in_1_bits_payload_manager_xact_id(gntNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_1_bits_payload_is_builtin_type(gntNet_io_in_1_bits_payload_is_builtin_type),
    .io_in_1_bits_payload_g_type(gntNet_io_in_1_bits_payload_g_type),
    .io_in_1_bits_payload_data(gntNet_io_in_1_bits_payload_data),
    .io_in_2_ready(gntNet_io_in_2_ready),
    .io_in_2_valid(gntNet_io_in_2_valid),
    .io_in_2_bits_header_src(gntNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(gntNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_addr_beat(gntNet_io_in_2_bits_payload_addr_beat),
    .io_in_2_bits_payload_client_xact_id(gntNet_io_in_2_bits_payload_client_xact_id),
    .io_in_2_bits_payload_manager_xact_id(gntNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_2_bits_payload_is_builtin_type(gntNet_io_in_2_bits_payload_is_builtin_type),
    .io_in_2_bits_payload_g_type(gntNet_io_in_2_bits_payload_g_type),
    .io_in_2_bits_payload_data(gntNet_io_in_2_bits_payload_data),
    .io_in_3_ready(gntNet_io_in_3_ready),
    .io_in_3_valid(gntNet_io_in_3_valid),
    .io_in_3_bits_header_src(gntNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(gntNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_addr_beat(gntNet_io_in_3_bits_payload_addr_beat),
    .io_in_3_bits_payload_client_xact_id(gntNet_io_in_3_bits_payload_client_xact_id),
    .io_in_3_bits_payload_manager_xact_id(gntNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_3_bits_payload_is_builtin_type(gntNet_io_in_3_bits_payload_is_builtin_type),
    .io_in_3_bits_payload_g_type(gntNet_io_in_3_bits_payload_g_type),
    .io_in_3_bits_payload_data(gntNet_io_in_3_bits_payload_data),
    .io_in_4_ready(gntNet_io_in_4_ready),
    .io_in_4_valid(gntNet_io_in_4_valid),
    .io_in_4_bits_header_src(gntNet_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(gntNet_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_addr_beat(gntNet_io_in_4_bits_payload_addr_beat),
    .io_in_4_bits_payload_client_xact_id(gntNet_io_in_4_bits_payload_client_xact_id),
    .io_in_4_bits_payload_manager_xact_id(gntNet_io_in_4_bits_payload_manager_xact_id),
    .io_in_4_bits_payload_is_builtin_type(gntNet_io_in_4_bits_payload_is_builtin_type),
    .io_in_4_bits_payload_g_type(gntNet_io_in_4_bits_payload_g_type),
    .io_in_4_bits_payload_data(gntNet_io_in_4_bits_payload_data),
    .io_out_0_ready(gntNet_io_out_0_ready),
    .io_out_0_valid(gntNet_io_out_0_valid),
    .io_out_0_bits_header_src(gntNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(gntNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_addr_beat(gntNet_io_out_0_bits_payload_addr_beat),
    .io_out_0_bits_payload_client_xact_id(gntNet_io_out_0_bits_payload_client_xact_id),
    .io_out_0_bits_payload_manager_xact_id(gntNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_0_bits_payload_is_builtin_type(gntNet_io_out_0_bits_payload_is_builtin_type),
    .io_out_0_bits_payload_g_type(gntNet_io_out_0_bits_payload_g_type),
    .io_out_0_bits_payload_data(gntNet_io_out_0_bits_payload_data),
    .io_out_1_ready(gntNet_io_out_1_ready),
    .io_out_1_valid(gntNet_io_out_1_valid),
    .io_out_1_bits_header_src(gntNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(gntNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_addr_beat(gntNet_io_out_1_bits_payload_addr_beat),
    .io_out_1_bits_payload_client_xact_id(gntNet_io_out_1_bits_payload_client_xact_id),
    .io_out_1_bits_payload_manager_xact_id(gntNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_1_bits_payload_is_builtin_type(gntNet_io_out_1_bits_payload_is_builtin_type),
    .io_out_1_bits_payload_g_type(gntNet_io_out_1_bits_payload_g_type),
    .io_out_1_bits_payload_data(gntNet_io_out_1_bits_payload_data),
    .io_out_2_ready(gntNet_io_out_2_ready),
    .io_out_2_valid(gntNet_io_out_2_valid),
    .io_out_2_bits_header_src(gntNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(gntNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_addr_beat(gntNet_io_out_2_bits_payload_addr_beat),
    .io_out_2_bits_payload_client_xact_id(gntNet_io_out_2_bits_payload_client_xact_id),
    .io_out_2_bits_payload_manager_xact_id(gntNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_2_bits_payload_is_builtin_type(gntNet_io_out_2_bits_payload_is_builtin_type),
    .io_out_2_bits_payload_g_type(gntNet_io_out_2_bits_payload_g_type),
    .io_out_2_bits_payload_data(gntNet_io_out_2_bits_payload_data),
    .io_out_3_ready(gntNet_io_out_3_ready),
    .io_out_3_valid(gntNet_io_out_3_valid),
    .io_out_3_bits_header_src(gntNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(gntNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_addr_beat(gntNet_io_out_3_bits_payload_addr_beat),
    .io_out_3_bits_payload_client_xact_id(gntNet_io_out_3_bits_payload_client_xact_id),
    .io_out_3_bits_payload_manager_xact_id(gntNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_3_bits_payload_is_builtin_type(gntNet_io_out_3_bits_payload_is_builtin_type),
    .io_out_3_bits_payload_g_type(gntNet_io_out_3_bits_payload_g_type),
    .io_out_3_bits_payload_data(gntNet_io_out_3_bits_payload_data),
    .io_out_4_ready(gntNet_io_out_4_ready),
    .io_out_4_valid(gntNet_io_out_4_valid),
    .io_out_4_bits_header_src(gntNet_io_out_4_bits_header_src),
    .io_out_4_bits_header_dst(gntNet_io_out_4_bits_header_dst),
    .io_out_4_bits_payload_addr_beat(gntNet_io_out_4_bits_payload_addr_beat),
    .io_out_4_bits_payload_client_xact_id(gntNet_io_out_4_bits_payload_client_xact_id),
    .io_out_4_bits_payload_manager_xact_id(gntNet_io_out_4_bits_payload_manager_xact_id),
    .io_out_4_bits_payload_is_builtin_type(gntNet_io_out_4_bits_payload_is_builtin_type),
    .io_out_4_bits_payload_g_type(gntNet_io_out_4_bits_payload_g_type),
    .io_out_4_bits_payload_data(gntNet_io_out_4_bits_payload_data)
  );
  BasicBus_26 ackNet (
    .clk(ackNet_clk),
    .reset(ackNet_reset),
    .io_in_0_ready(ackNet_io_in_0_ready),
    .io_in_0_valid(ackNet_io_in_0_valid),
    .io_in_0_bits_header_src(ackNet_io_in_0_bits_header_src),
    .io_in_0_bits_header_dst(ackNet_io_in_0_bits_header_dst),
    .io_in_0_bits_payload_manager_xact_id(ackNet_io_in_0_bits_payload_manager_xact_id),
    .io_in_1_ready(ackNet_io_in_1_ready),
    .io_in_1_valid(ackNet_io_in_1_valid),
    .io_in_1_bits_header_src(ackNet_io_in_1_bits_header_src),
    .io_in_1_bits_header_dst(ackNet_io_in_1_bits_header_dst),
    .io_in_1_bits_payload_manager_xact_id(ackNet_io_in_1_bits_payload_manager_xact_id),
    .io_in_2_ready(ackNet_io_in_2_ready),
    .io_in_2_valid(ackNet_io_in_2_valid),
    .io_in_2_bits_header_src(ackNet_io_in_2_bits_header_src),
    .io_in_2_bits_header_dst(ackNet_io_in_2_bits_header_dst),
    .io_in_2_bits_payload_manager_xact_id(ackNet_io_in_2_bits_payload_manager_xact_id),
    .io_in_3_ready(ackNet_io_in_3_ready),
    .io_in_3_valid(ackNet_io_in_3_valid),
    .io_in_3_bits_header_src(ackNet_io_in_3_bits_header_src),
    .io_in_3_bits_header_dst(ackNet_io_in_3_bits_header_dst),
    .io_in_3_bits_payload_manager_xact_id(ackNet_io_in_3_bits_payload_manager_xact_id),
    .io_in_4_ready(ackNet_io_in_4_ready),
    .io_in_4_valid(ackNet_io_in_4_valid),
    .io_in_4_bits_header_src(ackNet_io_in_4_bits_header_src),
    .io_in_4_bits_header_dst(ackNet_io_in_4_bits_header_dst),
    .io_in_4_bits_payload_manager_xact_id(ackNet_io_in_4_bits_payload_manager_xact_id),
    .io_out_0_ready(ackNet_io_out_0_ready),
    .io_out_0_valid(ackNet_io_out_0_valid),
    .io_out_0_bits_header_src(ackNet_io_out_0_bits_header_src),
    .io_out_0_bits_header_dst(ackNet_io_out_0_bits_header_dst),
    .io_out_0_bits_payload_manager_xact_id(ackNet_io_out_0_bits_payload_manager_xact_id),
    .io_out_1_ready(ackNet_io_out_1_ready),
    .io_out_1_valid(ackNet_io_out_1_valid),
    .io_out_1_bits_header_src(ackNet_io_out_1_bits_header_src),
    .io_out_1_bits_header_dst(ackNet_io_out_1_bits_header_dst),
    .io_out_1_bits_payload_manager_xact_id(ackNet_io_out_1_bits_payload_manager_xact_id),
    .io_out_2_ready(ackNet_io_out_2_ready),
    .io_out_2_valid(ackNet_io_out_2_valid),
    .io_out_2_bits_header_src(ackNet_io_out_2_bits_header_src),
    .io_out_2_bits_header_dst(ackNet_io_out_2_bits_header_dst),
    .io_out_2_bits_payload_manager_xact_id(ackNet_io_out_2_bits_payload_manager_xact_id),
    .io_out_3_ready(ackNet_io_out_3_ready),
    .io_out_3_valid(ackNet_io_out_3_valid),
    .io_out_3_bits_header_src(ackNet_io_out_3_bits_header_src),
    .io_out_3_bits_header_dst(ackNet_io_out_3_bits_header_dst),
    .io_out_3_bits_payload_manager_xact_id(ackNet_io_out_3_bits_payload_manager_xact_id),
    .io_out_4_ready(ackNet_io_out_4_ready),
    .io_out_4_valid(ackNet_io_out_4_valid),
    .io_out_4_bits_header_src(ackNet_io_out_4_bits_header_src),
    .io_out_4_bits_header_dst(ackNet_io_out_4_bits_header_dst),
    .io_out_4_bits_payload_manager_xact_id(ackNet_io_out_4_bits_payload_manager_xact_id)
  );
  assign io_clients_cached_0_acquire_ready = ClientTileLinkNetworkPort_14128_io_client_acquire_ready;
  assign io_clients_cached_0_probe_valid = ClientTileLinkNetworkPort_14128_io_client_probe_valid;
  assign io_clients_cached_0_probe_bits_addr_block = ClientTileLinkNetworkPort_14128_io_client_probe_bits_addr_block;
  assign io_clients_cached_0_probe_bits_p_type = ClientTileLinkNetworkPort_14128_io_client_probe_bits_p_type;
  assign io_clients_cached_0_release_ready = ClientTileLinkNetworkPort_14128_io_client_release_ready;
  assign io_clients_cached_0_grant_valid = ClientTileLinkNetworkPort_14128_io_client_grant_valid;
  assign io_clients_cached_0_grant_bits_addr_beat = ClientTileLinkNetworkPort_14128_io_client_grant_bits_addr_beat;
  assign io_clients_cached_0_grant_bits_client_xact_id = ClientTileLinkNetworkPort_14128_io_client_grant_bits_client_xact_id;
  assign io_clients_cached_0_grant_bits_manager_xact_id = ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_xact_id;
  assign io_clients_cached_0_grant_bits_is_builtin_type = ClientTileLinkNetworkPort_14128_io_client_grant_bits_is_builtin_type;
  assign io_clients_cached_0_grant_bits_g_type = ClientTileLinkNetworkPort_14128_io_client_grant_bits_g_type;
  assign io_clients_cached_0_grant_bits_data = ClientTileLinkNetworkPort_14128_io_client_grant_bits_data;
  assign io_clients_cached_0_grant_bits_manager_id = ClientTileLinkNetworkPort_14128_io_client_grant_bits_manager_id;
  assign io_clients_cached_0_finish_ready = ClientTileLinkNetworkPort_14128_io_client_finish_ready;
  assign io_clients_uncached_0_acquire_ready = ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_ready;
  assign io_clients_uncached_0_grant_valid = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_valid;
  assign io_clients_uncached_0_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_0_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_0_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_0_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_0_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_g_type;
  assign io_clients_uncached_0_grant_bits_data = ClientUncachedTileLinkNetworkPort_14130_io_client_grant_bits_data;
  assign io_clients_uncached_1_acquire_ready = ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_ready;
  assign io_clients_uncached_1_grant_valid = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_valid;
  assign io_clients_uncached_1_grant_bits_addr_beat = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_addr_beat;
  assign io_clients_uncached_1_grant_bits_client_xact_id = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_client_xact_id;
  assign io_clients_uncached_1_grant_bits_manager_xact_id = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_manager_xact_id;
  assign io_clients_uncached_1_grant_bits_is_builtin_type = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_is_builtin_type;
  assign io_clients_uncached_1_grant_bits_g_type = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_g_type;
  assign io_clients_uncached_1_grant_bits_data = ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_bits_data;
  assign io_managers_0_acquire_valid = ManagerTileLinkNetworkPort_14133_io_manager_acquire_valid;
  assign io_managers_0_acquire_bits_addr_block = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_block;
  assign io_managers_0_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_xact_id;
  assign io_managers_0_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_addr_beat;
  assign io_managers_0_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_0_acquire_bits_a_type = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_a_type;
  assign io_managers_0_acquire_bits_union = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_union;
  assign io_managers_0_acquire_bits_data = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_data;
  assign io_managers_0_acquire_bits_client_id = ManagerTileLinkNetworkPort_14133_io_manager_acquire_bits_client_id;
  assign io_managers_0_grant_ready = ManagerTileLinkNetworkPort_14133_io_manager_grant_ready;
  assign io_managers_0_finish_valid = ManagerTileLinkNetworkPort_14133_io_manager_finish_valid;
  assign io_managers_0_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_14133_io_manager_finish_bits_manager_xact_id;
  assign io_managers_0_probe_ready = ManagerTileLinkNetworkPort_14133_io_manager_probe_ready;
  assign io_managers_0_release_valid = ManagerTileLinkNetworkPort_14133_io_manager_release_valid;
  assign io_managers_0_release_bits_addr_beat = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_beat;
  assign io_managers_0_release_bits_addr_block = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_addr_block;
  assign io_managers_0_release_bits_client_xact_id = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_xact_id;
  assign io_managers_0_release_bits_voluntary = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_voluntary;
  assign io_managers_0_release_bits_r_type = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_r_type;
  assign io_managers_0_release_bits_data = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_data;
  assign io_managers_0_release_bits_client_id = ManagerTileLinkNetworkPort_14133_io_manager_release_bits_client_id;
  assign io_managers_1_acquire_valid = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_valid;
  assign io_managers_1_acquire_bits_addr_block = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_block;
  assign io_managers_1_acquire_bits_client_xact_id = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_xact_id;
  assign io_managers_1_acquire_bits_addr_beat = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_addr_beat;
  assign io_managers_1_acquire_bits_is_builtin_type = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_is_builtin_type;
  assign io_managers_1_acquire_bits_a_type = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_a_type;
  assign io_managers_1_acquire_bits_union = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_union;
  assign io_managers_1_acquire_bits_data = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_data;
  assign io_managers_1_acquire_bits_client_id = ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_bits_client_id;
  assign io_managers_1_grant_ready = ManagerTileLinkNetworkPort_18_14135_io_manager_grant_ready;
  assign io_managers_1_finish_valid = ManagerTileLinkNetworkPort_18_14135_io_manager_finish_valid;
  assign io_managers_1_finish_bits_manager_xact_id = ManagerTileLinkNetworkPort_18_14135_io_manager_finish_bits_manager_xact_id;
  assign io_managers_1_probe_ready = ManagerTileLinkNetworkPort_18_14135_io_manager_probe_ready;
  assign io_managers_1_release_valid = ManagerTileLinkNetworkPort_18_14135_io_manager_release_valid;
  assign io_managers_1_release_bits_addr_beat = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_beat;
  assign io_managers_1_release_bits_addr_block = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_addr_block;
  assign io_managers_1_release_bits_client_xact_id = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_xact_id;
  assign io_managers_1_release_bits_voluntary = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_voluntary;
  assign io_managers_1_release_bits_r_type = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_r_type;
  assign io_managers_1_release_bits_data = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_data;
  assign io_managers_1_release_bits_client_id = ManagerTileLinkNetworkPort_18_14135_io_manager_release_bits_client_id;
  assign TileLinkEnqueuer_14127_clk = clk;
  assign TileLinkEnqueuer_14127_reset = reset;
  assign TileLinkEnqueuer_14127_io_client_acquire_valid = ClientTileLinkNetworkPort_14128_io_network_acquire_valid;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_header_src = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_header_dst = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_block = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_client_xact_id = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_addr_beat = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_is_builtin_type = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_a_type = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_union = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_14127_io_client_acquire_bits_payload_data = ClientTileLinkNetworkPort_14128_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_14127_io_client_grant_ready = ClientTileLinkNetworkPort_14128_io_network_grant_ready;
  assign TileLinkEnqueuer_14127_io_client_finish_valid = ClientTileLinkNetworkPort_14128_io_network_finish_valid;
  assign TileLinkEnqueuer_14127_io_client_finish_bits_header_src = ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_14127_io_client_finish_bits_header_dst = ClientTileLinkNetworkPort_14128_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_14127_io_client_finish_bits_payload_manager_xact_id = ClientTileLinkNetworkPort_14128_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_14127_io_client_probe_ready = ClientTileLinkNetworkPort_14128_io_network_probe_ready;
  assign TileLinkEnqueuer_14127_io_client_release_valid = ClientTileLinkNetworkPort_14128_io_network_release_valid;
  assign TileLinkEnqueuer_14127_io_client_release_bits_header_src = ClientTileLinkNetworkPort_14128_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_14127_io_client_release_bits_header_dst = ClientTileLinkNetworkPort_14128_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_beat = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_addr_block = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_client_xact_id = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_voluntary = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_r_type = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_14127_io_client_release_bits_payload_data = ClientTileLinkNetworkPort_14128_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_14127_io_manager_acquire_ready = T_15723_ready;
  assign TileLinkEnqueuer_14127_io_manager_grant_valid = T_20911_valid;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_header_src = T_20911_bits_header_src;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_header_dst = T_20911_bits_header_dst;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_addr_beat = T_20911_bits_payload_addr_beat;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_client_xact_id = T_20911_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_manager_xact_id = T_20911_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_is_builtin_type = T_20911_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_g_type = T_20911_bits_payload_g_type;
  assign TileLinkEnqueuer_14127_io_manager_grant_bits_payload_data = T_20911_bits_payload_data;
  assign TileLinkEnqueuer_14127_io_manager_finish_ready = T_23770_ready;
  assign TileLinkEnqueuer_14127_io_manager_probe_valid = T_18679_valid;
  assign TileLinkEnqueuer_14127_io_manager_probe_bits_header_src = T_18679_bits_header_src;
  assign TileLinkEnqueuer_14127_io_manager_probe_bits_header_dst = T_18679_bits_header_dst;
  assign TileLinkEnqueuer_14127_io_manager_probe_bits_payload_addr_block = T_18679_bits_payload_addr_block;
  assign TileLinkEnqueuer_14127_io_manager_probe_bits_payload_p_type = T_18679_bits_payload_p_type;
  assign TileLinkEnqueuer_14127_io_manager_release_ready = T_17555_ready;
  assign ClientTileLinkNetworkPort_14128_clk = clk;
  assign ClientTileLinkNetworkPort_14128_reset = reset;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_valid = io_clients_cached_0_acquire_valid;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_block = io_clients_cached_0_acquire_bits_addr_block;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_client_xact_id = io_clients_cached_0_acquire_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_addr_beat = io_clients_cached_0_acquire_bits_addr_beat;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_is_builtin_type = io_clients_cached_0_acquire_bits_is_builtin_type;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_a_type = io_clients_cached_0_acquire_bits_a_type;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_union = io_clients_cached_0_acquire_bits_union;
  assign ClientTileLinkNetworkPort_14128_io_client_acquire_bits_data = io_clients_cached_0_acquire_bits_data;
  assign ClientTileLinkNetworkPort_14128_io_client_probe_ready = io_clients_cached_0_probe_ready;
  assign ClientTileLinkNetworkPort_14128_io_client_release_valid = io_clients_cached_0_release_valid;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_beat = io_clients_cached_0_release_bits_addr_beat;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_addr_block = io_clients_cached_0_release_bits_addr_block;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_client_xact_id = io_clients_cached_0_release_bits_client_xact_id;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_voluntary = io_clients_cached_0_release_bits_voluntary;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_r_type = io_clients_cached_0_release_bits_r_type;
  assign ClientTileLinkNetworkPort_14128_io_client_release_bits_data = io_clients_cached_0_release_bits_data;
  assign ClientTileLinkNetworkPort_14128_io_client_grant_ready = io_clients_cached_0_grant_ready;
  assign ClientTileLinkNetworkPort_14128_io_client_finish_valid = io_clients_cached_0_finish_valid;
  assign ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_xact_id = io_clients_cached_0_finish_bits_manager_xact_id;
  assign ClientTileLinkNetworkPort_14128_io_client_finish_bits_manager_id = io_clients_cached_0_finish_bits_manager_id;
  assign ClientTileLinkNetworkPort_14128_io_network_acquire_ready = TileLinkEnqueuer_14127_io_client_acquire_ready;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_valid = TileLinkEnqueuer_14127_io_client_grant_valid;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_src = TileLinkEnqueuer_14127_io_client_grant_bits_header_src;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_header_dst = TileLinkEnqueuer_14127_io_client_grant_bits_header_dst;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_14127_io_client_grant_bits_payload_addr_beat;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_14127_io_client_grant_bits_payload_client_xact_id;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_14127_io_client_grant_bits_payload_manager_xact_id;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_14127_io_client_grant_bits_payload_is_builtin_type;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_14127_io_client_grant_bits_payload_g_type;
  assign ClientTileLinkNetworkPort_14128_io_network_grant_bits_payload_data = TileLinkEnqueuer_14127_io_client_grant_bits_payload_data;
  assign ClientTileLinkNetworkPort_14128_io_network_finish_ready = TileLinkEnqueuer_14127_io_client_finish_ready;
  assign ClientTileLinkNetworkPort_14128_io_network_probe_valid = TileLinkEnqueuer_14127_io_client_probe_valid;
  assign ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_src = TileLinkEnqueuer_14127_io_client_probe_bits_header_src;
  assign ClientTileLinkNetworkPort_14128_io_network_probe_bits_header_dst = TileLinkEnqueuer_14127_io_client_probe_bits_header_dst;
  assign ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_14127_io_client_probe_bits_payload_addr_block;
  assign ClientTileLinkNetworkPort_14128_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_14127_io_client_probe_bits_payload_p_type;
  assign ClientTileLinkNetworkPort_14128_io_network_release_ready = TileLinkEnqueuer_14127_io_client_release_ready;
  assign TileLinkEnqueuer_4_14129_clk = clk;
  assign TileLinkEnqueuer_4_14129_reset = reset;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_valid;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_4_14129_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_4_14129_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_14130_io_network_grant_ready;
  assign TileLinkEnqueuer_4_14129_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_14130_io_network_finish_valid;
  assign TileLinkEnqueuer_4_14129_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_4_14129_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_4_14129_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_14130_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_14129_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_14130_io_network_probe_ready;
  assign TileLinkEnqueuer_4_14129_io_client_release_valid = ClientUncachedTileLinkNetworkPort_14130_io_network_release_valid;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_4_14129_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_14130_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_4_14129_io_manager_acquire_ready = T_15908_ready;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_valid = T_21551_valid;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_src = T_21551_bits_header_src;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_header_dst = T_21551_bits_header_dst;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_addr_beat = T_21551_bits_payload_addr_beat;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_client_xact_id = T_21551_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_manager_xact_id = T_21551_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_is_builtin_type = T_21551_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_g_type = T_21551_bits_payload_g_type;
  assign TileLinkEnqueuer_4_14129_io_manager_grant_bits_payload_data = T_21551_bits_payload_data;
  assign TileLinkEnqueuer_4_14129_io_manager_finish_ready = T_23925_ready;
  assign TileLinkEnqueuer_4_14129_io_manager_probe_valid = T_19299_valid;
  assign TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_src = T_19299_bits_header_src;
  assign TileLinkEnqueuer_4_14129_io_manager_probe_bits_header_dst = T_19299_bits_header_dst;
  assign TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_addr_block = T_19299_bits_payload_addr_block;
  assign TileLinkEnqueuer_4_14129_io_manager_probe_bits_payload_p_type = T_19299_bits_payload_p_type;
  assign TileLinkEnqueuer_4_14129_io_manager_release_ready = T_17735_ready;
  assign ClientUncachedTileLinkNetworkPort_14130_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_14130_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_valid = io_clients_uncached_0_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_block = io_clients_uncached_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_client_xact_id = io_clients_uncached_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_addr_beat = io_clients_uncached_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_is_builtin_type = io_clients_uncached_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_a_type = io_clients_uncached_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_union = io_clients_uncached_0_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_acquire_bits_data = io_clients_uncached_0_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_14130_io_client_grant_ready = io_clients_uncached_0_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_acquire_ready = TileLinkEnqueuer_4_14129_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_valid = TileLinkEnqueuer_4_14129_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_src = TileLinkEnqueuer_4_14129_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_header_dst = TileLinkEnqueuer_4_14129_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_grant_bits_payload_data = TileLinkEnqueuer_4_14129_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_finish_ready = TileLinkEnqueuer_4_14129_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_probe_valid = TileLinkEnqueuer_4_14129_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_src = TileLinkEnqueuer_4_14129_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_header_dst = TileLinkEnqueuer_4_14129_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_4_14129_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_14130_io_network_release_ready = TileLinkEnqueuer_4_14129_io_client_release_ready;
  assign TileLinkEnqueuer_9_14131_clk = clk;
  assign TileLinkEnqueuer_9_14131_reset = reset;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_valid = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_valid;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_src = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_src;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_header_dst = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_header_dst;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_block;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_addr_beat;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_is_builtin_type = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_a_type = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_a_type;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_union = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_union;
  assign TileLinkEnqueuer_9_14131_io_client_acquire_bits_payload_data = ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_bits_payload_data;
  assign TileLinkEnqueuer_9_14131_io_client_grant_ready = ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_ready;
  assign TileLinkEnqueuer_9_14131_io_client_finish_valid = ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_valid;
  assign TileLinkEnqueuer_9_14131_io_client_finish_bits_header_src = ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_src;
  assign TileLinkEnqueuer_9_14131_io_client_finish_bits_header_dst = ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_header_dst;
  assign TileLinkEnqueuer_9_14131_io_client_finish_bits_payload_manager_xact_id = ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_9_14131_io_client_probe_ready = ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_ready;
  assign TileLinkEnqueuer_9_14131_io_client_release_valid = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_valid;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_header_src = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_src;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_header_dst = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_header_dst;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_beat = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_beat;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_addr_block = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_addr_block;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_client_xact_id = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_voluntary = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_voluntary;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_r_type = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_r_type;
  assign TileLinkEnqueuer_9_14131_io_client_release_bits_payload_data = ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_bits_payload_data;
  assign TileLinkEnqueuer_9_14131_io_manager_acquire_ready = T_16093_ready;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_valid = T_22191_valid;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_src = T_22191_bits_header_src;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_header_dst = T_22191_bits_header_dst;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_addr_beat = T_22191_bits_payload_addr_beat;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_client_xact_id = T_22191_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_manager_xact_id = T_22191_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_is_builtin_type = T_22191_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_g_type = T_22191_bits_payload_g_type;
  assign TileLinkEnqueuer_9_14131_io_manager_grant_bits_payload_data = T_22191_bits_payload_data;
  assign TileLinkEnqueuer_9_14131_io_manager_finish_ready = T_24080_ready;
  assign TileLinkEnqueuer_9_14131_io_manager_probe_valid = T_19919_valid;
  assign TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_src = T_19919_bits_header_src;
  assign TileLinkEnqueuer_9_14131_io_manager_probe_bits_header_dst = T_19919_bits_header_dst;
  assign TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_addr_block = T_19919_bits_payload_addr_block;
  assign TileLinkEnqueuer_9_14131_io_manager_probe_bits_payload_p_type = T_19919_bits_payload_p_type;
  assign TileLinkEnqueuer_9_14131_io_manager_release_ready = T_17915_ready;
  assign ClientUncachedTileLinkNetworkPort_14_14132_clk = clk;
  assign ClientUncachedTileLinkNetworkPort_14_14132_reset = reset;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_valid = io_clients_uncached_1_acquire_valid;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_block = io_clients_uncached_1_acquire_bits_addr_block;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_client_xact_id = io_clients_uncached_1_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_addr_beat = io_clients_uncached_1_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_is_builtin_type = io_clients_uncached_1_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_a_type = io_clients_uncached_1_acquire_bits_a_type;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_union = io_clients_uncached_1_acquire_bits_union;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_acquire_bits_data = io_clients_uncached_1_acquire_bits_data;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_client_grant_ready = io_clients_uncached_1_grant_ready;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_acquire_ready = TileLinkEnqueuer_9_14131_io_client_acquire_ready;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_valid = TileLinkEnqueuer_9_14131_io_client_grant_valid;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_src = TileLinkEnqueuer_9_14131_io_client_grant_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_header_dst = TileLinkEnqueuer_9_14131_io_client_grant_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_addr_beat = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_addr_beat;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_client_xact_id = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_client_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_manager_xact_id = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_manager_xact_id;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_is_builtin_type = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_is_builtin_type;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_g_type = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_g_type;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_grant_bits_payload_data = TileLinkEnqueuer_9_14131_io_client_grant_bits_payload_data;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_finish_ready = TileLinkEnqueuer_9_14131_io_client_finish_ready;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_valid = TileLinkEnqueuer_9_14131_io_client_probe_valid;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_src = TileLinkEnqueuer_9_14131_io_client_probe_bits_header_src;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_header_dst = TileLinkEnqueuer_9_14131_io_client_probe_bits_header_dst;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_addr_block = TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_addr_block;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_probe_bits_payload_p_type = TileLinkEnqueuer_9_14131_io_client_probe_bits_payload_p_type;
  assign ClientUncachedTileLinkNetworkPort_14_14132_io_network_release_ready = TileLinkEnqueuer_9_14131_io_client_release_ready;
  assign ManagerTileLinkNetworkPort_14133_clk = clk;
  assign ManagerTileLinkNetworkPort_14133_reset = reset;
  assign ManagerTileLinkNetworkPort_14133_io_manager_acquire_ready = io_managers_0_acquire_ready;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_valid = io_managers_0_grant_valid;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_addr_beat = io_managers_0_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_xact_id = io_managers_0_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_manager_xact_id = io_managers_0_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_is_builtin_type = io_managers_0_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_g_type = io_managers_0_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_data = io_managers_0_grant_bits_data;
  assign ManagerTileLinkNetworkPort_14133_io_manager_grant_bits_client_id = io_managers_0_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_14133_io_manager_finish_ready = io_managers_0_finish_ready;
  assign ManagerTileLinkNetworkPort_14133_io_manager_probe_valid = io_managers_0_probe_valid;
  assign ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_addr_block = io_managers_0_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_p_type = io_managers_0_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_14133_io_manager_probe_bits_client_id = io_managers_0_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_14133_io_manager_release_ready = io_managers_0_release_ready;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_valid = TileLinkEnqueuer_17_14134_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_src = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_header_dst = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_union = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_14133_io_network_acquire_bits_payload_data = TileLinkEnqueuer_17_14134_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_14133_io_network_grant_ready = TileLinkEnqueuer_17_14134_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_14133_io_network_finish_valid = TileLinkEnqueuer_17_14134_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_src = TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_14133_io_network_finish_bits_header_dst = TileLinkEnqueuer_17_14134_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_14133_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_17_14134_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_14133_io_network_probe_ready = TileLinkEnqueuer_17_14134_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_valid = TileLinkEnqueuer_17_14134_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_src = TileLinkEnqueuer_17_14134_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_header_dst = TileLinkEnqueuer_17_14134_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_r_type = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_14133_io_network_release_bits_payload_data = TileLinkEnqueuer_17_14134_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_17_14134_clk = clk;
  assign TileLinkEnqueuer_17_14134_reset = reset;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_valid = T_14709_valid;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_src = T_14709_bits_header_src;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_header_dst = T_14709_bits_header_dst;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_block = T_14709_bits_payload_addr_block;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_client_xact_id = T_14709_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_addr_beat = T_14709_bits_payload_addr_beat;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_is_builtin_type = T_14709_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_a_type = T_14709_bits_payload_a_type;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_union = T_14709_bits_payload_union;
  assign TileLinkEnqueuer_17_14134_io_client_acquire_bits_payload_data = T_14709_bits_payload_data;
  assign TileLinkEnqueuer_17_14134_io_client_grant_ready = T_20275_ready;
  assign TileLinkEnqueuer_17_14134_io_client_finish_valid = T_22816_valid;
  assign TileLinkEnqueuer_17_14134_io_client_finish_bits_header_src = T_22816_bits_header_src;
  assign TileLinkEnqueuer_17_14134_io_client_finish_bits_header_dst = T_22816_bits_header_dst;
  assign TileLinkEnqueuer_17_14134_io_client_finish_bits_payload_manager_xact_id = T_22816_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_17_14134_io_client_probe_ready = T_18083_ready;
  assign TileLinkEnqueuer_17_14134_io_client_release_valid = T_16551_valid;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_header_src = T_16551_bits_header_src;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_header_dst = T_16551_bits_header_dst;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_beat = T_16551_bits_payload_addr_beat;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_addr_block = T_16551_bits_payload_addr_block;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_client_xact_id = T_16551_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_voluntary = T_16551_bits_payload_voluntary;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_r_type = T_16551_bits_payload_r_type;
  assign TileLinkEnqueuer_17_14134_io_client_release_bits_payload_data = T_16551_bits_payload_data;
  assign TileLinkEnqueuer_17_14134_io_manager_acquire_ready = ManagerTileLinkNetworkPort_14133_io_network_acquire_ready;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_valid = ManagerTileLinkNetworkPort_14133_io_network_grant_valid;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_17_14134_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_14133_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_17_14134_io_manager_finish_ready = ManagerTileLinkNetworkPort_14133_io_network_finish_ready;
  assign TileLinkEnqueuer_17_14134_io_manager_probe_valid = ManagerTileLinkNetworkPort_14133_io_network_probe_valid;
  assign TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_17_14134_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_14133_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_17_14134_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_14133_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_17_14134_io_manager_release_ready = ManagerTileLinkNetworkPort_14133_io_network_release_ready;
  assign ManagerTileLinkNetworkPort_18_14135_clk = clk;
  assign ManagerTileLinkNetworkPort_18_14135_reset = reset;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_acquire_ready = io_managers_1_acquire_ready;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_valid = io_managers_1_grant_valid;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_addr_beat = io_managers_1_grant_bits_addr_beat;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_xact_id = io_managers_1_grant_bits_client_xact_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_manager_xact_id = io_managers_1_grant_bits_manager_xact_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_is_builtin_type = io_managers_1_grant_bits_is_builtin_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_g_type = io_managers_1_grant_bits_g_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_data = io_managers_1_grant_bits_data;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_grant_bits_client_id = io_managers_1_grant_bits_client_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_finish_ready = io_managers_1_finish_ready;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_probe_valid = io_managers_1_probe_valid;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_addr_block = io_managers_1_probe_bits_addr_block;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_p_type = io_managers_1_probe_bits_p_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_probe_bits_client_id = io_managers_1_probe_bits_client_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_manager_release_ready = io_managers_1_release_ready;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_valid = TileLinkEnqueuer_19_14136_io_manager_acquire_valid;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_src = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_src;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_header_dst = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_header_dst;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_block = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_client_xact_id = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_addr_beat = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_is_builtin_type = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_is_builtin_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_a_type = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_a_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_union = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_union;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_acquire_bits_payload_data = TileLinkEnqueuer_19_14136_io_manager_acquire_bits_payload_data;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_grant_ready = TileLinkEnqueuer_19_14136_io_manager_grant_ready;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_finish_valid = TileLinkEnqueuer_19_14136_io_manager_finish_valid;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_src = TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_src;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_header_dst = TileLinkEnqueuer_19_14136_io_manager_finish_bits_header_dst;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_finish_bits_payload_manager_xact_id = TileLinkEnqueuer_19_14136_io_manager_finish_bits_payload_manager_xact_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_probe_ready = TileLinkEnqueuer_19_14136_io_manager_probe_ready;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_valid = TileLinkEnqueuer_19_14136_io_manager_release_valid;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_src = TileLinkEnqueuer_19_14136_io_manager_release_bits_header_src;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_header_dst = TileLinkEnqueuer_19_14136_io_manager_release_bits_header_dst;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_beat = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_beat;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_addr_block = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_addr_block;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_client_xact_id = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_client_xact_id;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_voluntary = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_voluntary;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_r_type = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_r_type;
  assign ManagerTileLinkNetworkPort_18_14135_io_network_release_bits_payload_data = TileLinkEnqueuer_19_14136_io_manager_release_bits_payload_data;
  assign TileLinkEnqueuer_19_14136_clk = clk;
  assign TileLinkEnqueuer_19_14136_reset = reset;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_valid = T_15354_valid;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_src = T_15354_bits_header_src;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_header_dst = T_15354_bits_header_dst;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_block = T_15354_bits_payload_addr_block;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_client_xact_id = T_15354_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_addr_beat = T_15354_bits_payload_addr_beat;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_is_builtin_type = T_15354_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_a_type = T_15354_bits_payload_a_type;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_union = T_15354_bits_payload_union;
  assign TileLinkEnqueuer_19_14136_io_client_acquire_bits_payload_data = T_15354_bits_payload_data;
  assign TileLinkEnqueuer_19_14136_io_client_grant_ready = T_20455_ready;
  assign TileLinkEnqueuer_19_14136_io_client_finish_valid = T_23431_valid;
  assign TileLinkEnqueuer_19_14136_io_client_finish_bits_header_src = T_23431_bits_header_src;
  assign TileLinkEnqueuer_19_14136_io_client_finish_bits_header_dst = T_23431_bits_header_dst;
  assign TileLinkEnqueuer_19_14136_io_client_finish_bits_payload_manager_xact_id = T_23431_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_19_14136_io_client_probe_ready = T_18243_ready;
  assign TileLinkEnqueuer_19_14136_io_client_release_valid = T_17191_valid;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_header_src = T_17191_bits_header_src;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_header_dst = T_17191_bits_header_dst;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_beat = T_17191_bits_payload_addr_beat;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_addr_block = T_17191_bits_payload_addr_block;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_client_xact_id = T_17191_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_voluntary = T_17191_bits_payload_voluntary;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_r_type = T_17191_bits_payload_r_type;
  assign TileLinkEnqueuer_19_14136_io_client_release_bits_payload_data = T_17191_bits_payload_data;
  assign TileLinkEnqueuer_19_14136_io_manager_acquire_ready = ManagerTileLinkNetworkPort_18_14135_io_network_acquire_ready;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_valid = ManagerTileLinkNetworkPort_18_14135_io_network_grant_valid;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_src = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_src;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_header_dst = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_header_dst;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_addr_beat = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_addr_beat;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_client_xact_id = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_client_xact_id;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_manager_xact_id = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_manager_xact_id;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_is_builtin_type = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_is_builtin_type;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_g_type = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_g_type;
  assign TileLinkEnqueuer_19_14136_io_manager_grant_bits_payload_data = ManagerTileLinkNetworkPort_18_14135_io_network_grant_bits_payload_data;
  assign TileLinkEnqueuer_19_14136_io_manager_finish_ready = ManagerTileLinkNetworkPort_18_14135_io_network_finish_ready;
  assign TileLinkEnqueuer_19_14136_io_manager_probe_valid = ManagerTileLinkNetworkPort_18_14135_io_network_probe_valid;
  assign TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_src = ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_src;
  assign TileLinkEnqueuer_19_14136_io_manager_probe_bits_header_dst = ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_header_dst;
  assign TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_addr_block = ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_addr_block;
  assign TileLinkEnqueuer_19_14136_io_manager_probe_bits_payload_p_type = ManagerTileLinkNetworkPort_18_14135_io_network_probe_bits_payload_p_type;
  assign TileLinkEnqueuer_19_14136_io_manager_release_ready = ManagerTileLinkNetworkPort_18_14135_io_network_release_ready;
  assign acqNet_clk = clk;
  assign acqNet_reset = reset;
  assign acqNet_io_in_0_valid = 1'h0;
  assign acqNet_io_in_0_bits_header_src = GEN_1;
  assign acqNet_io_in_0_bits_header_dst = GEN_2;
  assign acqNet_io_in_0_bits_payload_addr_block = GEN_3;
  assign acqNet_io_in_0_bits_payload_client_xact_id = GEN_4;
  assign acqNet_io_in_0_bits_payload_addr_beat = GEN_5;
  assign acqNet_io_in_0_bits_payload_is_builtin_type = GEN_6;
  assign acqNet_io_in_0_bits_payload_a_type = GEN_7;
  assign acqNet_io_in_0_bits_payload_union = GEN_8;
  assign acqNet_io_in_0_bits_payload_data = GEN_9;
  assign acqNet_io_in_1_valid = 1'h0;
  assign acqNet_io_in_1_bits_header_src = GEN_10;
  assign acqNet_io_in_1_bits_header_dst = GEN_11;
  assign acqNet_io_in_1_bits_payload_addr_block = GEN_12;
  assign acqNet_io_in_1_bits_payload_client_xact_id = GEN_13;
  assign acqNet_io_in_1_bits_payload_addr_beat = GEN_14;
  assign acqNet_io_in_1_bits_payload_is_builtin_type = GEN_15;
  assign acqNet_io_in_1_bits_payload_a_type = GEN_16;
  assign acqNet_io_in_1_bits_payload_union = GEN_17;
  assign acqNet_io_in_1_bits_payload_data = GEN_18;
  assign acqNet_io_in_2_valid = T_15723_valid;
  assign acqNet_io_in_2_bits_header_src = T_15723_bits_header_src;
  assign acqNet_io_in_2_bits_header_dst = T_15723_bits_header_dst;
  assign acqNet_io_in_2_bits_payload_addr_block = T_15723_bits_payload_addr_block;
  assign acqNet_io_in_2_bits_payload_client_xact_id = T_15723_bits_payload_client_xact_id;
  assign acqNet_io_in_2_bits_payload_addr_beat = T_15723_bits_payload_addr_beat;
  assign acqNet_io_in_2_bits_payload_is_builtin_type = T_15723_bits_payload_is_builtin_type;
  assign acqNet_io_in_2_bits_payload_a_type = T_15723_bits_payload_a_type;
  assign acqNet_io_in_2_bits_payload_union = T_15723_bits_payload_union;
  assign acqNet_io_in_2_bits_payload_data = T_15723_bits_payload_data;
  assign acqNet_io_in_3_valid = T_15908_valid;
  assign acqNet_io_in_3_bits_header_src = T_15908_bits_header_src;
  assign acqNet_io_in_3_bits_header_dst = T_15908_bits_header_dst;
  assign acqNet_io_in_3_bits_payload_addr_block = T_15908_bits_payload_addr_block;
  assign acqNet_io_in_3_bits_payload_client_xact_id = T_15908_bits_payload_client_xact_id;
  assign acqNet_io_in_3_bits_payload_addr_beat = T_15908_bits_payload_addr_beat;
  assign acqNet_io_in_3_bits_payload_is_builtin_type = T_15908_bits_payload_is_builtin_type;
  assign acqNet_io_in_3_bits_payload_a_type = T_15908_bits_payload_a_type;
  assign acqNet_io_in_3_bits_payload_union = T_15908_bits_payload_union;
  assign acqNet_io_in_3_bits_payload_data = T_15908_bits_payload_data;
  assign acqNet_io_in_4_valid = T_16093_valid;
  assign acqNet_io_in_4_bits_header_src = T_16093_bits_header_src;
  assign acqNet_io_in_4_bits_header_dst = T_16093_bits_header_dst;
  assign acqNet_io_in_4_bits_payload_addr_block = T_16093_bits_payload_addr_block;
  assign acqNet_io_in_4_bits_payload_client_xact_id = T_16093_bits_payload_client_xact_id;
  assign acqNet_io_in_4_bits_payload_addr_beat = T_16093_bits_payload_addr_beat;
  assign acqNet_io_in_4_bits_payload_is_builtin_type = T_16093_bits_payload_is_builtin_type;
  assign acqNet_io_in_4_bits_payload_a_type = T_16093_bits_payload_a_type;
  assign acqNet_io_in_4_bits_payload_union = T_16093_bits_payload_union;
  assign acqNet_io_in_4_bits_payload_data = T_16093_bits_payload_data;
  assign acqNet_io_out_0_ready = T_14709_ready;
  assign acqNet_io_out_1_ready = T_15354_ready;
  assign acqNet_io_out_2_ready = 1'h0;
  assign acqNet_io_out_3_ready = 1'h0;
  assign acqNet_io_out_4_ready = 1'h0;
  assign relNet_clk = clk;
  assign relNet_reset = reset;
  assign relNet_io_in_0_valid = 1'h0;
  assign relNet_io_in_0_bits_header_src = GEN_19;
  assign relNet_io_in_0_bits_header_dst = GEN_20;
  assign relNet_io_in_0_bits_payload_addr_beat = GEN_21;
  assign relNet_io_in_0_bits_payload_addr_block = GEN_22;
  assign relNet_io_in_0_bits_payload_client_xact_id = GEN_23;
  assign relNet_io_in_0_bits_payload_voluntary = GEN_24;
  assign relNet_io_in_0_bits_payload_r_type = GEN_25;
  assign relNet_io_in_0_bits_payload_data = GEN_26;
  assign relNet_io_in_1_valid = 1'h0;
  assign relNet_io_in_1_bits_header_src = GEN_27;
  assign relNet_io_in_1_bits_header_dst = GEN_28;
  assign relNet_io_in_1_bits_payload_addr_beat = GEN_29;
  assign relNet_io_in_1_bits_payload_addr_block = GEN_30;
  assign relNet_io_in_1_bits_payload_client_xact_id = GEN_31;
  assign relNet_io_in_1_bits_payload_voluntary = GEN_32;
  assign relNet_io_in_1_bits_payload_r_type = GEN_33;
  assign relNet_io_in_1_bits_payload_data = GEN_34;
  assign relNet_io_in_2_valid = T_17555_valid;
  assign relNet_io_in_2_bits_header_src = T_17555_bits_header_src;
  assign relNet_io_in_2_bits_header_dst = T_17555_bits_header_dst;
  assign relNet_io_in_2_bits_payload_addr_beat = T_17555_bits_payload_addr_beat;
  assign relNet_io_in_2_bits_payload_addr_block = T_17555_bits_payload_addr_block;
  assign relNet_io_in_2_bits_payload_client_xact_id = T_17555_bits_payload_client_xact_id;
  assign relNet_io_in_2_bits_payload_voluntary = T_17555_bits_payload_voluntary;
  assign relNet_io_in_2_bits_payload_r_type = T_17555_bits_payload_r_type;
  assign relNet_io_in_2_bits_payload_data = T_17555_bits_payload_data;
  assign relNet_io_in_3_valid = T_17735_valid;
  assign relNet_io_in_3_bits_header_src = T_17735_bits_header_src;
  assign relNet_io_in_3_bits_header_dst = T_17735_bits_header_dst;
  assign relNet_io_in_3_bits_payload_addr_beat = T_17735_bits_payload_addr_beat;
  assign relNet_io_in_3_bits_payload_addr_block = T_17735_bits_payload_addr_block;
  assign relNet_io_in_3_bits_payload_client_xact_id = T_17735_bits_payload_client_xact_id;
  assign relNet_io_in_3_bits_payload_voluntary = T_17735_bits_payload_voluntary;
  assign relNet_io_in_3_bits_payload_r_type = T_17735_bits_payload_r_type;
  assign relNet_io_in_3_bits_payload_data = T_17735_bits_payload_data;
  assign relNet_io_in_4_valid = T_17915_valid;
  assign relNet_io_in_4_bits_header_src = T_17915_bits_header_src;
  assign relNet_io_in_4_bits_header_dst = T_17915_bits_header_dst;
  assign relNet_io_in_4_bits_payload_addr_beat = T_17915_bits_payload_addr_beat;
  assign relNet_io_in_4_bits_payload_addr_block = T_17915_bits_payload_addr_block;
  assign relNet_io_in_4_bits_payload_client_xact_id = T_17915_bits_payload_client_xact_id;
  assign relNet_io_in_4_bits_payload_voluntary = T_17915_bits_payload_voluntary;
  assign relNet_io_in_4_bits_payload_r_type = T_17915_bits_payload_r_type;
  assign relNet_io_in_4_bits_payload_data = T_17915_bits_payload_data;
  assign relNet_io_out_0_ready = T_16551_ready;
  assign relNet_io_out_1_ready = T_17191_ready;
  assign relNet_io_out_2_ready = 1'h0;
  assign relNet_io_out_3_ready = 1'h0;
  assign relNet_io_out_4_ready = 1'h0;
  assign prbNet_clk = clk;
  assign prbNet_reset = reset;
  assign prbNet_io_in_0_valid = T_18083_valid;
  assign prbNet_io_in_0_bits_header_src = T_18083_bits_header_src;
  assign prbNet_io_in_0_bits_header_dst = T_18083_bits_header_dst;
  assign prbNet_io_in_0_bits_payload_addr_block = T_18083_bits_payload_addr_block;
  assign prbNet_io_in_0_bits_payload_p_type = T_18083_bits_payload_p_type;
  assign prbNet_io_in_1_valid = T_18243_valid;
  assign prbNet_io_in_1_bits_header_src = T_18243_bits_header_src;
  assign prbNet_io_in_1_bits_header_dst = T_18243_bits_header_dst;
  assign prbNet_io_in_1_bits_payload_addr_block = T_18243_bits_payload_addr_block;
  assign prbNet_io_in_1_bits_payload_p_type = T_18243_bits_payload_p_type;
  assign prbNet_io_in_2_valid = 1'h0;
  assign prbNet_io_in_2_bits_header_src = GEN_35;
  assign prbNet_io_in_2_bits_header_dst = GEN_36;
  assign prbNet_io_in_2_bits_payload_addr_block = GEN_37;
  assign prbNet_io_in_2_bits_payload_p_type = GEN_38;
  assign prbNet_io_in_3_valid = 1'h0;
  assign prbNet_io_in_3_bits_header_src = GEN_39;
  assign prbNet_io_in_3_bits_header_dst = GEN_40;
  assign prbNet_io_in_3_bits_payload_addr_block = GEN_41;
  assign prbNet_io_in_3_bits_payload_p_type = GEN_42;
  assign prbNet_io_in_4_valid = 1'h0;
  assign prbNet_io_in_4_bits_header_src = GEN_43;
  assign prbNet_io_in_4_bits_header_dst = GEN_44;
  assign prbNet_io_in_4_bits_payload_addr_block = GEN_45;
  assign prbNet_io_in_4_bits_payload_p_type = GEN_46;
  assign prbNet_io_out_0_ready = 1'h0;
  assign prbNet_io_out_1_ready = 1'h0;
  assign prbNet_io_out_2_ready = T_18679_ready;
  assign prbNet_io_out_3_ready = T_19299_ready;
  assign prbNet_io_out_4_ready = T_19919_ready;
  assign gntNet_clk = clk;
  assign gntNet_reset = reset;
  assign gntNet_io_in_0_valid = T_20275_valid;
  assign gntNet_io_in_0_bits_header_src = T_20275_bits_header_src;
  assign gntNet_io_in_0_bits_header_dst = T_20275_bits_header_dst;
  assign gntNet_io_in_0_bits_payload_addr_beat = T_20275_bits_payload_addr_beat;
  assign gntNet_io_in_0_bits_payload_client_xact_id = T_20275_bits_payload_client_xact_id;
  assign gntNet_io_in_0_bits_payload_manager_xact_id = T_20275_bits_payload_manager_xact_id;
  assign gntNet_io_in_0_bits_payload_is_builtin_type = T_20275_bits_payload_is_builtin_type;
  assign gntNet_io_in_0_bits_payload_g_type = T_20275_bits_payload_g_type;
  assign gntNet_io_in_0_bits_payload_data = T_20275_bits_payload_data;
  assign gntNet_io_in_1_valid = T_20455_valid;
  assign gntNet_io_in_1_bits_header_src = T_20455_bits_header_src;
  assign gntNet_io_in_1_bits_header_dst = T_20455_bits_header_dst;
  assign gntNet_io_in_1_bits_payload_addr_beat = T_20455_bits_payload_addr_beat;
  assign gntNet_io_in_1_bits_payload_client_xact_id = T_20455_bits_payload_client_xact_id;
  assign gntNet_io_in_1_bits_payload_manager_xact_id = T_20455_bits_payload_manager_xact_id;
  assign gntNet_io_in_1_bits_payload_is_builtin_type = T_20455_bits_payload_is_builtin_type;
  assign gntNet_io_in_1_bits_payload_g_type = T_20455_bits_payload_g_type;
  assign gntNet_io_in_1_bits_payload_data = T_20455_bits_payload_data;
  assign gntNet_io_in_2_valid = 1'h0;
  assign gntNet_io_in_2_bits_header_src = GEN_47;
  assign gntNet_io_in_2_bits_header_dst = GEN_48;
  assign gntNet_io_in_2_bits_payload_addr_beat = GEN_49;
  assign gntNet_io_in_2_bits_payload_client_xact_id = GEN_50;
  assign gntNet_io_in_2_bits_payload_manager_xact_id = GEN_51;
  assign gntNet_io_in_2_bits_payload_is_builtin_type = GEN_52;
  assign gntNet_io_in_2_bits_payload_g_type = GEN_53;
  assign gntNet_io_in_2_bits_payload_data = GEN_54;
  assign gntNet_io_in_3_valid = 1'h0;
  assign gntNet_io_in_3_bits_header_src = GEN_55;
  assign gntNet_io_in_3_bits_header_dst = GEN_56;
  assign gntNet_io_in_3_bits_payload_addr_beat = GEN_57;
  assign gntNet_io_in_3_bits_payload_client_xact_id = GEN_58;
  assign gntNet_io_in_3_bits_payload_manager_xact_id = GEN_59;
  assign gntNet_io_in_3_bits_payload_is_builtin_type = GEN_60;
  assign gntNet_io_in_3_bits_payload_g_type = GEN_61;
  assign gntNet_io_in_3_bits_payload_data = GEN_62;
  assign gntNet_io_in_4_valid = 1'h0;
  assign gntNet_io_in_4_bits_header_src = GEN_63;
  assign gntNet_io_in_4_bits_header_dst = GEN_64;
  assign gntNet_io_in_4_bits_payload_addr_beat = GEN_65;
  assign gntNet_io_in_4_bits_payload_client_xact_id = GEN_66;
  assign gntNet_io_in_4_bits_payload_manager_xact_id = GEN_67;
  assign gntNet_io_in_4_bits_payload_is_builtin_type = GEN_68;
  assign gntNet_io_in_4_bits_payload_g_type = GEN_69;
  assign gntNet_io_in_4_bits_payload_data = GEN_70;
  assign gntNet_io_out_0_ready = 1'h0;
  assign gntNet_io_out_1_ready = 1'h0;
  assign gntNet_io_out_2_ready = T_20911_ready;
  assign gntNet_io_out_3_ready = T_21551_ready;
  assign gntNet_io_out_4_ready = T_22191_ready;
  assign ackNet_clk = clk;
  assign ackNet_reset = reset;
  assign ackNet_io_in_0_valid = 1'h0;
  assign ackNet_io_in_0_bits_header_src = GEN_71;
  assign ackNet_io_in_0_bits_header_dst = GEN_72;
  assign ackNet_io_in_0_bits_payload_manager_xact_id = GEN_73;
  assign ackNet_io_in_1_valid = 1'h0;
  assign ackNet_io_in_1_bits_header_src = GEN_74;
  assign ackNet_io_in_1_bits_header_dst = GEN_75;
  assign ackNet_io_in_1_bits_payload_manager_xact_id = GEN_76;
  assign ackNet_io_in_2_valid = T_23770_valid;
  assign ackNet_io_in_2_bits_header_src = T_23770_bits_header_src;
  assign ackNet_io_in_2_bits_header_dst = T_23770_bits_header_dst;
  assign ackNet_io_in_2_bits_payload_manager_xact_id = T_23770_bits_payload_manager_xact_id;
  assign ackNet_io_in_3_valid = T_23925_valid;
  assign ackNet_io_in_3_bits_header_src = T_23925_bits_header_src;
  assign ackNet_io_in_3_bits_header_dst = T_23925_bits_header_dst;
  assign ackNet_io_in_3_bits_payload_manager_xact_id = T_23925_bits_payload_manager_xact_id;
  assign ackNet_io_in_4_valid = T_24080_valid;
  assign ackNet_io_in_4_bits_header_src = T_24080_bits_header_src;
  assign ackNet_io_in_4_bits_header_dst = T_24080_bits_header_dst;
  assign ackNet_io_in_4_bits_payload_manager_xact_id = T_24080_bits_payload_manager_xact_id;
  assign ackNet_io_out_0_ready = T_22816_ready;
  assign ackNet_io_out_1_ready = T_23431_ready;
  assign ackNet_io_out_2_ready = 1'h0;
  assign ackNet_io_out_3_ready = 1'h0;
  assign ackNet_io_out_4_ready = 1'h0;
  assign T_14709_ready = TileLinkEnqueuer_17_14134_io_client_acquire_ready;
  assign T_14709_valid = acqNet_io_out_0_valid;
  assign T_14709_bits_header_src = T_14968;
  assign T_14709_bits_header_dst = acqNet_io_out_0_bits_header_dst;
  assign T_14709_bits_payload_addr_block = acqNet_io_out_0_bits_payload_addr_block;
  assign T_14709_bits_payload_client_xact_id = acqNet_io_out_0_bits_payload_client_xact_id;
  assign T_14709_bits_payload_addr_beat = acqNet_io_out_0_bits_payload_addr_beat;
  assign T_14709_bits_payload_is_builtin_type = acqNet_io_out_0_bits_payload_is_builtin_type;
  assign T_14709_bits_payload_a_type = acqNet_io_out_0_bits_payload_a_type;
  assign T_14709_bits_payload_union = acqNet_io_out_0_bits_payload_union;
  assign T_14709_bits_payload_data = acqNet_io_out_0_bits_payload_data;
  assign GEN_0 = {{1'd0}, 2'h2};
  assign T_14967 = acqNet_io_out_0_bits_header_src - GEN_0;
  assign T_14968 = T_14967[2:0];
  assign T_15354_ready = TileLinkEnqueuer_19_14136_io_client_acquire_ready;
  assign T_15354_valid = acqNet_io_out_1_valid;
  assign T_15354_bits_header_src = T_15613;
  assign T_15354_bits_header_dst = acqNet_io_out_1_bits_header_dst;
  assign T_15354_bits_payload_addr_block = acqNet_io_out_1_bits_payload_addr_block;
  assign T_15354_bits_payload_client_xact_id = acqNet_io_out_1_bits_payload_client_xact_id;
  assign T_15354_bits_payload_addr_beat = acqNet_io_out_1_bits_payload_addr_beat;
  assign T_15354_bits_payload_is_builtin_type = acqNet_io_out_1_bits_payload_is_builtin_type;
  assign T_15354_bits_payload_a_type = acqNet_io_out_1_bits_payload_a_type;
  assign T_15354_bits_payload_union = acqNet_io_out_1_bits_payload_union;
  assign T_15354_bits_payload_data = acqNet_io_out_1_bits_payload_data;
  assign T_15612 = acqNet_io_out_1_bits_header_src - GEN_0;
  assign T_15613 = T_15612[2:0];
  assign T_15723_ready = acqNet_io_in_2_ready;
  assign T_15723_valid = TileLinkEnqueuer_14127_io_manager_acquire_valid;
  assign T_15723_bits_header_src = T_15798;
  assign T_15723_bits_header_dst = TileLinkEnqueuer_14127_io_manager_acquire_bits_header_dst;
  assign T_15723_bits_payload_addr_block = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_block;
  assign T_15723_bits_payload_client_xact_id = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_client_xact_id;
  assign T_15723_bits_payload_addr_beat = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_addr_beat;
  assign T_15723_bits_payload_is_builtin_type = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_15723_bits_payload_a_type = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_a_type;
  assign T_15723_bits_payload_union = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_union;
  assign T_15723_bits_payload_data = TileLinkEnqueuer_14127_io_manager_acquire_bits_payload_data;
  assign T_15797 = TileLinkEnqueuer_14127_io_manager_acquire_bits_header_src + 3'h2;
  assign T_15798 = T_15797[2:0];
  assign T_15908_ready = acqNet_io_in_3_ready;
  assign T_15908_valid = TileLinkEnqueuer_4_14129_io_manager_acquire_valid;
  assign T_15908_bits_header_src = T_15983;
  assign T_15908_bits_header_dst = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_dst;
  assign T_15908_bits_payload_addr_block = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_block;
  assign T_15908_bits_payload_client_xact_id = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_client_xact_id;
  assign T_15908_bits_payload_addr_beat = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_addr_beat;
  assign T_15908_bits_payload_is_builtin_type = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_15908_bits_payload_a_type = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_a_type;
  assign T_15908_bits_payload_union = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_union;
  assign T_15908_bits_payload_data = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_payload_data;
  assign T_15982 = TileLinkEnqueuer_4_14129_io_manager_acquire_bits_header_src + 3'h2;
  assign T_15983 = T_15982[2:0];
  assign T_16093_ready = acqNet_io_in_4_ready;
  assign T_16093_valid = TileLinkEnqueuer_9_14131_io_manager_acquire_valid;
  assign T_16093_bits_header_src = T_16168;
  assign T_16093_bits_header_dst = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_dst;
  assign T_16093_bits_payload_addr_block = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_block;
  assign T_16093_bits_payload_client_xact_id = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_client_xact_id;
  assign T_16093_bits_payload_addr_beat = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_addr_beat;
  assign T_16093_bits_payload_is_builtin_type = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_is_builtin_type;
  assign T_16093_bits_payload_a_type = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_a_type;
  assign T_16093_bits_payload_union = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_union;
  assign T_16093_bits_payload_data = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_payload_data;
  assign T_16167 = TileLinkEnqueuer_9_14131_io_manager_acquire_bits_header_src + 3'h2;
  assign T_16168 = T_16167[2:0];
  assign T_16551_ready = TileLinkEnqueuer_17_14134_io_client_release_ready;
  assign T_16551_valid = relNet_io_out_0_valid;
  assign T_16551_bits_header_src = T_16808;
  assign T_16551_bits_header_dst = relNet_io_out_0_bits_header_dst;
  assign T_16551_bits_payload_addr_beat = relNet_io_out_0_bits_payload_addr_beat;
  assign T_16551_bits_payload_addr_block = relNet_io_out_0_bits_payload_addr_block;
  assign T_16551_bits_payload_client_xact_id = relNet_io_out_0_bits_payload_client_xact_id;
  assign T_16551_bits_payload_voluntary = relNet_io_out_0_bits_payload_voluntary;
  assign T_16551_bits_payload_r_type = relNet_io_out_0_bits_payload_r_type;
  assign T_16551_bits_payload_data = relNet_io_out_0_bits_payload_data;
  assign T_16807 = relNet_io_out_0_bits_header_src - GEN_0;
  assign T_16808 = T_16807[2:0];
  assign T_17191_ready = TileLinkEnqueuer_19_14136_io_client_release_ready;
  assign T_17191_valid = relNet_io_out_1_valid;
  assign T_17191_bits_header_src = T_17448;
  assign T_17191_bits_header_dst = relNet_io_out_1_bits_header_dst;
  assign T_17191_bits_payload_addr_beat = relNet_io_out_1_bits_payload_addr_beat;
  assign T_17191_bits_payload_addr_block = relNet_io_out_1_bits_payload_addr_block;
  assign T_17191_bits_payload_client_xact_id = relNet_io_out_1_bits_payload_client_xact_id;
  assign T_17191_bits_payload_voluntary = relNet_io_out_1_bits_payload_voluntary;
  assign T_17191_bits_payload_r_type = relNet_io_out_1_bits_payload_r_type;
  assign T_17191_bits_payload_data = relNet_io_out_1_bits_payload_data;
  assign T_17447 = relNet_io_out_1_bits_header_src - GEN_0;
  assign T_17448 = T_17447[2:0];
  assign T_17555_ready = relNet_io_in_2_ready;
  assign T_17555_valid = TileLinkEnqueuer_14127_io_manager_release_valid;
  assign T_17555_bits_header_src = T_17628;
  assign T_17555_bits_header_dst = TileLinkEnqueuer_14127_io_manager_release_bits_header_dst;
  assign T_17555_bits_payload_addr_beat = TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_beat;
  assign T_17555_bits_payload_addr_block = TileLinkEnqueuer_14127_io_manager_release_bits_payload_addr_block;
  assign T_17555_bits_payload_client_xact_id = TileLinkEnqueuer_14127_io_manager_release_bits_payload_client_xact_id;
  assign T_17555_bits_payload_voluntary = TileLinkEnqueuer_14127_io_manager_release_bits_payload_voluntary;
  assign T_17555_bits_payload_r_type = TileLinkEnqueuer_14127_io_manager_release_bits_payload_r_type;
  assign T_17555_bits_payload_data = TileLinkEnqueuer_14127_io_manager_release_bits_payload_data;
  assign T_17627 = TileLinkEnqueuer_14127_io_manager_release_bits_header_src + 3'h2;
  assign T_17628 = T_17627[2:0];
  assign T_17735_ready = relNet_io_in_3_ready;
  assign T_17735_valid = TileLinkEnqueuer_4_14129_io_manager_release_valid;
  assign T_17735_bits_header_src = T_17808;
  assign T_17735_bits_header_dst = TileLinkEnqueuer_4_14129_io_manager_release_bits_header_dst;
  assign T_17735_bits_payload_addr_beat = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_beat;
  assign T_17735_bits_payload_addr_block = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_addr_block;
  assign T_17735_bits_payload_client_xact_id = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_client_xact_id;
  assign T_17735_bits_payload_voluntary = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_voluntary;
  assign T_17735_bits_payload_r_type = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_r_type;
  assign T_17735_bits_payload_data = TileLinkEnqueuer_4_14129_io_manager_release_bits_payload_data;
  assign T_17807 = TileLinkEnqueuer_4_14129_io_manager_release_bits_header_src + 3'h2;
  assign T_17808 = T_17807[2:0];
  assign T_17915_ready = relNet_io_in_4_ready;
  assign T_17915_valid = TileLinkEnqueuer_9_14131_io_manager_release_valid;
  assign T_17915_bits_header_src = T_17988;
  assign T_17915_bits_header_dst = TileLinkEnqueuer_9_14131_io_manager_release_bits_header_dst;
  assign T_17915_bits_payload_addr_beat = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_beat;
  assign T_17915_bits_payload_addr_block = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_addr_block;
  assign T_17915_bits_payload_client_xact_id = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_client_xact_id;
  assign T_17915_bits_payload_voluntary = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_voluntary;
  assign T_17915_bits_payload_r_type = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_r_type;
  assign T_17915_bits_payload_data = TileLinkEnqueuer_9_14131_io_manager_release_bits_payload_data;
  assign T_17987 = TileLinkEnqueuer_9_14131_io_manager_release_bits_header_src + 3'h2;
  assign T_17988 = T_17987[2:0];
  assign T_18083_ready = prbNet_io_in_0_ready;
  assign T_18083_valid = TileLinkEnqueuer_17_14134_io_client_probe_valid;
  assign T_18083_bits_header_src = TileLinkEnqueuer_17_14134_io_client_probe_bits_header_src;
  assign T_18083_bits_header_dst = T_18148;
  assign T_18083_bits_payload_addr_block = TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_addr_block;
  assign T_18083_bits_payload_p_type = TileLinkEnqueuer_17_14134_io_client_probe_bits_payload_p_type;
  assign T_18147 = TileLinkEnqueuer_17_14134_io_client_probe_bits_header_dst + 3'h2;
  assign T_18148 = T_18147[2:0];
  assign T_18243_ready = prbNet_io_in_1_ready;
  assign T_18243_valid = TileLinkEnqueuer_19_14136_io_client_probe_valid;
  assign T_18243_bits_header_src = TileLinkEnqueuer_19_14136_io_client_probe_bits_header_src;
  assign T_18243_bits_header_dst = T_18308;
  assign T_18243_bits_payload_addr_block = TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_addr_block;
  assign T_18243_bits_payload_p_type = TileLinkEnqueuer_19_14136_io_client_probe_bits_payload_p_type;
  assign T_18307 = TileLinkEnqueuer_19_14136_io_client_probe_bits_header_dst + 3'h2;
  assign T_18308 = T_18307[2:0];
  assign T_18679_ready = TileLinkEnqueuer_14127_io_manager_probe_ready;
  assign T_18679_valid = prbNet_io_out_2_valid;
  assign T_18679_bits_header_src = prbNet_io_out_2_bits_header_src;
  assign T_18679_bits_header_dst = T_18928;
  assign T_18679_bits_payload_addr_block = prbNet_io_out_2_bits_payload_addr_block;
  assign T_18679_bits_payload_p_type = prbNet_io_out_2_bits_payload_p_type;
  assign T_18927 = prbNet_io_out_2_bits_header_dst - GEN_0;
  assign T_18928 = T_18927[2:0];
  assign T_19299_ready = TileLinkEnqueuer_4_14129_io_manager_probe_ready;
  assign T_19299_valid = prbNet_io_out_3_valid;
  assign T_19299_bits_header_src = prbNet_io_out_3_bits_header_src;
  assign T_19299_bits_header_dst = T_19548;
  assign T_19299_bits_payload_addr_block = prbNet_io_out_3_bits_payload_addr_block;
  assign T_19299_bits_payload_p_type = prbNet_io_out_3_bits_payload_p_type;
  assign T_19547 = prbNet_io_out_3_bits_header_dst - GEN_0;
  assign T_19548 = T_19547[2:0];
  assign T_19919_ready = TileLinkEnqueuer_9_14131_io_manager_probe_ready;
  assign T_19919_valid = prbNet_io_out_4_valid;
  assign T_19919_bits_header_src = prbNet_io_out_4_bits_header_src;
  assign T_19919_bits_header_dst = T_20168;
  assign T_19919_bits_payload_addr_block = prbNet_io_out_4_bits_payload_addr_block;
  assign T_19919_bits_payload_p_type = prbNet_io_out_4_bits_payload_p_type;
  assign T_20167 = prbNet_io_out_4_bits_header_dst - GEN_0;
  assign T_20168 = T_20167[2:0];
  assign T_20275_ready = gntNet_io_in_0_ready;
  assign T_20275_valid = TileLinkEnqueuer_17_14134_io_client_grant_valid;
  assign T_20275_bits_header_src = TileLinkEnqueuer_17_14134_io_client_grant_bits_header_src;
  assign T_20275_bits_header_dst = T_20348;
  assign T_20275_bits_payload_addr_beat = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_addr_beat;
  assign T_20275_bits_payload_client_xact_id = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_client_xact_id;
  assign T_20275_bits_payload_manager_xact_id = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_manager_xact_id;
  assign T_20275_bits_payload_is_builtin_type = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_is_builtin_type;
  assign T_20275_bits_payload_g_type = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_g_type;
  assign T_20275_bits_payload_data = TileLinkEnqueuer_17_14134_io_client_grant_bits_payload_data;
  assign T_20347 = TileLinkEnqueuer_17_14134_io_client_grant_bits_header_dst + 3'h2;
  assign T_20348 = T_20347[2:0];
  assign T_20455_ready = gntNet_io_in_1_ready;
  assign T_20455_valid = TileLinkEnqueuer_19_14136_io_client_grant_valid;
  assign T_20455_bits_header_src = TileLinkEnqueuer_19_14136_io_client_grant_bits_header_src;
  assign T_20455_bits_header_dst = T_20528;
  assign T_20455_bits_payload_addr_beat = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_addr_beat;
  assign T_20455_bits_payload_client_xact_id = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_client_xact_id;
  assign T_20455_bits_payload_manager_xact_id = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_manager_xact_id;
  assign T_20455_bits_payload_is_builtin_type = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_is_builtin_type;
  assign T_20455_bits_payload_g_type = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_g_type;
  assign T_20455_bits_payload_data = TileLinkEnqueuer_19_14136_io_client_grant_bits_payload_data;
  assign T_20527 = TileLinkEnqueuer_19_14136_io_client_grant_bits_header_dst + 3'h2;
  assign T_20528 = T_20527[2:0];
  assign T_20911_ready = TileLinkEnqueuer_14127_io_manager_grant_ready;
  assign T_20911_valid = gntNet_io_out_2_valid;
  assign T_20911_bits_header_src = gntNet_io_out_2_bits_header_src;
  assign T_20911_bits_header_dst = T_21168;
  assign T_20911_bits_payload_addr_beat = gntNet_io_out_2_bits_payload_addr_beat;
  assign T_20911_bits_payload_client_xact_id = gntNet_io_out_2_bits_payload_client_xact_id;
  assign T_20911_bits_payload_manager_xact_id = gntNet_io_out_2_bits_payload_manager_xact_id;
  assign T_20911_bits_payload_is_builtin_type = gntNet_io_out_2_bits_payload_is_builtin_type;
  assign T_20911_bits_payload_g_type = gntNet_io_out_2_bits_payload_g_type;
  assign T_20911_bits_payload_data = gntNet_io_out_2_bits_payload_data;
  assign T_21167 = gntNet_io_out_2_bits_header_dst - GEN_0;
  assign T_21168 = T_21167[2:0];
  assign T_21551_ready = TileLinkEnqueuer_4_14129_io_manager_grant_ready;
  assign T_21551_valid = gntNet_io_out_3_valid;
  assign T_21551_bits_header_src = gntNet_io_out_3_bits_header_src;
  assign T_21551_bits_header_dst = T_21808;
  assign T_21551_bits_payload_addr_beat = gntNet_io_out_3_bits_payload_addr_beat;
  assign T_21551_bits_payload_client_xact_id = gntNet_io_out_3_bits_payload_client_xact_id;
  assign T_21551_bits_payload_manager_xact_id = gntNet_io_out_3_bits_payload_manager_xact_id;
  assign T_21551_bits_payload_is_builtin_type = gntNet_io_out_3_bits_payload_is_builtin_type;
  assign T_21551_bits_payload_g_type = gntNet_io_out_3_bits_payload_g_type;
  assign T_21551_bits_payload_data = gntNet_io_out_3_bits_payload_data;
  assign T_21807 = gntNet_io_out_3_bits_header_dst - GEN_0;
  assign T_21808 = T_21807[2:0];
  assign T_22191_ready = TileLinkEnqueuer_9_14131_io_manager_grant_ready;
  assign T_22191_valid = gntNet_io_out_4_valid;
  assign T_22191_bits_header_src = gntNet_io_out_4_bits_header_src;
  assign T_22191_bits_header_dst = T_22448;
  assign T_22191_bits_payload_addr_beat = gntNet_io_out_4_bits_payload_addr_beat;
  assign T_22191_bits_payload_client_xact_id = gntNet_io_out_4_bits_payload_client_xact_id;
  assign T_22191_bits_payload_manager_xact_id = gntNet_io_out_4_bits_payload_manager_xact_id;
  assign T_22191_bits_payload_is_builtin_type = gntNet_io_out_4_bits_payload_is_builtin_type;
  assign T_22191_bits_payload_g_type = gntNet_io_out_4_bits_payload_g_type;
  assign T_22191_bits_payload_data = gntNet_io_out_4_bits_payload_data;
  assign T_22447 = gntNet_io_out_4_bits_header_dst - GEN_0;
  assign T_22448 = T_22447[2:0];
  assign T_22816_ready = TileLinkEnqueuer_17_14134_io_client_finish_ready;
  assign T_22816_valid = ackNet_io_out_0_valid;
  assign T_22816_bits_header_src = T_23063;
  assign T_22816_bits_header_dst = ackNet_io_out_0_bits_header_dst;
  assign T_22816_bits_payload_manager_xact_id = ackNet_io_out_0_bits_payload_manager_xact_id;
  assign T_23062 = ackNet_io_out_0_bits_header_src - GEN_0;
  assign T_23063 = T_23062[2:0];
  assign T_23431_ready = TileLinkEnqueuer_19_14136_io_client_finish_ready;
  assign T_23431_valid = ackNet_io_out_1_valid;
  assign T_23431_bits_header_src = T_23678;
  assign T_23431_bits_header_dst = ackNet_io_out_1_bits_header_dst;
  assign T_23431_bits_payload_manager_xact_id = ackNet_io_out_1_bits_payload_manager_xact_id;
  assign T_23677 = ackNet_io_out_1_bits_header_src - GEN_0;
  assign T_23678 = T_23677[2:0];
  assign T_23770_ready = ackNet_io_in_2_ready;
  assign T_23770_valid = TileLinkEnqueuer_14127_io_manager_finish_valid;
  assign T_23770_bits_header_src = T_23833;
  assign T_23770_bits_header_dst = TileLinkEnqueuer_14127_io_manager_finish_bits_header_dst;
  assign T_23770_bits_payload_manager_xact_id = TileLinkEnqueuer_14127_io_manager_finish_bits_payload_manager_xact_id;
  assign T_23832 = TileLinkEnqueuer_14127_io_manager_finish_bits_header_src + 3'h2;
  assign T_23833 = T_23832[2:0];
  assign T_23925_ready = ackNet_io_in_3_ready;
  assign T_23925_valid = TileLinkEnqueuer_4_14129_io_manager_finish_valid;
  assign T_23925_bits_header_src = T_23988;
  assign T_23925_bits_header_dst = TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_dst;
  assign T_23925_bits_payload_manager_xact_id = TileLinkEnqueuer_4_14129_io_manager_finish_bits_payload_manager_xact_id;
  assign T_23987 = TileLinkEnqueuer_4_14129_io_manager_finish_bits_header_src + 3'h2;
  assign T_23988 = T_23987[2:0];
  assign T_24080_ready = ackNet_io_in_4_ready;
  assign T_24080_valid = TileLinkEnqueuer_9_14131_io_manager_finish_valid;
  assign T_24080_bits_header_src = T_24143;
  assign T_24080_bits_header_dst = TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_dst;
  assign T_24080_bits_payload_manager_xact_id = TileLinkEnqueuer_9_14131_io_manager_finish_bits_payload_manager_xact_id;
  assign T_24142 = TileLinkEnqueuer_9_14131_io_manager_finish_bits_header_src + 3'h2;
  assign T_24143 = T_24142[2:0];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_77 = {1{$random}};
  GEN_1 = GEN_77[2:0];
  GEN_78 = {1{$random}};
  GEN_2 = GEN_78[2:0];
  GEN_79 = {1{$random}};
  GEN_3 = GEN_79[25:0];
  GEN_80 = {1{$random}};
  GEN_4 = GEN_80[1:0];
  GEN_81 = {1{$random}};
  GEN_5 = GEN_81[2:0];
  GEN_82 = {1{$random}};
  GEN_6 = GEN_82[0:0];
  GEN_83 = {1{$random}};
  GEN_7 = GEN_83[2:0];
  GEN_84 = {1{$random}};
  GEN_8 = GEN_84[11:0];
  GEN_85 = {2{$random}};
  GEN_9 = GEN_85[63:0];
  GEN_86 = {1{$random}};
  GEN_10 = GEN_86[2:0];
  GEN_87 = {1{$random}};
  GEN_11 = GEN_87[2:0];
  GEN_88 = {1{$random}};
  GEN_12 = GEN_88[25:0];
  GEN_89 = {1{$random}};
  GEN_13 = GEN_89[1:0];
  GEN_90 = {1{$random}};
  GEN_14 = GEN_90[2:0];
  GEN_91 = {1{$random}};
  GEN_15 = GEN_91[0:0];
  GEN_92 = {1{$random}};
  GEN_16 = GEN_92[2:0];
  GEN_93 = {1{$random}};
  GEN_17 = GEN_93[11:0];
  GEN_94 = {2{$random}};
  GEN_18 = GEN_94[63:0];
  GEN_95 = {1{$random}};
  GEN_19 = GEN_95[2:0];
  GEN_96 = {1{$random}};
  GEN_20 = GEN_96[2:0];
  GEN_97 = {1{$random}};
  GEN_21 = GEN_97[2:0];
  GEN_98 = {1{$random}};
  GEN_22 = GEN_98[25:0];
  GEN_99 = {1{$random}};
  GEN_23 = GEN_99[1:0];
  GEN_100 = {1{$random}};
  GEN_24 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  GEN_25 = GEN_101[2:0];
  GEN_102 = {2{$random}};
  GEN_26 = GEN_102[63:0];
  GEN_103 = {1{$random}};
  GEN_27 = GEN_103[2:0];
  GEN_104 = {1{$random}};
  GEN_28 = GEN_104[2:0];
  GEN_105 = {1{$random}};
  GEN_29 = GEN_105[2:0];
  GEN_106 = {1{$random}};
  GEN_30 = GEN_106[25:0];
  GEN_107 = {1{$random}};
  GEN_31 = GEN_107[1:0];
  GEN_108 = {1{$random}};
  GEN_32 = GEN_108[0:0];
  GEN_109 = {1{$random}};
  GEN_33 = GEN_109[2:0];
  GEN_110 = {2{$random}};
  GEN_34 = GEN_110[63:0];
  GEN_111 = {1{$random}};
  GEN_35 = GEN_111[2:0];
  GEN_112 = {1{$random}};
  GEN_36 = GEN_112[2:0];
  GEN_113 = {1{$random}};
  GEN_37 = GEN_113[25:0];
  GEN_114 = {1{$random}};
  GEN_38 = GEN_114[1:0];
  GEN_115 = {1{$random}};
  GEN_39 = GEN_115[2:0];
  GEN_116 = {1{$random}};
  GEN_40 = GEN_116[2:0];
  GEN_117 = {1{$random}};
  GEN_41 = GEN_117[25:0];
  GEN_118 = {1{$random}};
  GEN_42 = GEN_118[1:0];
  GEN_119 = {1{$random}};
  GEN_43 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  GEN_44 = GEN_120[2:0];
  GEN_121 = {1{$random}};
  GEN_45 = GEN_121[25:0];
  GEN_122 = {1{$random}};
  GEN_46 = GEN_122[1:0];
  GEN_123 = {1{$random}};
  GEN_47 = GEN_123[2:0];
  GEN_124 = {1{$random}};
  GEN_48 = GEN_124[2:0];
  GEN_125 = {1{$random}};
  GEN_49 = GEN_125[2:0];
  GEN_126 = {1{$random}};
  GEN_50 = GEN_126[1:0];
  GEN_127 = {1{$random}};
  GEN_51 = GEN_127[2:0];
  GEN_128 = {1{$random}};
  GEN_52 = GEN_128[0:0];
  GEN_129 = {1{$random}};
  GEN_53 = GEN_129[3:0];
  GEN_130 = {2{$random}};
  GEN_54 = GEN_130[63:0];
  GEN_131 = {1{$random}};
  GEN_55 = GEN_131[2:0];
  GEN_132 = {1{$random}};
  GEN_56 = GEN_132[2:0];
  GEN_133 = {1{$random}};
  GEN_57 = GEN_133[2:0];
  GEN_134 = {1{$random}};
  GEN_58 = GEN_134[1:0];
  GEN_135 = {1{$random}};
  GEN_59 = GEN_135[2:0];
  GEN_136 = {1{$random}};
  GEN_60 = GEN_136[0:0];
  GEN_137 = {1{$random}};
  GEN_61 = GEN_137[3:0];
  GEN_138 = {2{$random}};
  GEN_62 = GEN_138[63:0];
  GEN_139 = {1{$random}};
  GEN_63 = GEN_139[2:0];
  GEN_140 = {1{$random}};
  GEN_64 = GEN_140[2:0];
  GEN_141 = {1{$random}};
  GEN_65 = GEN_141[2:0];
  GEN_142 = {1{$random}};
  GEN_66 = GEN_142[1:0];
  GEN_143 = {1{$random}};
  GEN_67 = GEN_143[2:0];
  GEN_144 = {1{$random}};
  GEN_68 = GEN_144[0:0];
  GEN_145 = {1{$random}};
  GEN_69 = GEN_145[3:0];
  GEN_146 = {2{$random}};
  GEN_70 = GEN_146[63:0];
  GEN_147 = {1{$random}};
  GEN_71 = GEN_147[2:0];
  GEN_148 = {1{$random}};
  GEN_72 = GEN_148[2:0];
  GEN_149 = {1{$random}};
  GEN_73 = GEN_149[2:0];
  GEN_150 = {1{$random}};
  GEN_74 = GEN_150[2:0];
  GEN_151 = {1{$random}};
  GEN_75 = GEN_151[2:0];
  GEN_152 = {1{$random}};
  GEN_76 = GEN_152[2:0];
  end
`endif
endmodule
module BroadcastVoluntaryReleaseTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [4:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [4:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [4:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [4:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [4:0] io_outer_grant_bits_data,
  output  io_matches_iacq,
  output  io_matches_irel,
  output  io_matches_oprb,
  input   io_alloc_iacq,
  input   io_alloc_irel,
  input   io_alloc_oprb
);
  reg  state;
  reg [31:0] GEN_29;
  reg [2:0] xact_addr_beat;
  reg [31:0] GEN_38;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_39;
  reg [1:0] xact_client_xact_id;
  reg [31:0] GEN_40;
  reg  xact_voluntary;
  reg [31:0] GEN_41;
  reg [2:0] xact_r_type;
  reg [31:0] GEN_42;
  reg [4:0] xact_data_buffer_0;
  reg [31:0] GEN_43;
  reg [4:0] xact_data_buffer_1;
  reg [31:0] GEN_45;
  reg [4:0] xact_data_buffer_2;
  reg [31:0] GEN_46;
  reg [4:0] xact_data_buffer_3;
  reg [31:0] GEN_47;
  reg [4:0] xact_data_buffer_4;
  reg [31:0] GEN_53;
  reg [4:0] xact_data_buffer_5;
  reg [31:0] GEN_56;
  reg [4:0] xact_data_buffer_6;
  reg [31:0] GEN_62;
  reg [4:0] xact_data_buffer_7;
  reg [31:0] GEN_64;
  reg [7:0] xact_wmask_buffer_0;
  reg [31:0] GEN_65;
  reg [7:0] xact_wmask_buffer_1;
  reg [31:0] GEN_67;
  reg [7:0] xact_wmask_buffer_2;
  reg [31:0] GEN_68;
  reg [7:0] xact_wmask_buffer_3;
  reg [31:0] GEN_69;
  reg [7:0] xact_wmask_buffer_4;
  reg [31:0] GEN_70;
  reg [7:0] xact_wmask_buffer_5;
  reg [31:0] GEN_72;
  reg [7:0] xact_wmask_buffer_6;
  reg [31:0] GEN_74;
  reg [7:0] xact_wmask_buffer_7;
  reg [31:0] GEN_75;
  reg [1:0] xact_client_id;
  reg [31:0] GEN_76;
  wire  coh_sharers;
  reg [7:0] pending_irels;
  reg [31:0] GEN_77;
  reg [7:0] pending_writes;
  reg [31:0] GEN_78;
  reg  pending_ignt;
  reg [31:0] GEN_79;
  wire [7:0] GEN_52;
  wire  T_286;
  wire  T_288;
  wire  T_289;
  wire  T_290;
  wire  all_pending_done;
  wire  T_292;
  wire [2:0] T_298_0;
  wire [2:0] T_298_1;
  wire [2:0] T_298_2;
  wire  T_300;
  wire  T_301;
  wire  T_302;
  wire  T_305;
  wire  T_306;
  wire  T_307;
  wire [7:0] GEN_54;
  wire [8:0] T_309;
  wire [7:0] T_310;
  wire [7:0] T_311;
  wire [7:0] GEN_55;
  wire [7:0] T_313;
  wire [7:0] T_314;
  wire [7:0] T_315;
  wire [7:0] T_316;
  wire  T_317;
  wire  T_318;
  wire  T_321;
  wire [4:0] GEN_0;
  wire [2:0] GEN_57;
  wire [4:0] GEN_2;
  wire [2:0] GEN_58;
  wire [4:0] GEN_3;
  wire [2:0] GEN_59;
  wire [4:0] GEN_4;
  wire [2:0] GEN_60;
  wire [4:0] GEN_5;
  wire [4:0] GEN_6;
  wire [4:0] GEN_7;
  wire [4:0] GEN_8;
  wire [4:0] GEN_9;
  wire [4:0] GEN_11;
  wire [4:0] GEN_12;
  wire [4:0] GEN_13;
  wire [4:0] GEN_14;
  wire [4:0] GEN_15;
  wire [4:0] GEN_16;
  wire [4:0] GEN_17;
  wire [4:0] GEN_18;
  wire  T_323;
  wire [2:0] T_332_0;
  wire [2:0] T_332_1;
  wire [2:0] T_332_2;
  wire  T_334;
  wire  T_335;
  wire  T_336;
  wire  T_339;
  wire  T_340;
  wire  T_341;
  wire  T_342;
  wire [7:0] GEN_61;
  wire [8:0] T_344;
  wire [7:0] T_345;
  wire [7:0] T_346;
  wire [7:0] T_348;
  wire [7:0] T_349;
  wire [7:0] T_350;
  wire [7:0] T_351;
  wire [2:0] T_359_0;
  wire [2:0] T_359_1;
  wire [2:0] T_359_2;
  wire  T_361;
  wire  T_362;
  wire  T_363;
  wire  T_366;
  wire  T_367;
  wire  T_368;
  wire [7:0] GEN_63;
  wire [8:0] T_371;
  wire [7:0] T_372;
  wire [7:0] T_375;
  wire [7:0] T_376;
  wire  T_377;
  wire  T_378;
  wire  T_379;
  wire  T_380;
  wire  T_381;
  wire  T_382;
  wire  T_383;
  wire [2:0] T_393;
  wire [2:0] T_394;
  wire [2:0] T_395;
  wire [2:0] T_396;
  wire [2:0] T_397;
  wire [2:0] T_398;
  wire [2:0] curr_write_beat;
  wire  T_402;
  wire [7:0] GEN_66;
  wire [7:0] T_407;
  wire [8:0] T_432;
  wire [11:0] T_450;
  wire [25:0] T_465_addr_block;
  wire [1:0] T_465_client_xact_id;
  wire [2:0] T_465_addr_beat;
  wire  T_465_is_builtin_type;
  wire [2:0] T_465_a_type;
  wire [11:0] T_465_union;
  wire [4:0] T_465_data;
  wire [4:0] GEN_1;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [4:0] GEN_25;
  wire  T_474;
  wire  T_476;
  wire  T_477;
  wire  T_478;
  wire [2:0] T_492_addr_beat;
  wire [1:0] T_492_client_xact_id;
  wire [2:0] T_492_manager_xact_id;
  wire  T_492_is_builtin_type;
  wire [3:0] T_492_g_type;
  wire [4:0] T_492_data;
  wire [1:0] T_492_client_id;
  wire  T_500;
  wire  GEN_26;
  wire  T_503;
  wire  T_505;
  wire  T_506;
  wire [2:0] T_513_0;
  wire [2:0] T_513_1;
  wire [2:0] T_513_2;
  wire  T_515;
  wire  T_516;
  wire  T_517;
  wire  T_520;
  wire  T_521;
  wire [2:0] T_529_0;
  wire [2:0] T_529_1;
  wire [2:0] T_529_2;
  wire  T_531;
  wire  T_532;
  wire  T_533;
  wire  T_536;
  wire  T_537;
  wire  T_538;
  wire [7:0] GEN_71;
  wire [8:0] T_540;
  wire [7:0] T_541;
  wire [7:0] T_542;
  wire [7:0] T_546;
  wire [7:0] GEN_30;
  wire  T_548;
  wire [7:0] GEN_31;
  wire [2:0] T_557_0;
  wire [2:0] T_557_1;
  wire [2:0] T_557_2;
  wire  T_559;
  wire  T_560;
  wire  T_561;
  wire  T_564;
  wire  T_565;
  wire  T_566;
  wire [7:0] GEN_73;
  wire [8:0] T_569;
  wire [7:0] T_570;
  wire [7:0] T_573;
  wire [2:0] GEN_32;
  wire [25:0] GEN_33;
  wire [1:0] GEN_34;
  wire  GEN_35;
  wire [2:0] GEN_36;
  wire [1:0] GEN_37;
  wire [7:0] GEN_44;
  wire [7:0] GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  T_578;
  wire  GEN_51;
  wire  T_580;
  wire  T_581;
  wire  T_583;
  wire  T_584;
  wire  T_585;
  wire  T_589;
  wire  T_591;
  wire  T_592;
  wire  T_594;
  wire  T_595;
  wire  T_597;
  reg [25:0] GEN_10;
  reg [31:0] GEN_80;
  reg [1:0] GEN_27;
  reg [31:0] GEN_81;
  reg [1:0] GEN_28;
  reg [31:0] GEN_82;
  assign io_inner_acquire_ready = 1'h0;
  assign io_inner_grant_valid = T_478;
  assign io_inner_grant_bits_addr_beat = T_492_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_492_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_492_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_492_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_492_g_type;
  assign io_inner_grant_bits_data = T_492_data;
  assign io_inner_grant_bits_client_id = T_492_client_id;
  assign io_inner_finish_ready = 1'h0;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_10;
  assign io_inner_probe_bits_p_type = GEN_27;
  assign io_inner_probe_bits_client_id = GEN_28;
  assign io_inner_release_ready = T_321;
  assign io_outer_acquire_valid = T_402;
  assign io_outer_acquire_bits_addr_block = T_465_addr_block;
  assign io_outer_acquire_bits_client_xact_id = {{1'd0}, T_465_client_xact_id};
  assign io_outer_acquire_bits_addr_beat = T_465_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_465_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_465_a_type;
  assign io_outer_acquire_bits_union = T_465_union;
  assign io_outer_acquire_bits_data = T_465_data;
  assign io_outer_grant_ready = T_503;
  assign io_matches_iacq = T_581;
  assign io_matches_irel = T_585;
  assign io_matches_oprb = 1'h0;
  assign coh_sharers = 1'h0;
  assign GEN_52 = {{7'd0}, 1'h0};
  assign T_286 = pending_irels != GEN_52;
  assign T_288 = pending_writes != GEN_52;
  assign T_289 = T_286 | T_288;
  assign T_290 = T_289 | pending_ignt;
  assign all_pending_done = T_290 == 1'h0;
  assign T_292 = io_inner_release_ready & io_inner_release_valid;
  assign T_298_0 = 3'h0;
  assign T_298_1 = 3'h1;
  assign T_298_2 = 3'h2;
  assign T_300 = T_298_0 == io_inner_release_bits_r_type;
  assign T_301 = T_298_1 == io_inner_release_bits_r_type;
  assign T_302 = T_298_2 == io_inner_release_bits_r_type;
  assign T_305 = T_300 | T_301;
  assign T_306 = T_305 | T_302;
  assign T_307 = T_292 & T_306;
  assign GEN_54 = {{7'd0}, T_307};
  assign T_309 = 8'h0 - GEN_54;
  assign T_310 = T_309[7:0];
  assign T_311 = ~ T_310;
  assign GEN_55 = {{7'd0}, 1'h1};
  assign T_313 = GEN_55 << io_inner_release_bits_addr_beat;
  assign T_314 = ~ T_313;
  assign T_315 = T_311 | T_314;
  assign T_316 = pending_irels & T_315;
  assign T_317 = state == 1'h0;
  assign T_318 = T_317 & io_inner_release_bits_voluntary;
  assign T_321 = T_318 | T_286;
  assign GEN_0 = io_inner_release_bits_data;
  assign GEN_57 = {{2'd0}, 1'h0};
  assign GEN_2 = GEN_57 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_0;
  assign GEN_58 = {{2'd0}, 1'h1};
  assign GEN_3 = GEN_58 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_1;
  assign GEN_59 = {{1'd0}, 2'h2};
  assign GEN_4 = GEN_59 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_2;
  assign GEN_60 = {{1'd0}, 2'h3};
  assign GEN_5 = GEN_60 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_3;
  assign GEN_6 = 3'h4 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_4;
  assign GEN_7 = 3'h5 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_5;
  assign GEN_8 = 3'h6 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_6;
  assign GEN_9 = 3'h7 == io_inner_release_bits_addr_beat ? GEN_0 : xact_data_buffer_7;
  assign GEN_11 = T_292 ? GEN_2 : xact_data_buffer_0;
  assign GEN_12 = T_292 ? GEN_3 : xact_data_buffer_1;
  assign GEN_13 = T_292 ? GEN_4 : xact_data_buffer_2;
  assign GEN_14 = T_292 ? GEN_5 : xact_data_buffer_3;
  assign GEN_15 = T_292 ? GEN_6 : xact_data_buffer_4;
  assign GEN_16 = T_292 ? GEN_7 : xact_data_buffer_5;
  assign GEN_17 = T_292 ? GEN_8 : xact_data_buffer_6;
  assign GEN_18 = T_292 ? GEN_9 : xact_data_buffer_7;
  assign T_323 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_332_0 = 3'h2;
  assign T_332_1 = 3'h3;
  assign T_332_2 = 3'h4;
  assign T_334 = T_332_0 == io_outer_acquire_bits_a_type;
  assign T_335 = T_332_1 == io_outer_acquire_bits_a_type;
  assign T_336 = T_332_2 == io_outer_acquire_bits_a_type;
  assign T_339 = T_334 | T_335;
  assign T_340 = T_339 | T_336;
  assign T_341 = io_outer_acquire_bits_is_builtin_type & T_340;
  assign T_342 = T_323 & T_341;
  assign GEN_61 = {{7'd0}, T_342};
  assign T_344 = 8'h0 - GEN_61;
  assign T_345 = T_344[7:0];
  assign T_346 = ~ T_345;
  assign T_348 = GEN_55 << io_outer_acquire_bits_addr_beat;
  assign T_349 = ~ T_348;
  assign T_350 = T_346 | T_349;
  assign T_351 = pending_writes & T_350;
  assign T_359_0 = 3'h0;
  assign T_359_1 = 3'h1;
  assign T_359_2 = 3'h2;
  assign T_361 = T_359_0 == io_inner_release_bits_r_type;
  assign T_362 = T_359_1 == io_inner_release_bits_r_type;
  assign T_363 = T_359_2 == io_inner_release_bits_r_type;
  assign T_366 = T_361 | T_362;
  assign T_367 = T_366 | T_363;
  assign T_368 = T_292 & T_367;
  assign GEN_63 = {{7'd0}, T_368};
  assign T_371 = 8'h0 - GEN_63;
  assign T_372 = T_371[7:0];
  assign T_375 = T_372 & T_313;
  assign T_376 = T_351 | T_375;
  assign T_377 = pending_writes[0];
  assign T_378 = pending_writes[1];
  assign T_379 = pending_writes[2];
  assign T_380 = pending_writes[3];
  assign T_381 = pending_writes[4];
  assign T_382 = pending_writes[5];
  assign T_383 = pending_writes[6];
  assign T_393 = T_383 ? 3'h6 : 3'h7;
  assign T_394 = T_382 ? 3'h5 : T_393;
  assign T_395 = T_381 ? 3'h4 : T_394;
  assign T_396 = T_380 ? {{1'd0}, 2'h3} : T_395;
  assign T_397 = T_379 ? {{1'd0}, 2'h2} : T_396;
  assign T_398 = T_378 ? {{2'd0}, 1'h1} : T_397;
  assign curr_write_beat = T_377 ? {{2'd0}, 1'h0} : T_398;
  assign T_402 = state & T_288;
  assign GEN_66 = $signed(8'hff);
  assign T_407 = $unsigned(GEN_66);
  assign T_432 = {T_407,1'h1};
  assign T_450 = 1'h1 ? {{3'd0}, T_432} : 12'h0;
  assign T_465_addr_block = xact_addr_block;
  assign T_465_client_xact_id = {{1'd0}, 1'h0};
  assign T_465_addr_beat = curr_write_beat;
  assign T_465_is_builtin_type = 1'h1;
  assign T_465_a_type = 3'h3;
  assign T_465_union = T_450;
  assign T_465_data = GEN_1;
  assign GEN_1 = GEN_25;
  assign GEN_19 = GEN_58 == curr_write_beat ? xact_data_buffer_1 : xact_data_buffer_0;
  assign GEN_20 = GEN_59 == curr_write_beat ? xact_data_buffer_2 : GEN_19;
  assign GEN_21 = GEN_60 == curr_write_beat ? xact_data_buffer_3 : GEN_20;
  assign GEN_22 = 3'h4 == curr_write_beat ? xact_data_buffer_4 : GEN_21;
  assign GEN_23 = 3'h5 == curr_write_beat ? xact_data_buffer_5 : GEN_22;
  assign GEN_24 = 3'h6 == curr_write_beat ? xact_data_buffer_6 : GEN_23;
  assign GEN_25 = 3'h7 == curr_write_beat ? xact_data_buffer_7 : GEN_24;
  assign T_474 = state & pending_ignt;
  assign T_476 = pending_irels == GEN_52;
  assign T_477 = T_474 & T_476;
  assign T_478 = T_477 & io_outer_grant_valid;
  assign T_492_addr_beat = {{2'd0}, 1'h0};
  assign T_492_client_xact_id = xact_client_xact_id;
  assign T_492_manager_xact_id = {{2'd0}, 1'h0};
  assign T_492_is_builtin_type = 1'h1;
  assign T_492_g_type = {{1'd0}, 3'h0};
  assign T_492_data = {{4'd0}, 1'h0};
  assign T_492_client_id = xact_client_id;
  assign T_500 = io_inner_grant_ready & io_inner_grant_valid;
  assign GEN_26 = T_500 ? 1'h0 : pending_ignt;
  assign T_503 = state & io_inner_grant_ready;
  assign T_505 = T_317 & io_inner_release_valid;
  assign T_506 = T_505 & io_alloc_irel;
  assign T_513_0 = 3'h0;
  assign T_513_1 = 3'h1;
  assign T_513_2 = 3'h2;
  assign T_515 = T_513_0 == io_inner_release_bits_r_type;
  assign T_516 = T_513_1 == io_inner_release_bits_r_type;
  assign T_517 = T_513_2 == io_inner_release_bits_r_type;
  assign T_520 = T_515 | T_516;
  assign T_521 = T_520 | T_517;
  assign T_529_0 = 3'h0;
  assign T_529_1 = 3'h1;
  assign T_529_2 = 3'h2;
  assign T_531 = T_529_0 == io_inner_release_bits_r_type;
  assign T_532 = T_529_1 == io_inner_release_bits_r_type;
  assign T_533 = T_529_2 == io_inner_release_bits_r_type;
  assign T_536 = T_531 | T_532;
  assign T_537 = T_536 | T_533;
  assign T_538 = T_292 & T_537;
  assign GEN_71 = {{7'd0}, T_538};
  assign T_540 = 8'h0 - GEN_71;
  assign T_541 = T_540[7:0];
  assign T_542 = ~ T_541;
  assign T_546 = T_542 | T_314;
  assign GEN_30 = T_521 ? T_546 : T_316;
  assign T_548 = T_521 == 1'h0;
  assign GEN_31 = T_548 ? {{7'd0}, 1'h0} : GEN_30;
  assign T_557_0 = 3'h0;
  assign T_557_1 = 3'h1;
  assign T_557_2 = 3'h2;
  assign T_559 = T_557_0 == io_inner_release_bits_r_type;
  assign T_560 = T_557_1 == io_inner_release_bits_r_type;
  assign T_561 = T_557_2 == io_inner_release_bits_r_type;
  assign T_564 = T_559 | T_560;
  assign T_565 = T_564 | T_561;
  assign T_566 = T_292 & T_565;
  assign GEN_73 = {{7'd0}, T_566};
  assign T_569 = 8'h0 - GEN_73;
  assign T_570 = T_569[7:0];
  assign T_573 = T_570 & T_313;
  assign GEN_32 = T_506 ? io_inner_release_bits_addr_beat : xact_addr_beat;
  assign GEN_33 = T_506 ? io_inner_release_bits_addr_block : xact_addr_block;
  assign GEN_34 = T_506 ? io_inner_release_bits_client_xact_id : xact_client_xact_id;
  assign GEN_35 = T_506 ? io_inner_release_bits_voluntary : xact_voluntary;
  assign GEN_36 = T_506 ? io_inner_release_bits_r_type : xact_r_type;
  assign GEN_37 = T_506 ? io_inner_release_bits_client_id : xact_client_id;
  assign GEN_44 = T_506 ? GEN_31 : T_316;
  assign GEN_48 = T_506 ? T_573 : T_376;
  assign GEN_49 = T_506 ? 1'h1 : GEN_26;
  assign GEN_50 = T_506 ? 1'h1 : state;
  assign T_578 = state & all_pending_done;
  assign GEN_51 = T_578 ? 1'h0 : GEN_50;
  assign T_580 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign T_581 = state & T_580;
  assign T_583 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T_584 = state & T_583;
  assign T_585 = T_584 & io_inner_release_bits_voluntary;
  assign T_589 = T_317 & T_292;
  assign T_591 = io_inner_release_bits_voluntary == 1'h0;
  assign T_592 = T_589 & T_591;
  assign T_594 = T_592 == 1'h0;
  assign T_595 = T_594 | reset;
  assign T_597 = T_595 == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_29 = {1{$random}};
  state = GEN_29[0:0];
  GEN_38 = {1{$random}};
  xact_addr_beat = GEN_38[2:0];
  GEN_39 = {1{$random}};
  xact_addr_block = GEN_39[25:0];
  GEN_40 = {1{$random}};
  xact_client_xact_id = GEN_40[1:0];
  GEN_41 = {1{$random}};
  xact_voluntary = GEN_41[0:0];
  GEN_42 = {1{$random}};
  xact_r_type = GEN_42[2:0];
  GEN_43 = {1{$random}};
  xact_data_buffer_0 = GEN_43[4:0];
  GEN_45 = {1{$random}};
  xact_data_buffer_1 = GEN_45[4:0];
  GEN_46 = {1{$random}};
  xact_data_buffer_2 = GEN_46[4:0];
  GEN_47 = {1{$random}};
  xact_data_buffer_3 = GEN_47[4:0];
  GEN_53 = {1{$random}};
  xact_data_buffer_4 = GEN_53[4:0];
  GEN_56 = {1{$random}};
  xact_data_buffer_5 = GEN_56[4:0];
  GEN_62 = {1{$random}};
  xact_data_buffer_6 = GEN_62[4:0];
  GEN_64 = {1{$random}};
  xact_data_buffer_7 = GEN_64[4:0];
  GEN_65 = {1{$random}};
  xact_wmask_buffer_0 = GEN_65[7:0];
  GEN_67 = {1{$random}};
  xact_wmask_buffer_1 = GEN_67[7:0];
  GEN_68 = {1{$random}};
  xact_wmask_buffer_2 = GEN_68[7:0];
  GEN_69 = {1{$random}};
  xact_wmask_buffer_3 = GEN_69[7:0];
  GEN_70 = {1{$random}};
  xact_wmask_buffer_4 = GEN_70[7:0];
  GEN_72 = {1{$random}};
  xact_wmask_buffer_5 = GEN_72[7:0];
  GEN_74 = {1{$random}};
  xact_wmask_buffer_6 = GEN_74[7:0];
  GEN_75 = {1{$random}};
  xact_wmask_buffer_7 = GEN_75[7:0];
  GEN_76 = {1{$random}};
  xact_client_id = GEN_76[1:0];
  GEN_77 = {1{$random}};
  pending_irels = GEN_77[7:0];
  GEN_78 = {1{$random}};
  pending_writes = GEN_78[7:0];
  GEN_79 = {1{$random}};
  pending_ignt = GEN_79[0:0];
  GEN_80 = {1{$random}};
  GEN_10 = GEN_80[25:0];
  GEN_81 = {1{$random}};
  GEN_27 = GEN_81[1:0];
  GEN_82 = {1{$random}};
  GEN_28 = GEN_82[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 1'h0;
    end else begin
      state <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      xact_addr_beat <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      xact_addr_block <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      xact_client_xact_id <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      xact_voluntary <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      xact_r_type <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_0 <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_1 <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_2 <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_3 <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_4 <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_5 <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_6 <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_7 <= GEN_18;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      xact_client_id <= GEN_37;
    end
    if(reset) begin
      pending_irels <= 8'h0;
    end else begin
      pending_irels <= GEN_44;
    end
    if(reset) begin
      pending_writes <= 8'h0;
    end else begin
      pending_writes <= GEN_48;
    end
    if(reset) begin
      pending_ignt <= 1'h0;
    end else begin
      pending_ignt <= GEN_49;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_597) begin
          $fwrite(32'h80000002,"Assertion failed: VoluntaryReleaseTracker accepted Release that wasn't voluntary!\n    at broadcast.scala:191 assert(!(state === s_idle && io.inner.release.fire() && !io.irel().isVoluntary()),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_597) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module BroadcastAcquireTracker(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [4:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [4:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [4:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [4:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [4:0] io_outer_grant_bits_data,
  output  io_matches_iacq,
  output  io_matches_irel,
  output  io_matches_oprb,
  input   io_alloc_iacq,
  input   io_alloc_irel,
  input   io_alloc_oprb
);
  reg [2:0] state;
  reg [31:0] GEN_41;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_50;
  reg [1:0] xact_client_xact_id;
  reg [31:0] GEN_51;
  reg [2:0] xact_addr_beat;
  reg [31:0] GEN_62;
  reg  xact_is_builtin_type;
  reg [31:0] GEN_63;
  reg [2:0] xact_a_type;
  reg [31:0] GEN_72;
  reg [11:0] xact_union;
  reg [31:0] GEN_73;
  reg [4:0] xact_data_buffer_0;
  reg [31:0] GEN_85;
  reg [4:0] xact_data_buffer_1;
  reg [31:0] GEN_87;
  reg [4:0] xact_data_buffer_2;
  reg [31:0] GEN_88;
  reg [4:0] xact_data_buffer_3;
  reg [31:0] GEN_89;
  reg [4:0] xact_data_buffer_4;
  reg [31:0] GEN_90;
  reg [4:0] xact_data_buffer_5;
  reg [31:0] GEN_91;
  reg [4:0] xact_data_buffer_6;
  reg [31:0] GEN_92;
  reg [4:0] xact_data_buffer_7;
  reg [31:0] GEN_93;
  reg [7:0] xact_wmask_buffer_0;
  reg [31:0] GEN_94;
  reg [7:0] xact_wmask_buffer_1;
  reg [31:0] GEN_95;
  reg [7:0] xact_wmask_buffer_2;
  reg [31:0] GEN_96;
  reg [7:0] xact_wmask_buffer_3;
  reg [31:0] GEN_97;
  reg [7:0] xact_wmask_buffer_4;
  reg [31:0] GEN_98;
  reg [7:0] xact_wmask_buffer_5;
  reg [31:0] GEN_99;
  reg [7:0] xact_wmask_buffer_6;
  reg [31:0] GEN_100;
  reg [7:0] xact_wmask_buffer_7;
  reg [31:0] GEN_101;
  reg [1:0] xact_client_id;
  reg [31:0] GEN_102;
  wire  coh_sharers;
  wire  T_284;
  wire  T_285;
  wire [2:0] T_294_0;
  wire [2:0] T_294_1;
  wire [2:0] T_294_2;
  wire  T_296;
  wire  T_297;
  wire  T_298;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_305;
  wire  T_306;
  wire  T_308;
  reg  release_count;
  reg [31:0] GEN_112;
  reg  pending_probes;
  reg [31:0] GEN_114;
  wire  GEN_229;
  wire  T_313;
  wire [3:0] GEN_230;
  wire [3:0] T_316;
  wire  T_318;
  wire [3:0] GEN_232;
  wire [3:0] T_319;
  wire [3:0] T_320;
  wire  T_321;
  wire [3:0] GEN_233;
  wire [3:0] mask_incoherent;
  reg  collect_iacq_data;
  reg [31:0] GEN_115;
  reg [7:0] iacq_data_valid;
  reg [31:0] GEN_116;
  wire  T_324;
  wire [2:0] T_334_0;
  wire  T_336;
  wire  T_339;
  wire  T_340;
  reg [2:0] T_342;
  reg [31:0] GEN_117;
  wire  T_344;
  wire [2:0] GEN_234;
  wire [3:0] T_346;
  wire [2:0] T_347;
  wire [2:0] GEN_6;
  wire  T_348;
  wire  iacq_data_done;
  wire  T_350;
  wire [2:0] T_358_0;
  wire [2:0] T_358_1;
  wire [2:0] T_358_2;
  wire  T_360;
  wire  T_361;
  wire  T_362;
  wire  T_365;
  wire  T_366;
  wire  T_368;
  reg [2:0] T_370;
  reg [31:0] GEN_118;
  wire [3:0] T_374;
  wire [2:0] T_375;
  wire [2:0] GEN_7;
  wire  T_379;
  wire [2:0] T_387_0;
  wire [3:0] GEN_236;
  wire  T_389;
  wire [1:0] T_397_0;
  wire [1:0] T_397_1;
  wire [3:0] GEN_237;
  wire  T_399;
  wire [3:0] GEN_238;
  wire  T_400;
  wire  T_403;
  wire  T_404;
  wire  T_406;
  reg [2:0] T_408;
  reg [31:0] GEN_119;
  wire  T_410;
  wire [3:0] T_412;
  wire [2:0] T_413;
  wire [2:0] GEN_8;
  wire  T_414;
  wire  ignt_data_done;
  wire  T_416;
  wire [2:0] T_425_0;
  wire  T_427;
  wire  T_430;
  wire  T_431;
  reg [2:0] T_433;
  reg [31:0] GEN_120;
  wire  T_435;
  wire [3:0] T_437;
  wire [2:0] T_438;
  wire [2:0] GEN_9;
  wire  T_439;
  wire [2:0] oacq_data_cnt;
  wire  oacq_data_done;
  wire  T_440;
  wire [2:0] T_449_0;
  wire [3:0] GEN_241;
  wire  T_451;
  wire  T_459_0;
  wire [3:0] GEN_242;
  wire  T_461;
  wire  T_464;
  wire  T_466;
  reg [2:0] T_468;
  reg [31:0] GEN_121;
  wire [3:0] T_472;
  wire [2:0] T_473;
  wire [2:0] GEN_10;
  reg  pending_ognt_ack;
  reg [31:0] GEN_122;
  wire [2:0] T_485_0;
  wire [2:0] T_485_1;
  wire [2:0] T_485_2;
  wire  T_487;
  wire  T_488;
  wire  T_489;
  wire  T_492;
  wire  T_493;
  wire  pending_outer_write;
  wire [2:0] T_502_0;
  wire [2:0] T_502_1;
  wire [2:0] T_502_2;
  wire  T_504;
  wire  T_505;
  wire  T_506;
  wire  T_509;
  wire  T_510;
  wire  pending_outer_write_;
  wire [2:0] T_518_0;
  wire [2:0] T_518_1;
  wire [3:0] GEN_244;
  wire  T_520;
  wire [3:0] GEN_245;
  wire  T_521;
  wire  T_524;
  wire [1:0] T_530_0;
  wire [1:0] T_530_1;
  wire [3:0] GEN_246;
  wire  T_532;
  wire [3:0] GEN_247;
  wire  T_533;
  wire  T_536;
  wire  pending_outer_read;
  wire  T_555;
  wire [2:0] T_556;
  wire  T_557;
  wire [2:0] T_558;
  wire  T_559;
  wire [2:0] T_560;
  wire  T_561;
  wire [2:0] T_562;
  wire  T_563;
  wire [2:0] T_564;
  wire  T_565;
  wire [2:0] T_566;
  wire  T_567;
  wire [2:0] T_568;
  wire [2:0] GEN_248;
  wire  T_569;
  wire [1:0] T_574;
  wire [2:0] T_575;
  wire [2:0] T_584_addr_beat;
  wire [1:0] T_584_client_xact_id;
  wire [2:0] T_584_manager_xact_id;
  wire  T_584_is_builtin_type;
  wire [3:0] T_584_g_type;
  wire [4:0] T_584_data;
  wire [1:0] T_584_client_id;
  wire [2:0] T_599_0;
  wire [2:0] T_599_1;
  wire [3:0] GEN_249;
  wire  T_601;
  wire [3:0] GEN_250;
  wire  T_602;
  wire  T_605;
  wire [1:0] T_611_0;
  wire [1:0] T_611_1;
  wire [3:0] GEN_251;
  wire  T_613;
  wire [3:0] GEN_252;
  wire  T_614;
  wire  T_617;
  wire  pending_outer_read_;
  wire [2:0] T_626_0;
  wire [2:0] T_626_1;
  wire [2:0] T_626_2;
  wire  T_628;
  wire  T_629;
  wire  T_630;
  wire  T_633;
  wire  T_634;
  wire  subblock_type;
  wire  T_636;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire  T_642;
  wire  T_643;
  wire [7:0] GEN_253;
  wire [7:0] T_649;
  wire [8:0] T_674;
  wire [11:0] T_692;
  wire [25:0] oacq_probe_addr_block;
  wire [2:0] oacq_probe_client_xact_id;
  wire [2:0] oacq_probe_addr_beat;
  wire  oacq_probe_is_builtin_type;
  wire [2:0] oacq_probe_a_type;
  wire [11:0] oacq_probe_union;
  wire [4:0] oacq_probe_data;
  wire  T_716;
  wire  T_717;
  wire [7:0] GEN_254;
  wire [8:0] T_721;
  wire [7:0] T_722;
  wire [7:0] T_728_0;
  wire  T_731;
  wire  T_732;
  wire  T_734;
  wire  T_735;
  wire  T_736;
  wire [7:0] T_737;
  wire [7:0] T_739;
  wire [7:0] T_740;
  wire [8:0] T_767;
  wire [11:0] T_787;
  wire [25:0] oacq_write_beat_addr_block;
  wire [2:0] oacq_write_beat_client_xact_id;
  wire [2:0] oacq_write_beat_addr_beat;
  wire  oacq_write_beat_is_builtin_type;
  wire [2:0] oacq_write_beat_a_type;
  wire [11:0] oacq_write_beat_union;
  wire [4:0] oacq_write_beat_data;
  wire [7:0] GEN_0;
  wire [7:0] GEN_11;
  wire [2:0] GEN_256;
  wire [7:0] GEN_12;
  wire [2:0] GEN_257;
  wire [7:0] GEN_13;
  wire [7:0] GEN_14;
  wire [7:0] GEN_15;
  wire [7:0] GEN_16;
  wire [7:0] GEN_17;
  wire [8:0] T_834;
  wire [11:0] T_852;
  wire [25:0] oacq_write_block_addr_block;
  wire [2:0] oacq_write_block_client_xact_id;
  wire [2:0] oacq_write_block_addr_beat;
  wire  oacq_write_block_is_builtin_type;
  wire [2:0] oacq_write_block_a_type;
  wire [11:0] oacq_write_block_union;
  wire [4:0] oacq_write_block_data;
  wire [4:0] GEN_1;
  wire [4:0] GEN_18;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [2:0] T_875;
  wire [2:0] T_876;
  wire [5:0] T_897;
  wire [11:0] T_898;
  wire [25:0] oacq_read_beat_addr_block;
  wire [2:0] oacq_read_beat_client_xact_id;
  wire [2:0] oacq_read_beat_addr_beat;
  wire  oacq_read_beat_is_builtin_type;
  wire [2:0] oacq_read_beat_a_type;
  wire [11:0] oacq_read_beat_union;
  wire [4:0] oacq_read_beat_data;
  wire [25:0] oacq_read_block_addr_block;
  wire [2:0] oacq_read_block_client_xact_id;
  wire [2:0] oacq_read_block_addr_beat;
  wire  oacq_read_block_is_builtin_type;
  wire [2:0] oacq_read_block_a_type;
  wire [11:0] oacq_read_block_union;
  wire [4:0] oacq_read_block_data;
  wire  T_1013;
  wire  T_1014;
  wire [25:0] T_1015_addr_block;
  wire [2:0] T_1015_client_xact_id;
  wire [2:0] T_1015_addr_beat;
  wire  T_1015_is_builtin_type;
  wire [2:0] T_1015_a_type;
  wire [11:0] T_1015_union;
  wire [4:0] T_1015_data;
  wire [25:0] T_1023_addr_block;
  wire [2:0] T_1023_client_xact_id;
  wire [2:0] T_1023_addr_beat;
  wire  T_1023_is_builtin_type;
  wire [2:0] T_1023_a_type;
  wire [11:0] T_1023_union;
  wire [4:0] T_1023_data;
  wire [25:0] T_1031_addr_block;
  wire [2:0] T_1031_client_xact_id;
  wire [2:0] T_1031_addr_beat;
  wire  T_1031_is_builtin_type;
  wire [2:0] T_1031_a_type;
  wire [11:0] T_1031_union;
  wire [4:0] T_1031_data;
  wire [25:0] T_1039_addr_block;
  wire [2:0] T_1039_client_xact_id;
  wire [2:0] T_1039_addr_beat;
  wire  T_1039_is_builtin_type;
  wire [2:0] T_1039_a_type;
  wire [11:0] T_1039_union;
  wire [4:0] T_1039_data;
  wire  T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire  T_1060;
  wire [1:0] T_1061;
  wire  T_1062;
  wire [1:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire  T_1066;
  wire [1:0] T_1067;
  wire  T_1068;
  wire [1:0] T_1069;
  wire  T_1070;
  wire [1:0] T_1071;
  wire  T_1072;
  wire [1:0] T_1073;
  wire [1:0] T_1074;
  wire [25:0] T_1079_addr_block;
  wire [1:0] T_1079_p_type;
  wire [1:0] T_1079_client_id;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1107;
  wire [2:0] T_1109;
  wire [2:0] T_1111;
  wire [2:0] T_1113;
  wire [2:0] T_1115;
  wire  T_1116;
  wire [1:0] T_1121;
  wire [2:0] T_1122;
  wire [2:0] T_1131_addr_beat;
  wire [1:0] T_1131_client_xact_id;
  wire [2:0] T_1131_manager_xact_id;
  wire  T_1131_is_builtin_type;
  wire [3:0] T_1131_g_type;
  wire [4:0] T_1131_data;
  wire [1:0] T_1131_client_id;
  wire  T_1143;
  wire  T_1145;
  wire  T_1146;
  wire  T_1147;
  wire  T_1149;
  wire  T_1150;
  wire  T_1152;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire [2:0] T_1176_0;
  wire  T_1178;
  wire  T_1181;
  wire  T_1182;
  wire  T_1184;
  wire  T_1185;
  wire  T_1187;
  wire  T_1188;
  wire  T_1190;
  wire [4:0] GEN_2;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire [4:0] GEN_29;
  wire [4:0] GEN_30;
  wire [4:0] GEN_31;
  wire [4:0] GEN_32;
  wire  T_1193;
  wire  T_1194;
  wire [7:0] T_1205_0;
  wire  T_1208;
  wire  T_1209;
  wire  T_1211;
  wire  T_1212;
  wire  T_1213;
  wire [7:0] T_1214;
  wire [7:0] T_1216;
  wire [7:0] T_1217;
  wire [7:0] GEN_3;
  wire [7:0] GEN_33;
  wire [7:0] GEN_34;
  wire [7:0] GEN_35;
  wire [7:0] GEN_36;
  wire [7:0] GEN_37;
  wire [7:0] GEN_38;
  wire [7:0] GEN_39;
  wire [7:0] GEN_40;
  wire [7:0] T_1220;
  wire [7:0] T_1221;
  wire [4:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [4:0] GEN_45;
  wire [4:0] GEN_46;
  wire [4:0] GEN_47;
  wire [4:0] GEN_48;
  wire [4:0] GEN_49;
  wire [7:0] GEN_52;
  wire [7:0] GEN_53;
  wire [7:0] GEN_54;
  wire [7:0] GEN_55;
  wire [7:0] GEN_56;
  wire [7:0] GEN_57;
  wire [7:0] GEN_58;
  wire [7:0] GEN_59;
  wire [7:0] GEN_60;
  wire  GEN_61;
  wire [4:0] GEN_64;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] GEN_71;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire [7:0] GEN_78;
  wire [7:0] GEN_79;
  wire [7:0] GEN_80;
  wire [7:0] GEN_81;
  wire [7:0] GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_86;
  wire  T_1229;
  wire  T_1231;
  wire [4:0] GEN_4;
  wire [7:0] T_1247_0;
  wire [7:0] T_1259;
  wire [7:0] GEN_5;
  wire [2:0] T_1268_0;
  wire  T_1270;
  wire  T_1273;
  wire [2:0] T_1282_0;
  wire [2:0] T_1282_1;
  wire [2:0] T_1282_2;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1289;
  wire  T_1290;
  wire  T_1291;
  wire [7:0] GEN_276;
  wire [7:0] T_1292;
  wire [3:0] GEN_277;
  wire  T_1294;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire  T_1298;
  wire [1:0] T_1300;
  wire [1:0] GEN_278;
  wire [2:0] T_1301;
  wire [1:0] T_1302;
  wire [1:0] T_1305;
  wire [1:0] GEN_279;
  wire [2:0] T_1306;
  wire [1:0] T_1307;
  wire [2:0] T_1308;
  wire [2:0] GEN_280;
  wire [3:0] T_1309;
  wire [2:0] T_1310;
  wire [3:0] GEN_103;
  wire [2:0] GEN_104;
  wire [2:0] T_1311;
  wire [2:0] T_1312;
  wire [2:0] T_1313;
  wire [25:0] GEN_105;
  wire [1:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire [2:0] GEN_109;
  wire [11:0] GEN_110;
  wire [1:0] GEN_111;
  wire [4:0] GEN_113;
  wire [7:0] GEN_123;
  wire  GEN_132;
  wire [7:0] GEN_136;
  wire [3:0] GEN_137;
  wire [2:0] GEN_138;
  wire [2:0] GEN_139;
  wire  GEN_140;
  wire [25:0] GEN_141;
  wire [1:0] GEN_142;
  wire [2:0] GEN_143;
  wire  GEN_144;
  wire [2:0] GEN_145;
  wire [11:0] GEN_146;
  wire [1:0] GEN_147;
  wire [4:0] GEN_149;
  wire [7:0] GEN_159;
  wire  GEN_168;
  wire [7:0] GEN_172;
  wire [3:0] GEN_173;
  wire [2:0] GEN_174;
  wire [2:0] GEN_175;
  wire  T_1314;
  wire [1:0] GEN_281;
  wire [1:0] T_1318;
  wire [1:0] T_1319;
  wire [1:0] GEN_282;
  wire [1:0] T_1320;
  wire [3:0] GEN_176;
  wire [2:0] T_1326_0;
  wire [2:0] T_1326_1;
  wire [2:0] T_1326_2;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire  T_1339;
  wire [2:0] T_1345_0;
  wire [2:0] T_1345_1;
  wire [2:0] T_1345_2;
  wire  T_1347;
  wire  T_1348;
  wire  T_1349;
  wire  T_1352;
  wire  T_1353;
  wire [1:0] T_1357;
  wire  T_1358;
  wire [2:0] T_1361;
  wire [2:0] T_1362;
  wire [2:0] GEN_177;
  wire  GEN_178;
  wire [2:0] GEN_179;
  wire [2:0] GEN_180;
  wire  GEN_181;
  wire [2:0] GEN_182;
  wire [2:0] GEN_183;
  wire  GEN_185;
  wire [2:0] GEN_186;
  wire [2:0] GEN_187;
  wire  T_1364;
  wire [2:0] GEN_188;
  wire [2:0] GEN_189;
  wire [2:0] GEN_190;
  wire  GEN_194;
  wire  GEN_195;
  wire [2:0] GEN_196;
  wire [2:0] GEN_197;
  wire  GEN_198;
  wire [3:0] GEN_199;
  wire  GEN_203;
  wire  GEN_207;
  wire  GEN_208;
  wire [2:0] GEN_209;
  wire [2:0] GEN_210;
  wire  T_1372;
  wire  T_1374;
  wire  T_1376;
  wire [7:0] T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1380;
  wire [2:0] T_1382;
  wire  GEN_211;
  wire [2:0] GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire [2:0] GEN_215;
  wire  T_1383;
  wire [2:0] GEN_216;
  wire  GEN_217;
  wire [2:0] GEN_218;
  wire  T_1387;
  wire [3:0] GEN_283;
  wire  T_1392;
  wire  T_1393;
  wire  T_1395;
  wire [2:0] T_1397;
  wire [2:0] GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire [2:0] GEN_222;
  wire  T_1398;
  wire [2:0] GEN_223;
  wire  GEN_224;
  wire [2:0] GEN_225;
  wire  T_1410;
  wire [2:0] GEN_226;
  wire [2:0] GEN_228;
  assign io_inner_acquire_ready = GEN_140;
  assign io_inner_grant_valid = GEN_224;
  assign io_inner_grant_bits_addr_beat = T_1131_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1131_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1131_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1131_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1131_g_type;
  assign io_inner_grant_bits_data = T_1131_data;
  assign io_inner_grant_bits_client_id = T_1131_client_id;
  assign io_inner_finish_ready = T_1410;
  assign io_inner_probe_valid = GEN_198;
  assign io_inner_probe_bits_addr_block = T_1079_addr_block;
  assign io_inner_probe_bits_p_type = T_1079_p_type;
  assign io_inner_probe_bits_client_id = T_1079_client_id;
  assign io_inner_release_ready = GEN_203;
  assign io_outer_acquire_valid = GEN_217;
  assign io_outer_acquire_bits_addr_block = T_1039_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_1039_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_1039_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_1039_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_1039_a_type;
  assign io_outer_acquire_bits_union = T_1039_union;
  assign io_outer_acquire_bits_data = T_1039_data;
  assign io_outer_grant_ready = GEN_220;
  assign io_matches_iacq = T_637;
  assign io_matches_irel = T_643;
  assign io_matches_oprb = 1'h0;
  assign coh_sharers = 1'h0;
  assign T_284 = state != 3'h0;
  assign T_285 = T_284 & xact_is_builtin_type;
  assign T_294_0 = 3'h4;
  assign T_294_1 = 3'h5;
  assign T_294_2 = 3'h6;
  assign T_296 = T_294_0 == xact_a_type;
  assign T_297 = T_294_1 == xact_a_type;
  assign T_298 = T_294_2 == xact_a_type;
  assign T_301 = T_296 | T_297;
  assign T_302 = T_301 | T_298;
  assign T_303 = T_285 & T_302;
  assign T_305 = T_303 == 1'h0;
  assign T_306 = T_305 | reset;
  assign T_308 = T_306 == 1'h0;
  assign GEN_229 = $signed(1'h1);
  assign T_313 = $unsigned(GEN_229);
  assign GEN_230 = {{3'd0}, 1'h1};
  assign T_316 = GEN_230 << io_inner_acquire_bits_client_id;
  assign T_318 = ~ T_313;
  assign GEN_232 = {{3'd0}, T_318};
  assign T_319 = GEN_232 | T_316;
  assign T_320 = ~ T_319;
  assign T_321 = ~ io_incoherent_0;
  assign GEN_233 = {{3'd0}, T_321};
  assign mask_incoherent = T_320 & GEN_233;
  assign T_324 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_334_0 = 3'h3;
  assign T_336 = T_334_0 == io_inner_acquire_bits_a_type;
  assign T_339 = io_inner_acquire_bits_is_builtin_type & T_336;
  assign T_340 = T_324 & T_339;
  assign T_344 = T_342 == 3'h7;
  assign GEN_234 = {{2'd0}, 1'h1};
  assign T_346 = T_342 + GEN_234;
  assign T_347 = T_346[2:0];
  assign GEN_6 = T_340 ? T_347 : T_342;
  assign T_348 = T_340 & T_344;
  assign iacq_data_done = T_339 ? T_348 : T_324;
  assign T_350 = io_inner_release_ready & io_inner_release_valid;
  assign T_358_0 = 3'h0;
  assign T_358_1 = 3'h1;
  assign T_358_2 = 3'h2;
  assign T_360 = T_358_0 == io_inner_release_bits_r_type;
  assign T_361 = T_358_1 == io_inner_release_bits_r_type;
  assign T_362 = T_358_2 == io_inner_release_bits_r_type;
  assign T_365 = T_360 | T_361;
  assign T_366 = T_365 | T_362;
  assign T_368 = T_350 & T_366;
  assign T_374 = T_370 + GEN_234;
  assign T_375 = T_374[2:0];
  assign GEN_7 = T_368 ? T_375 : T_370;
  assign T_379 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_387_0 = 3'h5;
  assign GEN_236 = {{1'd0}, T_387_0};
  assign T_389 = GEN_236 == io_inner_grant_bits_g_type;
  assign T_397_0 = 2'h0;
  assign T_397_1 = 2'h1;
  assign GEN_237 = {{2'd0}, T_397_0};
  assign T_399 = GEN_237 == io_inner_grant_bits_g_type;
  assign GEN_238 = {{2'd0}, T_397_1};
  assign T_400 = GEN_238 == io_inner_grant_bits_g_type;
  assign T_403 = T_399 | T_400;
  assign T_404 = io_inner_grant_bits_is_builtin_type ? T_389 : T_403;
  assign T_406 = T_379 & T_404;
  assign T_410 = T_408 == 3'h7;
  assign T_412 = T_408 + GEN_234;
  assign T_413 = T_412[2:0];
  assign GEN_8 = T_406 ? T_413 : T_408;
  assign T_414 = T_406 & T_410;
  assign ignt_data_done = T_404 ? T_414 : T_379;
  assign T_416 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_425_0 = 3'h3;
  assign T_427 = T_425_0 == io_outer_acquire_bits_a_type;
  assign T_430 = io_outer_acquire_bits_is_builtin_type & T_427;
  assign T_431 = T_416 & T_430;
  assign T_435 = T_433 == 3'h7;
  assign T_437 = T_433 + GEN_234;
  assign T_438 = T_437[2:0];
  assign GEN_9 = T_431 ? T_438 : T_433;
  assign T_439 = T_431 & T_435;
  assign oacq_data_cnt = T_430 ? T_433 : {{2'd0}, 1'h0};
  assign oacq_data_done = T_430 ? T_439 : T_416;
  assign T_440 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_449_0 = 3'h5;
  assign GEN_241 = {{1'd0}, T_449_0};
  assign T_451 = GEN_241 == io_outer_grant_bits_g_type;
  assign T_459_0 = 1'h0;
  assign GEN_242 = {{3'd0}, T_459_0};
  assign T_461 = GEN_242 == io_outer_grant_bits_g_type;
  assign T_464 = io_outer_grant_bits_is_builtin_type ? T_451 : T_461;
  assign T_466 = T_440 & T_464;
  assign T_472 = T_468 + GEN_234;
  assign T_473 = T_472[2:0];
  assign GEN_10 = T_466 ? T_473 : T_468;
  assign T_485_0 = 3'h2;
  assign T_485_1 = 3'h3;
  assign T_485_2 = 3'h4;
  assign T_487 = T_485_0 == xact_a_type;
  assign T_488 = T_485_1 == xact_a_type;
  assign T_489 = T_485_2 == xact_a_type;
  assign T_492 = T_487 | T_488;
  assign T_493 = T_492 | T_489;
  assign pending_outer_write = xact_is_builtin_type & T_493;
  assign T_502_0 = 3'h2;
  assign T_502_1 = 3'h3;
  assign T_502_2 = 3'h4;
  assign T_504 = T_502_0 == io_inner_acquire_bits_a_type;
  assign T_505 = T_502_1 == io_inner_acquire_bits_a_type;
  assign T_506 = T_502_2 == io_inner_acquire_bits_a_type;
  assign T_509 = T_504 | T_505;
  assign T_510 = T_509 | T_506;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T_510;
  assign T_518_0 = 3'h5;
  assign T_518_1 = 3'h4;
  assign GEN_244 = {{1'd0}, T_518_0};
  assign T_520 = GEN_244 == io_inner_grant_bits_g_type;
  assign GEN_245 = {{1'd0}, T_518_1};
  assign T_521 = GEN_245 == io_inner_grant_bits_g_type;
  assign T_524 = T_520 | T_521;
  assign T_530_0 = 2'h0;
  assign T_530_1 = 2'h1;
  assign GEN_246 = {{2'd0}, T_530_0};
  assign T_532 = GEN_246 == io_inner_grant_bits_g_type;
  assign GEN_247 = {{2'd0}, T_530_1};
  assign T_533 = GEN_247 == io_inner_grant_bits_g_type;
  assign T_536 = T_532 | T_533;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T_524 : T_536;
  assign T_555 = 3'h6 == io_inner_acquire_bits_a_type;
  assign T_556 = T_555 ? 3'h1 : 3'h3;
  assign T_557 = 3'h5 == io_inner_acquire_bits_a_type;
  assign T_558 = T_557 ? 3'h1 : T_556;
  assign T_559 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T_560 = T_559 ? 3'h4 : T_558;
  assign T_561 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T_562 = T_561 ? 3'h3 : T_560;
  assign T_563 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T_564 = T_563 ? 3'h3 : T_562;
  assign T_565 = 3'h1 == io_inner_acquire_bits_a_type;
  assign T_566 = T_565 ? 3'h5 : T_564;
  assign T_567 = 3'h0 == io_inner_acquire_bits_a_type;
  assign T_568 = T_567 ? 3'h4 : T_566;
  assign GEN_248 = {{2'd0}, 1'h0};
  assign T_569 = io_inner_acquire_bits_a_type == GEN_248;
  assign T_574 = T_569 ? 2'h0 : 2'h1;
  assign T_575 = io_inner_acquire_bits_is_builtin_type ? T_568 : {{1'd0}, T_574};
  assign T_584_addr_beat = {{2'd0}, 1'h0};
  assign T_584_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign T_584_manager_xact_id = {{2'd0}, 1'h1};
  assign T_584_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign T_584_g_type = {{1'd0}, T_575};
  assign T_584_data = {{4'd0}, 1'h0};
  assign T_584_client_id = io_inner_acquire_bits_client_id;
  assign T_599_0 = 3'h5;
  assign T_599_1 = 3'h4;
  assign GEN_249 = {{1'd0}, T_599_0};
  assign T_601 = GEN_249 == T_584_g_type;
  assign GEN_250 = {{1'd0}, T_599_1};
  assign T_602 = GEN_250 == T_584_g_type;
  assign T_605 = T_601 | T_602;
  assign T_611_0 = 2'h0;
  assign T_611_1 = 2'h1;
  assign GEN_251 = {{2'd0}, T_611_0};
  assign T_613 = GEN_251 == T_584_g_type;
  assign GEN_252 = {{2'd0}, T_611_1};
  assign T_614 = GEN_252 == T_584_g_type;
  assign T_617 = T_613 | T_614;
  assign pending_outer_read_ = T_584_is_builtin_type ? T_605 : T_617;
  assign T_626_0 = 3'h2;
  assign T_626_1 = 3'h0;
  assign T_626_2 = 3'h4;
  assign T_628 = T_626_0 == xact_a_type;
  assign T_629 = T_626_1 == xact_a_type;
  assign T_630 = T_626_2 == xact_a_type;
  assign T_633 = T_628 | T_629;
  assign T_634 = T_633 | T_630;
  assign subblock_type = xact_is_builtin_type & T_634;
  assign T_636 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign T_637 = T_284 & T_636;
  assign T_639 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T_640 = T_284 & T_639;
  assign T_642 = io_inner_release_bits_voluntary == 1'h0;
  assign T_643 = T_640 & T_642;
  assign GEN_253 = $signed(8'hff);
  assign T_649 = $unsigned(GEN_253);
  assign T_674 = {T_649,1'h1};
  assign T_692 = 1'h1 ? {{3'd0}, T_674} : 12'h0;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign oacq_probe_client_xact_id = {{2'd0}, 1'h1};
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign oacq_probe_a_type = 3'h3;
  assign oacq_probe_union = T_692;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T_716 = xact_a_type == 3'h4;
  assign T_717 = xact_is_builtin_type & T_716;
  assign GEN_254 = {{7'd0}, 1'h1};
  assign T_721 = 8'h0 - GEN_254;
  assign T_722 = T_721[7:0];
  assign T_728_0 = T_722;
  assign T_731 = xact_a_type == 3'h3;
  assign T_732 = xact_is_builtin_type & T_731;
  assign T_734 = xact_a_type == 3'h2;
  assign T_735 = xact_is_builtin_type & T_734;
  assign T_736 = T_732 | T_735;
  assign T_737 = xact_union[8:1];
  assign T_739 = T_736 ? T_737 : {{7'd0}, 1'h0};
  assign T_740 = T_717 ? T_728_0 : T_739;
  assign T_767 = {T_740,1'h1};
  assign T_787 = 1'h1 ? {{3'd0}, T_767} : 12'h0;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_write_beat_client_xact_id = {{2'd0}, 1'h1};
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_write_beat_union = T_787;
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign GEN_0 = GEN_17;
  assign GEN_11 = GEN_234 == oacq_data_cnt ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign GEN_256 = {{1'd0}, 2'h2};
  assign GEN_12 = GEN_256 == oacq_data_cnt ? xact_wmask_buffer_2 : GEN_11;
  assign GEN_257 = {{1'd0}, 2'h3};
  assign GEN_13 = GEN_257 == oacq_data_cnt ? xact_wmask_buffer_3 : GEN_12;
  assign GEN_14 = 3'h4 == oacq_data_cnt ? xact_wmask_buffer_4 : GEN_13;
  assign GEN_15 = 3'h5 == oacq_data_cnt ? xact_wmask_buffer_5 : GEN_14;
  assign GEN_16 = 3'h6 == oacq_data_cnt ? xact_wmask_buffer_6 : GEN_15;
  assign GEN_17 = 3'h7 == oacq_data_cnt ? xact_wmask_buffer_7 : GEN_16;
  assign T_834 = {GEN_0,1'h1};
  assign T_852 = 1'h1 ? {{3'd0}, T_834} : 12'h0;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_block_client_xact_id = {{2'd0}, 1'h1};
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_block_union = T_852;
  assign oacq_write_block_data = GEN_1;
  assign GEN_1 = GEN_24;
  assign GEN_18 = GEN_234 == oacq_data_cnt ? xact_data_buffer_1 : xact_data_buffer_0;
  assign GEN_19 = GEN_256 == oacq_data_cnt ? xact_data_buffer_2 : GEN_18;
  assign GEN_20 = GEN_257 == oacq_data_cnt ? xact_data_buffer_3 : GEN_19;
  assign GEN_21 = 3'h4 == oacq_data_cnt ? xact_data_buffer_4 : GEN_20;
  assign GEN_22 = 3'h5 == oacq_data_cnt ? xact_data_buffer_5 : GEN_21;
  assign GEN_23 = 3'h6 == oacq_data_cnt ? xact_data_buffer_6 : GEN_22;
  assign GEN_24 = 3'h7 == oacq_data_cnt ? xact_data_buffer_7 : GEN_23;
  assign T_875 = xact_union[11:9];
  assign T_876 = xact_union[8:6];
  assign T_897 = {T_875,T_876};
  assign T_898 = {T_897,6'h0};
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign oacq_read_beat_client_xact_id = {{2'd0}, 1'h1};
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign oacq_read_beat_union = T_898;
  assign oacq_read_beat_data = {{4'd0}, 1'h0};
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_block_client_xact_id = {{2'd0}, 1'h1};
  assign oacq_read_block_addr_beat = {{2'd0}, 1'h0};
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_block_union = 12'h1c1;
  assign oacq_read_block_data = {{4'd0}, 1'h0};
  assign T_1013 = state == 3'h1;
  assign T_1014 = state == 3'h3;
  assign T_1015_addr_block = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign T_1015_client_xact_id = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign T_1015_addr_beat = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign T_1015_is_builtin_type = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign T_1015_a_type = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign T_1015_union = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign T_1015_data = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign T_1023_addr_block = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign T_1023_client_xact_id = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign T_1023_addr_beat = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign T_1023_is_builtin_type = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign T_1023_a_type = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign T_1023_union = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign T_1023_data = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign T_1031_addr_block = T_1014 ? T_1015_addr_block : T_1023_addr_block;
  assign T_1031_client_xact_id = T_1014 ? T_1015_client_xact_id : T_1023_client_xact_id;
  assign T_1031_addr_beat = T_1014 ? T_1015_addr_beat : T_1023_addr_beat;
  assign T_1031_is_builtin_type = T_1014 ? T_1015_is_builtin_type : T_1023_is_builtin_type;
  assign T_1031_a_type = T_1014 ? T_1015_a_type : T_1023_a_type;
  assign T_1031_union = T_1014 ? T_1015_union : T_1023_union;
  assign T_1031_data = T_1014 ? T_1015_data : T_1023_data;
  assign T_1039_addr_block = T_1013 ? oacq_probe_addr_block : T_1031_addr_block;
  assign T_1039_client_xact_id = T_1013 ? oacq_probe_client_xact_id : T_1031_client_xact_id;
  assign T_1039_addr_beat = T_1013 ? oacq_probe_addr_beat : T_1031_addr_beat;
  assign T_1039_is_builtin_type = T_1013 ? oacq_probe_is_builtin_type : T_1031_is_builtin_type;
  assign T_1039_a_type = T_1013 ? oacq_probe_a_type : T_1031_a_type;
  assign T_1039_union = T_1013 ? oacq_probe_union : T_1031_union;
  assign T_1039_data = T_1013 ? oacq_probe_data : T_1031_data;
  assign T_1056 = 3'h4 == xact_a_type;
  assign T_1057 = T_1056 ? 2'h0 : 2'h2;
  assign T_1058 = 3'h6 == xact_a_type;
  assign T_1059 = T_1058 ? 2'h0 : T_1057;
  assign T_1060 = 3'h5 == xact_a_type;
  assign T_1061 = T_1060 ? 2'h2 : T_1059;
  assign T_1062 = 3'h2 == xact_a_type;
  assign T_1063 = T_1062 ? 2'h0 : T_1061;
  assign T_1064 = 3'h0 == xact_a_type;
  assign T_1065 = T_1064 ? 2'h2 : T_1063;
  assign T_1066 = 3'h3 == xact_a_type;
  assign T_1067 = T_1066 ? 2'h0 : T_1065;
  assign T_1068 = 3'h1 == xact_a_type;
  assign T_1069 = T_1068 ? 2'h2 : T_1067;
  assign T_1070 = GEN_234 == xact_a_type;
  assign T_1071 = T_1070 ? 2'h0 : 2'h2;
  assign T_1072 = GEN_248 == xact_a_type;
  assign T_1073 = T_1072 ? 2'h1 : T_1071;
  assign T_1074 = xact_is_builtin_type ? T_1069 : T_1073;
  assign T_1079_addr_block = xact_addr_block;
  assign T_1079_p_type = T_1074;
  assign T_1079_client_id = {{1'd0}, 1'h0};
  assign T_1103 = T_1058 ? 3'h1 : 3'h3;
  assign T_1105 = T_1060 ? 3'h1 : T_1103;
  assign T_1107 = T_1056 ? 3'h4 : T_1105;
  assign T_1109 = T_1066 ? 3'h3 : T_1107;
  assign T_1111 = T_1062 ? 3'h3 : T_1109;
  assign T_1113 = T_1068 ? 3'h5 : T_1111;
  assign T_1115 = T_1064 ? 3'h4 : T_1113;
  assign T_1116 = xact_a_type == GEN_248;
  assign T_1121 = T_1116 ? 2'h0 : 2'h1;
  assign T_1122 = xact_is_builtin_type ? T_1115 : {{1'd0}, T_1121};
  assign T_1131_addr_beat = {{2'd0}, 1'h0};
  assign T_1131_client_xact_id = xact_client_xact_id;
  assign T_1131_manager_xact_id = {{2'd0}, 1'h1};
  assign T_1131_is_builtin_type = xact_is_builtin_type;
  assign T_1131_g_type = {{1'd0}, T_1122};
  assign T_1131_data = {{4'd0}, 1'h0};
  assign T_1131_client_id = xact_client_id;
  assign T_1143 = T_284 & collect_iacq_data;
  assign T_1145 = T_1143 & T_324;
  assign T_1146 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T_1147 = T_1145 & T_1146;
  assign T_1149 = T_1147 == 1'h0;
  assign T_1150 = T_1149 | reset;
  assign T_1152 = T_1150 == 1'h0;
  assign T_1157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T_1158 = T_1145 & T_1157;
  assign T_1160 = T_1158 == 1'h0;
  assign T_1161 = T_1160 | reset;
  assign T_1163 = T_1161 == 1'h0;
  assign T_1164 = state == 3'h0;
  assign T_1166 = T_1164 & T_324;
  assign T_1167 = T_1166 & io_alloc_iacq;
  assign T_1176_0 = 3'h3;
  assign T_1178 = T_1176_0 == io_inner_acquire_bits_a_type;
  assign T_1181 = io_inner_acquire_bits_is_builtin_type & T_1178;
  assign T_1182 = T_1167 & T_1181;
  assign T_1184 = io_inner_acquire_bits_addr_beat != GEN_248;
  assign T_1185 = T_1182 & T_1184;
  assign T_1187 = T_1185 == 1'h0;
  assign T_1188 = T_1187 | reset;
  assign T_1190 = T_1188 == 1'h0;
  assign GEN_2 = io_inner_acquire_bits_data;
  assign GEN_25 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_0;
  assign GEN_26 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_1;
  assign GEN_27 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_2;
  assign GEN_28 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_3;
  assign GEN_29 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_4;
  assign GEN_30 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_5;
  assign GEN_31 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_6;
  assign GEN_32 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_7;
  assign T_1193 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_1194 = io_inner_acquire_bits_is_builtin_type & T_1193;
  assign T_1205_0 = T_722;
  assign T_1208 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1209 = io_inner_acquire_bits_is_builtin_type & T_1208;
  assign T_1211 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1212 = io_inner_acquire_bits_is_builtin_type & T_1211;
  assign T_1213 = T_1209 | T_1212;
  assign T_1214 = io_inner_acquire_bits_union[8:1];
  assign T_1216 = T_1213 ? T_1214 : {{7'd0}, 1'h0};
  assign T_1217 = T_1194 ? T_1205_0 : T_1216;
  assign GEN_3 = T_1217;
  assign GEN_33 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_0;
  assign GEN_34 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_1;
  assign GEN_35 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_2;
  assign GEN_36 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_3;
  assign GEN_37 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_4;
  assign GEN_38 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_5;
  assign GEN_39 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_6;
  assign GEN_40 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_7;
  assign T_1220 = GEN_254 << io_inner_acquire_bits_addr_beat;
  assign T_1221 = iacq_data_valid | T_1220;
  assign GEN_42 = io_inner_acquire_valid ? GEN_25 : xact_data_buffer_0;
  assign GEN_43 = io_inner_acquire_valid ? GEN_26 : xact_data_buffer_1;
  assign GEN_44 = io_inner_acquire_valid ? GEN_27 : xact_data_buffer_2;
  assign GEN_45 = io_inner_acquire_valid ? GEN_28 : xact_data_buffer_3;
  assign GEN_46 = io_inner_acquire_valid ? GEN_29 : xact_data_buffer_4;
  assign GEN_47 = io_inner_acquire_valid ? GEN_30 : xact_data_buffer_5;
  assign GEN_48 = io_inner_acquire_valid ? GEN_31 : xact_data_buffer_6;
  assign GEN_49 = io_inner_acquire_valid ? GEN_32 : xact_data_buffer_7;
  assign GEN_52 = io_inner_acquire_valid ? GEN_33 : xact_wmask_buffer_0;
  assign GEN_53 = io_inner_acquire_valid ? GEN_34 : xact_wmask_buffer_1;
  assign GEN_54 = io_inner_acquire_valid ? GEN_35 : xact_wmask_buffer_2;
  assign GEN_55 = io_inner_acquire_valid ? GEN_36 : xact_wmask_buffer_3;
  assign GEN_56 = io_inner_acquire_valid ? GEN_37 : xact_wmask_buffer_4;
  assign GEN_57 = io_inner_acquire_valid ? GEN_38 : xact_wmask_buffer_5;
  assign GEN_58 = io_inner_acquire_valid ? GEN_39 : xact_wmask_buffer_6;
  assign GEN_59 = io_inner_acquire_valid ? GEN_40 : xact_wmask_buffer_7;
  assign GEN_60 = io_inner_acquire_valid ? T_1221 : iacq_data_valid;
  assign GEN_61 = iacq_data_done ? 1'h0 : collect_iacq_data;
  assign GEN_64 = collect_iacq_data ? GEN_42 : xact_data_buffer_0;
  assign GEN_65 = collect_iacq_data ? GEN_43 : xact_data_buffer_1;
  assign GEN_66 = collect_iacq_data ? GEN_44 : xact_data_buffer_2;
  assign GEN_67 = collect_iacq_data ? GEN_45 : xact_data_buffer_3;
  assign GEN_68 = collect_iacq_data ? GEN_46 : xact_data_buffer_4;
  assign GEN_69 = collect_iacq_data ? GEN_47 : xact_data_buffer_5;
  assign GEN_70 = collect_iacq_data ? GEN_48 : xact_data_buffer_6;
  assign GEN_71 = collect_iacq_data ? GEN_49 : xact_data_buffer_7;
  assign GEN_74 = collect_iacq_data ? GEN_52 : xact_wmask_buffer_0;
  assign GEN_75 = collect_iacq_data ? GEN_53 : xact_wmask_buffer_1;
  assign GEN_76 = collect_iacq_data ? GEN_54 : xact_wmask_buffer_2;
  assign GEN_77 = collect_iacq_data ? GEN_55 : xact_wmask_buffer_3;
  assign GEN_78 = collect_iacq_data ? GEN_56 : xact_wmask_buffer_4;
  assign GEN_79 = collect_iacq_data ? GEN_57 : xact_wmask_buffer_5;
  assign GEN_80 = collect_iacq_data ? GEN_58 : xact_wmask_buffer_6;
  assign GEN_81 = collect_iacq_data ? GEN_59 : xact_wmask_buffer_7;
  assign GEN_82 = collect_iacq_data ? GEN_60 : iacq_data_valid;
  assign GEN_83 = collect_iacq_data ? GEN_61 : collect_iacq_data;
  assign GEN_84 = io_outer_grant_valid ? 1'h0 : pending_ognt_ack;
  assign GEN_86 = pending_ognt_ack ? GEN_84 : pending_ognt_ack;
  assign T_1229 = 3'h0 == state;
  assign T_1231 = io_inner_acquire_valid & io_alloc_iacq;
  assign GEN_4 = io_inner_acquire_bits_data;
  assign T_1247_0 = T_722;
  assign T_1259 = T_1194 ? T_1247_0 : T_1216;
  assign GEN_5 = T_1259;
  assign T_1268_0 = 3'h3;
  assign T_1270 = T_1268_0 == io_inner_acquire_bits_a_type;
  assign T_1273 = io_inner_acquire_bits_is_builtin_type & T_1270;
  assign T_1282_0 = 3'h2;
  assign T_1282_1 = 3'h3;
  assign T_1282_2 = 3'h4;
  assign T_1284 = T_1282_0 == io_inner_acquire_bits_a_type;
  assign T_1285 = T_1282_1 == io_inner_acquire_bits_a_type;
  assign T_1286 = T_1282_2 == io_inner_acquire_bits_a_type;
  assign T_1289 = T_1284 | T_1285;
  assign T_1290 = T_1289 | T_1286;
  assign T_1291 = io_inner_acquire_bits_is_builtin_type & T_1290;
  assign GEN_276 = {{7'd0}, T_1291};
  assign T_1292 = GEN_276 << io_inner_acquire_bits_addr_beat;
  assign GEN_277 = {{3'd0}, 1'h0};
  assign T_1294 = mask_incoherent != GEN_277;
  assign T_1295 = mask_incoherent[0];
  assign T_1296 = mask_incoherent[1];
  assign T_1297 = mask_incoherent[2];
  assign T_1298 = mask_incoherent[3];
  assign T_1300 = {1'h0,T_1296};
  assign GEN_278 = {{1'd0}, T_1295};
  assign T_1301 = GEN_278 + T_1300;
  assign T_1302 = T_1301[1:0];
  assign T_1305 = {1'h0,T_1298};
  assign GEN_279 = {{1'd0}, T_1297};
  assign T_1306 = GEN_279 + T_1305;
  assign T_1307 = T_1306[1:0];
  assign T_1308 = {1'h0,T_1307};
  assign GEN_280 = {{1'd0}, T_1302};
  assign T_1309 = GEN_280 + T_1308;
  assign T_1310 = T_1309[2:0];
  assign GEN_103 = T_1294 ? mask_incoherent : {{3'd0}, pending_probes};
  assign GEN_104 = T_1294 ? T_1310 : {{2'd0}, release_count};
  assign T_1311 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign T_1312 = pending_outer_write_ ? 3'h3 : T_1311;
  assign T_1313 = T_1294 ? 3'h1 : T_1312;
  assign GEN_105 = T_1231 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_106 = T_1231 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign GEN_107 = T_1231 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign GEN_108 = T_1231 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign GEN_109 = T_1231 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign GEN_110 = T_1231 ? io_inner_acquire_bits_union : xact_union;
  assign GEN_111 = T_1231 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign GEN_113 = T_1231 ? GEN_4 : GEN_64;
  assign GEN_123 = T_1231 ? GEN_5 : GEN_74;
  assign GEN_132 = T_1231 ? T_1273 : GEN_83;
  assign GEN_136 = T_1231 ? T_1292 : GEN_82;
  assign GEN_137 = T_1231 ? GEN_103 : {{3'd0}, pending_probes};
  assign GEN_138 = T_1231 ? GEN_104 : {{2'd0}, release_count};
  assign GEN_139 = T_1231 ? T_1313 : state;
  assign GEN_140 = T_1229 ? 1'h1 : collect_iacq_data;
  assign GEN_141 = T_1229 ? GEN_105 : xact_addr_block;
  assign GEN_142 = T_1229 ? GEN_106 : xact_client_xact_id;
  assign GEN_143 = T_1229 ? GEN_107 : xact_addr_beat;
  assign GEN_144 = T_1229 ? GEN_108 : xact_is_builtin_type;
  assign GEN_145 = T_1229 ? GEN_109 : xact_a_type;
  assign GEN_146 = T_1229 ? GEN_110 : xact_union;
  assign GEN_147 = T_1229 ? GEN_111 : xact_client_id;
  assign GEN_149 = T_1229 ? GEN_113 : GEN_64;
  assign GEN_159 = T_1229 ? GEN_123 : GEN_74;
  assign GEN_168 = T_1229 ? GEN_132 : GEN_83;
  assign GEN_172 = T_1229 ? GEN_136 : GEN_82;
  assign GEN_173 = T_1229 ? GEN_137 : {{3'd0}, pending_probes};
  assign GEN_174 = T_1229 ? GEN_138 : {{2'd0}, release_count};
  assign GEN_175 = T_1229 ? GEN_139 : state;
  assign T_1314 = 3'h1 == state;
  assign GEN_281 = {{1'd0}, 1'h1};
  assign T_1318 = GEN_281 << 1'h0;
  assign T_1319 = ~ T_1318;
  assign GEN_282 = {{1'd0}, pending_probes};
  assign T_1320 = GEN_282 & T_1319;
  assign GEN_176 = io_inner_probe_ready ? {{2'd0}, T_1320} : GEN_173;
  assign T_1326_0 = 3'h0;
  assign T_1326_1 = 3'h1;
  assign T_1326_2 = 3'h2;
  assign T_1328 = T_1326_0 == io_inner_release_bits_r_type;
  assign T_1329 = T_1326_1 == io_inner_release_bits_r_type;
  assign T_1330 = T_1326_2 == io_inner_release_bits_r_type;
  assign T_1333 = T_1328 | T_1329;
  assign T_1334 = T_1333 | T_1330;
  assign T_1336 = T_1334 == 1'h0;
  assign T_1337 = T_1336 | io_outer_acquire_ready;
  assign T_1338 = T_1337 & io_matches_irel;
  assign T_1339 = io_inner_release_valid & io_matches_irel;
  assign T_1345_0 = 3'h0;
  assign T_1345_1 = 3'h1;
  assign T_1345_2 = 3'h2;
  assign T_1347 = T_1345_0 == io_inner_release_bits_r_type;
  assign T_1348 = T_1345_1 == io_inner_release_bits_r_type;
  assign T_1349 = T_1345_2 == io_inner_release_bits_r_type;
  assign T_1352 = T_1347 | T_1348;
  assign T_1353 = T_1352 | T_1349;
  assign T_1357 = release_count - 1'h1;
  assign T_1358 = T_1357[0:0];
  assign T_1361 = pending_outer_read ? 3'h2 : 3'h4;
  assign T_1362 = pending_outer_write ? 3'h3 : T_1361;
  assign GEN_177 = release_count ? T_1362 : GEN_175;
  assign GEN_178 = oacq_data_done ? 1'h1 : GEN_86;
  assign GEN_179 = oacq_data_done ? {{2'd0}, T_1358} : GEN_174;
  assign GEN_180 = oacq_data_done ? GEN_177 : GEN_175;
  assign GEN_181 = io_outer_acquire_ready ? GEN_178 : GEN_86;
  assign GEN_182 = io_outer_acquire_ready ? GEN_179 : GEN_174;
  assign GEN_183 = io_outer_acquire_ready ? GEN_180 : GEN_175;
  assign GEN_185 = T_1353 ? GEN_181 : GEN_86;
  assign GEN_186 = T_1353 ? GEN_182 : GEN_174;
  assign GEN_187 = T_1353 ? GEN_183 : GEN_175;
  assign T_1364 = T_1353 == 1'h0;
  assign GEN_188 = release_count ? T_1362 : GEN_187;
  assign GEN_189 = T_1364 ? {{2'd0}, T_1358} : GEN_186;
  assign GEN_190 = T_1364 ? GEN_188 : GEN_187;
  assign GEN_194 = T_1339 ? T_1353 : 1'h0;
  assign GEN_195 = T_1339 ? GEN_185 : GEN_86;
  assign GEN_196 = T_1339 ? GEN_189 : GEN_174;
  assign GEN_197 = T_1339 ? GEN_190 : GEN_175;
  assign GEN_198 = T_1314 ? pending_probes : 1'h0;
  assign GEN_199 = T_1314 ? GEN_176 : GEN_173;
  assign GEN_203 = T_1314 ? T_1338 : 1'h0;
  assign GEN_207 = T_1314 ? GEN_194 : 1'h0;
  assign GEN_208 = T_1314 ? GEN_195 : GEN_86;
  assign GEN_209 = T_1314 ? GEN_196 : GEN_174;
  assign GEN_210 = T_1314 ? GEN_197 : GEN_175;
  assign T_1372 = 3'h3 == state;
  assign T_1374 = pending_ognt_ack == 1'h0;
  assign T_1376 = collect_iacq_data == 1'h0;
  assign T_1377 = iacq_data_valid >> oacq_data_cnt;
  assign T_1378 = T_1377[0];
  assign T_1379 = T_1376 | T_1378;
  assign T_1380 = T_1374 & T_1379;
  assign T_1382 = pending_outer_read ? 3'h2 : 3'h5;
  assign GEN_211 = oacq_data_done ? 1'h1 : GEN_208;
  assign GEN_212 = oacq_data_done ? T_1382 : GEN_210;
  assign GEN_213 = T_1372 ? T_1380 : GEN_207;
  assign GEN_214 = T_1372 ? GEN_211 : GEN_208;
  assign GEN_215 = T_1372 ? GEN_212 : GEN_210;
  assign T_1383 = 3'h2 == state;
  assign GEN_216 = T_416 ? 3'h5 : GEN_215;
  assign GEN_217 = T_1383 ? T_1374 : GEN_213;
  assign GEN_218 = T_1383 ? GEN_216 : GEN_215;
  assign T_1387 = 3'h5 == state;
  assign GEN_283 = {{1'd0}, 3'h0};
  assign T_1392 = io_inner_grant_bits_g_type == GEN_283;
  assign T_1393 = io_inner_grant_bits_is_builtin_type & T_1392;
  assign T_1395 = T_1393 == 1'h0;
  assign T_1397 = T_1395 ? 3'h6 : 3'h0;
  assign GEN_219 = ignt_data_done ? T_1397 : GEN_218;
  assign GEN_220 = T_1387 ? io_inner_grant_ready : pending_ognt_ack;
  assign GEN_221 = T_1387 ? io_outer_grant_valid : 1'h0;
  assign GEN_222 = T_1387 ? GEN_219 : GEN_218;
  assign T_1398 = 3'h4 == state;
  assign GEN_223 = io_inner_grant_ready ? T_1397 : GEN_222;
  assign GEN_224 = T_1398 ? 1'h1 : GEN_221;
  assign GEN_225 = T_1398 ? GEN_223 : GEN_222;
  assign T_1410 = 3'h6 == state;
  assign GEN_226 = io_inner_finish_valid ? 3'h0 : GEN_225;
  assign GEN_228 = T_1410 ? GEN_226 : GEN_225;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_41 = {1{$random}};
  state = GEN_41[2:0];
  GEN_50 = {1{$random}};
  xact_addr_block = GEN_50[25:0];
  GEN_51 = {1{$random}};
  xact_client_xact_id = GEN_51[1:0];
  GEN_62 = {1{$random}};
  xact_addr_beat = GEN_62[2:0];
  GEN_63 = {1{$random}};
  xact_is_builtin_type = GEN_63[0:0];
  GEN_72 = {1{$random}};
  xact_a_type = GEN_72[2:0];
  GEN_73 = {1{$random}};
  xact_union = GEN_73[11:0];
  GEN_85 = {1{$random}};
  xact_data_buffer_0 = GEN_85[4:0];
  GEN_87 = {1{$random}};
  xact_data_buffer_1 = GEN_87[4:0];
  GEN_88 = {1{$random}};
  xact_data_buffer_2 = GEN_88[4:0];
  GEN_89 = {1{$random}};
  xact_data_buffer_3 = GEN_89[4:0];
  GEN_90 = {1{$random}};
  xact_data_buffer_4 = GEN_90[4:0];
  GEN_91 = {1{$random}};
  xact_data_buffer_5 = GEN_91[4:0];
  GEN_92 = {1{$random}};
  xact_data_buffer_6 = GEN_92[4:0];
  GEN_93 = {1{$random}};
  xact_data_buffer_7 = GEN_93[4:0];
  GEN_94 = {1{$random}};
  xact_wmask_buffer_0 = GEN_94[7:0];
  GEN_95 = {1{$random}};
  xact_wmask_buffer_1 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  xact_wmask_buffer_2 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  xact_wmask_buffer_3 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  xact_wmask_buffer_4 = GEN_98[7:0];
  GEN_99 = {1{$random}};
  xact_wmask_buffer_5 = GEN_99[7:0];
  GEN_100 = {1{$random}};
  xact_wmask_buffer_6 = GEN_100[7:0];
  GEN_101 = {1{$random}};
  xact_wmask_buffer_7 = GEN_101[7:0];
  GEN_102 = {1{$random}};
  xact_client_id = GEN_102[1:0];
  GEN_112 = {1{$random}};
  release_count = GEN_112[0:0];
  GEN_114 = {1{$random}};
  pending_probes = GEN_114[0:0];
  GEN_115 = {1{$random}};
  collect_iacq_data = GEN_115[0:0];
  GEN_116 = {1{$random}};
  iacq_data_valid = GEN_116[7:0];
  GEN_117 = {1{$random}};
  T_342 = GEN_117[2:0];
  GEN_118 = {1{$random}};
  T_370 = GEN_118[2:0];
  GEN_119 = {1{$random}};
  T_408 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  T_433 = GEN_120[2:0];
  GEN_121 = {1{$random}};
  T_468 = GEN_121[2:0];
  GEN_122 = {1{$random}};
  pending_ognt_ack = GEN_122[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_228;
    end
    if(1'h0) begin
    end else begin
      xact_addr_block <= GEN_141;
    end
    if(1'h0) begin
    end else begin
      xact_client_xact_id <= GEN_142;
    end
    if(1'h0) begin
    end else begin
      xact_addr_beat <= GEN_143;
    end
    if(1'h0) begin
    end else begin
      xact_is_builtin_type <= GEN_144;
    end
    if(1'h0) begin
    end else begin
      xact_a_type <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      xact_union <= GEN_146;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_0 <= GEN_149;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_1 <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_2 <= GEN_66;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_3 <= GEN_67;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_4 <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_5 <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_6 <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_7 <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_0 <= GEN_159;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_1 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_2 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_3 <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_4 <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_5 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_6 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_7 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      xact_client_id <= GEN_147;
    end
    if(reset) begin
      release_count <= 1'h0;
    end else begin
      release_count <= GEN_209[0];
    end
    if(reset) begin
      pending_probes <= 1'h0;
    end else begin
      pending_probes <= GEN_199[0];
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else begin
      collect_iacq_data <= GEN_168;
    end
    if(reset) begin
      iacq_data_valid <= 8'h0;
    end else begin
      iacq_data_valid <= GEN_172;
    end
    if(reset) begin
      T_342 <= 3'h0;
    end else begin
      T_342 <= GEN_6;
    end
    if(reset) begin
      T_370 <= 3'h0;
    end else begin
      T_370 <= GEN_7;
    end
    if(reset) begin
      T_408 <= 3'h0;
    end else begin
      T_408 <= GEN_8;
    end
    if(reset) begin
      T_433 <= 3'h0;
    end else begin
      T_433 <= GEN_9;
    end
    if(reset) begin
      T_468 <= 3'h0;
    end else begin
      T_468 <= GEN_10;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else begin
      pending_ognt_ack <= GEN_214;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics or prefetches\n    at broadcast.scala:203 assert(!(state =/= s_idle && xact.isBuiltInType() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different network source than initial request.\n    at broadcast.scala:285 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different client transaction than initial request.\n    at broadcast.scala:289 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at broadcast.scala:293 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module BroadcastAcquireTracker_28(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [4:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [4:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [4:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [4:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [4:0] io_outer_grant_bits_data,
  output  io_matches_iacq,
  output  io_matches_irel,
  output  io_matches_oprb,
  input   io_alloc_iacq,
  input   io_alloc_irel,
  input   io_alloc_oprb
);
  reg [2:0] state;
  reg [31:0] GEN_41;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_50;
  reg [1:0] xact_client_xact_id;
  reg [31:0] GEN_51;
  reg [2:0] xact_addr_beat;
  reg [31:0] GEN_62;
  reg  xact_is_builtin_type;
  reg [31:0] GEN_63;
  reg [2:0] xact_a_type;
  reg [31:0] GEN_72;
  reg [11:0] xact_union;
  reg [31:0] GEN_73;
  reg [4:0] xact_data_buffer_0;
  reg [31:0] GEN_85;
  reg [4:0] xact_data_buffer_1;
  reg [31:0] GEN_87;
  reg [4:0] xact_data_buffer_2;
  reg [31:0] GEN_88;
  reg [4:0] xact_data_buffer_3;
  reg [31:0] GEN_89;
  reg [4:0] xact_data_buffer_4;
  reg [31:0] GEN_90;
  reg [4:0] xact_data_buffer_5;
  reg [31:0] GEN_91;
  reg [4:0] xact_data_buffer_6;
  reg [31:0] GEN_92;
  reg [4:0] xact_data_buffer_7;
  reg [31:0] GEN_93;
  reg [7:0] xact_wmask_buffer_0;
  reg [31:0] GEN_94;
  reg [7:0] xact_wmask_buffer_1;
  reg [31:0] GEN_95;
  reg [7:0] xact_wmask_buffer_2;
  reg [31:0] GEN_96;
  reg [7:0] xact_wmask_buffer_3;
  reg [31:0] GEN_97;
  reg [7:0] xact_wmask_buffer_4;
  reg [31:0] GEN_98;
  reg [7:0] xact_wmask_buffer_5;
  reg [31:0] GEN_99;
  reg [7:0] xact_wmask_buffer_6;
  reg [31:0] GEN_100;
  reg [7:0] xact_wmask_buffer_7;
  reg [31:0] GEN_101;
  reg [1:0] xact_client_id;
  reg [31:0] GEN_102;
  wire  coh_sharers;
  wire  T_284;
  wire  T_285;
  wire [2:0] T_294_0;
  wire [2:0] T_294_1;
  wire [2:0] T_294_2;
  wire  T_296;
  wire  T_297;
  wire  T_298;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_305;
  wire  T_306;
  wire  T_308;
  reg  release_count;
  reg [31:0] GEN_112;
  reg  pending_probes;
  reg [31:0] GEN_114;
  wire  GEN_229;
  wire  T_313;
  wire [3:0] GEN_230;
  wire [3:0] T_316;
  wire  T_318;
  wire [3:0] GEN_232;
  wire [3:0] T_319;
  wire [3:0] T_320;
  wire  T_321;
  wire [3:0] GEN_233;
  wire [3:0] mask_incoherent;
  reg  collect_iacq_data;
  reg [31:0] GEN_115;
  reg [7:0] iacq_data_valid;
  reg [31:0] GEN_116;
  wire  T_324;
  wire [2:0] T_334_0;
  wire  T_336;
  wire  T_339;
  wire  T_340;
  reg [2:0] T_342;
  reg [31:0] GEN_117;
  wire  T_344;
  wire [2:0] GEN_234;
  wire [3:0] T_346;
  wire [2:0] T_347;
  wire [2:0] GEN_6;
  wire  T_348;
  wire  iacq_data_done;
  wire  T_350;
  wire [2:0] T_358_0;
  wire [2:0] T_358_1;
  wire [2:0] T_358_2;
  wire  T_360;
  wire  T_361;
  wire  T_362;
  wire  T_365;
  wire  T_366;
  wire  T_368;
  reg [2:0] T_370;
  reg [31:0] GEN_118;
  wire [3:0] T_374;
  wire [2:0] T_375;
  wire [2:0] GEN_7;
  wire  T_379;
  wire [2:0] T_387_0;
  wire [3:0] GEN_236;
  wire  T_389;
  wire [1:0] T_397_0;
  wire [1:0] T_397_1;
  wire [3:0] GEN_237;
  wire  T_399;
  wire [3:0] GEN_238;
  wire  T_400;
  wire  T_403;
  wire  T_404;
  wire  T_406;
  reg [2:0] T_408;
  reg [31:0] GEN_119;
  wire  T_410;
  wire [3:0] T_412;
  wire [2:0] T_413;
  wire [2:0] GEN_8;
  wire  T_414;
  wire  ignt_data_done;
  wire  T_416;
  wire [2:0] T_425_0;
  wire  T_427;
  wire  T_430;
  wire  T_431;
  reg [2:0] T_433;
  reg [31:0] GEN_120;
  wire  T_435;
  wire [3:0] T_437;
  wire [2:0] T_438;
  wire [2:0] GEN_9;
  wire  T_439;
  wire [2:0] oacq_data_cnt;
  wire  oacq_data_done;
  wire  T_440;
  wire [2:0] T_449_0;
  wire [3:0] GEN_241;
  wire  T_451;
  wire  T_459_0;
  wire [3:0] GEN_242;
  wire  T_461;
  wire  T_464;
  wire  T_466;
  reg [2:0] T_468;
  reg [31:0] GEN_121;
  wire [3:0] T_472;
  wire [2:0] T_473;
  wire [2:0] GEN_10;
  reg  pending_ognt_ack;
  reg [31:0] GEN_122;
  wire [2:0] T_485_0;
  wire [2:0] T_485_1;
  wire [2:0] T_485_2;
  wire  T_487;
  wire  T_488;
  wire  T_489;
  wire  T_492;
  wire  T_493;
  wire  pending_outer_write;
  wire [2:0] T_502_0;
  wire [2:0] T_502_1;
  wire [2:0] T_502_2;
  wire  T_504;
  wire  T_505;
  wire  T_506;
  wire  T_509;
  wire  T_510;
  wire  pending_outer_write_;
  wire [2:0] T_518_0;
  wire [2:0] T_518_1;
  wire [3:0] GEN_244;
  wire  T_520;
  wire [3:0] GEN_245;
  wire  T_521;
  wire  T_524;
  wire [1:0] T_530_0;
  wire [1:0] T_530_1;
  wire [3:0] GEN_246;
  wire  T_532;
  wire [3:0] GEN_247;
  wire  T_533;
  wire  T_536;
  wire  pending_outer_read;
  wire  T_555;
  wire [2:0] T_556;
  wire  T_557;
  wire [2:0] T_558;
  wire  T_559;
  wire [2:0] T_560;
  wire  T_561;
  wire [2:0] T_562;
  wire  T_563;
  wire [2:0] T_564;
  wire  T_565;
  wire [2:0] T_566;
  wire  T_567;
  wire [2:0] T_568;
  wire [2:0] GEN_248;
  wire  T_569;
  wire [1:0] T_574;
  wire [2:0] T_575;
  wire [2:0] T_584_addr_beat;
  wire [1:0] T_584_client_xact_id;
  wire [2:0] T_584_manager_xact_id;
  wire  T_584_is_builtin_type;
  wire [3:0] T_584_g_type;
  wire [4:0] T_584_data;
  wire [1:0] T_584_client_id;
  wire [2:0] T_599_0;
  wire [2:0] T_599_1;
  wire [3:0] GEN_249;
  wire  T_601;
  wire [3:0] GEN_250;
  wire  T_602;
  wire  T_605;
  wire [1:0] T_611_0;
  wire [1:0] T_611_1;
  wire [3:0] GEN_251;
  wire  T_613;
  wire [3:0] GEN_252;
  wire  T_614;
  wire  T_617;
  wire  pending_outer_read_;
  wire [2:0] T_626_0;
  wire [2:0] T_626_1;
  wire [2:0] T_626_2;
  wire  T_628;
  wire  T_629;
  wire  T_630;
  wire  T_633;
  wire  T_634;
  wire  subblock_type;
  wire  T_636;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire  T_642;
  wire  T_643;
  wire [7:0] GEN_253;
  wire [7:0] T_649;
  wire [8:0] T_674;
  wire [11:0] T_692;
  wire [25:0] oacq_probe_addr_block;
  wire [2:0] oacq_probe_client_xact_id;
  wire [2:0] oacq_probe_addr_beat;
  wire  oacq_probe_is_builtin_type;
  wire [2:0] oacq_probe_a_type;
  wire [11:0] oacq_probe_union;
  wire [4:0] oacq_probe_data;
  wire  T_716;
  wire  T_717;
  wire [7:0] GEN_254;
  wire [8:0] T_721;
  wire [7:0] T_722;
  wire [7:0] T_728_0;
  wire  T_731;
  wire  T_732;
  wire  T_734;
  wire  T_735;
  wire  T_736;
  wire [7:0] T_737;
  wire [7:0] T_739;
  wire [7:0] T_740;
  wire [8:0] T_767;
  wire [11:0] T_787;
  wire [25:0] oacq_write_beat_addr_block;
  wire [2:0] oacq_write_beat_client_xact_id;
  wire [2:0] oacq_write_beat_addr_beat;
  wire  oacq_write_beat_is_builtin_type;
  wire [2:0] oacq_write_beat_a_type;
  wire [11:0] oacq_write_beat_union;
  wire [4:0] oacq_write_beat_data;
  wire [7:0] GEN_0;
  wire [7:0] GEN_11;
  wire [2:0] GEN_256;
  wire [7:0] GEN_12;
  wire [2:0] GEN_257;
  wire [7:0] GEN_13;
  wire [7:0] GEN_14;
  wire [7:0] GEN_15;
  wire [7:0] GEN_16;
  wire [7:0] GEN_17;
  wire [8:0] T_834;
  wire [11:0] T_852;
  wire [25:0] oacq_write_block_addr_block;
  wire [2:0] oacq_write_block_client_xact_id;
  wire [2:0] oacq_write_block_addr_beat;
  wire  oacq_write_block_is_builtin_type;
  wire [2:0] oacq_write_block_a_type;
  wire [11:0] oacq_write_block_union;
  wire [4:0] oacq_write_block_data;
  wire [4:0] GEN_1;
  wire [4:0] GEN_18;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [2:0] T_875;
  wire [2:0] T_876;
  wire [5:0] T_897;
  wire [11:0] T_898;
  wire [25:0] oacq_read_beat_addr_block;
  wire [2:0] oacq_read_beat_client_xact_id;
  wire [2:0] oacq_read_beat_addr_beat;
  wire  oacq_read_beat_is_builtin_type;
  wire [2:0] oacq_read_beat_a_type;
  wire [11:0] oacq_read_beat_union;
  wire [4:0] oacq_read_beat_data;
  wire [25:0] oacq_read_block_addr_block;
  wire [2:0] oacq_read_block_client_xact_id;
  wire [2:0] oacq_read_block_addr_beat;
  wire  oacq_read_block_is_builtin_type;
  wire [2:0] oacq_read_block_a_type;
  wire [11:0] oacq_read_block_union;
  wire [4:0] oacq_read_block_data;
  wire  T_1013;
  wire  T_1014;
  wire [25:0] T_1015_addr_block;
  wire [2:0] T_1015_client_xact_id;
  wire [2:0] T_1015_addr_beat;
  wire  T_1015_is_builtin_type;
  wire [2:0] T_1015_a_type;
  wire [11:0] T_1015_union;
  wire [4:0] T_1015_data;
  wire [25:0] T_1023_addr_block;
  wire [2:0] T_1023_client_xact_id;
  wire [2:0] T_1023_addr_beat;
  wire  T_1023_is_builtin_type;
  wire [2:0] T_1023_a_type;
  wire [11:0] T_1023_union;
  wire [4:0] T_1023_data;
  wire [25:0] T_1031_addr_block;
  wire [2:0] T_1031_client_xact_id;
  wire [2:0] T_1031_addr_beat;
  wire  T_1031_is_builtin_type;
  wire [2:0] T_1031_a_type;
  wire [11:0] T_1031_union;
  wire [4:0] T_1031_data;
  wire [25:0] T_1039_addr_block;
  wire [2:0] T_1039_client_xact_id;
  wire [2:0] T_1039_addr_beat;
  wire  T_1039_is_builtin_type;
  wire [2:0] T_1039_a_type;
  wire [11:0] T_1039_union;
  wire [4:0] T_1039_data;
  wire  T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire  T_1060;
  wire [1:0] T_1061;
  wire  T_1062;
  wire [1:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire  T_1066;
  wire [1:0] T_1067;
  wire  T_1068;
  wire [1:0] T_1069;
  wire  T_1070;
  wire [1:0] T_1071;
  wire  T_1072;
  wire [1:0] T_1073;
  wire [1:0] T_1074;
  wire [25:0] T_1079_addr_block;
  wire [1:0] T_1079_p_type;
  wire [1:0] T_1079_client_id;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1107;
  wire [2:0] T_1109;
  wire [2:0] T_1111;
  wire [2:0] T_1113;
  wire [2:0] T_1115;
  wire  T_1116;
  wire [1:0] T_1121;
  wire [2:0] T_1122;
  wire [2:0] T_1131_addr_beat;
  wire [1:0] T_1131_client_xact_id;
  wire [2:0] T_1131_manager_xact_id;
  wire  T_1131_is_builtin_type;
  wire [3:0] T_1131_g_type;
  wire [4:0] T_1131_data;
  wire [1:0] T_1131_client_id;
  wire  T_1143;
  wire  T_1145;
  wire  T_1146;
  wire  T_1147;
  wire  T_1149;
  wire  T_1150;
  wire  T_1152;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire [2:0] T_1176_0;
  wire  T_1178;
  wire  T_1181;
  wire  T_1182;
  wire  T_1184;
  wire  T_1185;
  wire  T_1187;
  wire  T_1188;
  wire  T_1190;
  wire [4:0] GEN_2;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire [4:0] GEN_29;
  wire [4:0] GEN_30;
  wire [4:0] GEN_31;
  wire [4:0] GEN_32;
  wire  T_1193;
  wire  T_1194;
  wire [7:0] T_1205_0;
  wire  T_1208;
  wire  T_1209;
  wire  T_1211;
  wire  T_1212;
  wire  T_1213;
  wire [7:0] T_1214;
  wire [7:0] T_1216;
  wire [7:0] T_1217;
  wire [7:0] GEN_3;
  wire [7:0] GEN_33;
  wire [7:0] GEN_34;
  wire [7:0] GEN_35;
  wire [7:0] GEN_36;
  wire [7:0] GEN_37;
  wire [7:0] GEN_38;
  wire [7:0] GEN_39;
  wire [7:0] GEN_40;
  wire [7:0] T_1220;
  wire [7:0] T_1221;
  wire [4:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [4:0] GEN_45;
  wire [4:0] GEN_46;
  wire [4:0] GEN_47;
  wire [4:0] GEN_48;
  wire [4:0] GEN_49;
  wire [7:0] GEN_52;
  wire [7:0] GEN_53;
  wire [7:0] GEN_54;
  wire [7:0] GEN_55;
  wire [7:0] GEN_56;
  wire [7:0] GEN_57;
  wire [7:0] GEN_58;
  wire [7:0] GEN_59;
  wire [7:0] GEN_60;
  wire  GEN_61;
  wire [4:0] GEN_64;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] GEN_71;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire [7:0] GEN_78;
  wire [7:0] GEN_79;
  wire [7:0] GEN_80;
  wire [7:0] GEN_81;
  wire [7:0] GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_86;
  wire  T_1229;
  wire  T_1231;
  wire [4:0] GEN_4;
  wire [7:0] T_1247_0;
  wire [7:0] T_1259;
  wire [7:0] GEN_5;
  wire [2:0] T_1268_0;
  wire  T_1270;
  wire  T_1273;
  wire [2:0] T_1282_0;
  wire [2:0] T_1282_1;
  wire [2:0] T_1282_2;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1289;
  wire  T_1290;
  wire  T_1291;
  wire [7:0] GEN_276;
  wire [7:0] T_1292;
  wire [3:0] GEN_277;
  wire  T_1294;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire  T_1298;
  wire [1:0] T_1300;
  wire [1:0] GEN_278;
  wire [2:0] T_1301;
  wire [1:0] T_1302;
  wire [1:0] T_1305;
  wire [1:0] GEN_279;
  wire [2:0] T_1306;
  wire [1:0] T_1307;
  wire [2:0] T_1308;
  wire [2:0] GEN_280;
  wire [3:0] T_1309;
  wire [2:0] T_1310;
  wire [3:0] GEN_103;
  wire [2:0] GEN_104;
  wire [2:0] T_1311;
  wire [2:0] T_1312;
  wire [2:0] T_1313;
  wire [25:0] GEN_105;
  wire [1:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire [2:0] GEN_109;
  wire [11:0] GEN_110;
  wire [1:0] GEN_111;
  wire [4:0] GEN_113;
  wire [7:0] GEN_123;
  wire  GEN_132;
  wire [7:0] GEN_136;
  wire [3:0] GEN_137;
  wire [2:0] GEN_138;
  wire [2:0] GEN_139;
  wire  GEN_140;
  wire [25:0] GEN_141;
  wire [1:0] GEN_142;
  wire [2:0] GEN_143;
  wire  GEN_144;
  wire [2:0] GEN_145;
  wire [11:0] GEN_146;
  wire [1:0] GEN_147;
  wire [4:0] GEN_149;
  wire [7:0] GEN_159;
  wire  GEN_168;
  wire [7:0] GEN_172;
  wire [3:0] GEN_173;
  wire [2:0] GEN_174;
  wire [2:0] GEN_175;
  wire  T_1314;
  wire [1:0] GEN_281;
  wire [1:0] T_1318;
  wire [1:0] T_1319;
  wire [1:0] GEN_282;
  wire [1:0] T_1320;
  wire [3:0] GEN_176;
  wire [2:0] T_1326_0;
  wire [2:0] T_1326_1;
  wire [2:0] T_1326_2;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire  T_1339;
  wire [2:0] T_1345_0;
  wire [2:0] T_1345_1;
  wire [2:0] T_1345_2;
  wire  T_1347;
  wire  T_1348;
  wire  T_1349;
  wire  T_1352;
  wire  T_1353;
  wire [1:0] T_1357;
  wire  T_1358;
  wire [2:0] T_1361;
  wire [2:0] T_1362;
  wire [2:0] GEN_177;
  wire  GEN_178;
  wire [2:0] GEN_179;
  wire [2:0] GEN_180;
  wire  GEN_181;
  wire [2:0] GEN_182;
  wire [2:0] GEN_183;
  wire  GEN_185;
  wire [2:0] GEN_186;
  wire [2:0] GEN_187;
  wire  T_1364;
  wire [2:0] GEN_188;
  wire [2:0] GEN_189;
  wire [2:0] GEN_190;
  wire  GEN_194;
  wire  GEN_195;
  wire [2:0] GEN_196;
  wire [2:0] GEN_197;
  wire  GEN_198;
  wire [3:0] GEN_199;
  wire  GEN_203;
  wire  GEN_207;
  wire  GEN_208;
  wire [2:0] GEN_209;
  wire [2:0] GEN_210;
  wire  T_1372;
  wire  T_1374;
  wire  T_1376;
  wire [7:0] T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1380;
  wire [2:0] T_1382;
  wire  GEN_211;
  wire [2:0] GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire [2:0] GEN_215;
  wire  T_1383;
  wire [2:0] GEN_216;
  wire  GEN_217;
  wire [2:0] GEN_218;
  wire  T_1387;
  wire [3:0] GEN_283;
  wire  T_1392;
  wire  T_1393;
  wire  T_1395;
  wire [2:0] T_1397;
  wire [2:0] GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire [2:0] GEN_222;
  wire  T_1398;
  wire [2:0] GEN_223;
  wire  GEN_224;
  wire [2:0] GEN_225;
  wire  T_1410;
  wire [2:0] GEN_226;
  wire [2:0] GEN_228;
  assign io_inner_acquire_ready = GEN_140;
  assign io_inner_grant_valid = GEN_224;
  assign io_inner_grant_bits_addr_beat = T_1131_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1131_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1131_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1131_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1131_g_type;
  assign io_inner_grant_bits_data = T_1131_data;
  assign io_inner_grant_bits_client_id = T_1131_client_id;
  assign io_inner_finish_ready = T_1410;
  assign io_inner_probe_valid = GEN_198;
  assign io_inner_probe_bits_addr_block = T_1079_addr_block;
  assign io_inner_probe_bits_p_type = T_1079_p_type;
  assign io_inner_probe_bits_client_id = T_1079_client_id;
  assign io_inner_release_ready = GEN_203;
  assign io_outer_acquire_valid = GEN_217;
  assign io_outer_acquire_bits_addr_block = T_1039_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_1039_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_1039_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_1039_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_1039_a_type;
  assign io_outer_acquire_bits_union = T_1039_union;
  assign io_outer_acquire_bits_data = T_1039_data;
  assign io_outer_grant_ready = GEN_220;
  assign io_matches_iacq = T_637;
  assign io_matches_irel = T_643;
  assign io_matches_oprb = 1'h0;
  assign coh_sharers = 1'h0;
  assign T_284 = state != 3'h0;
  assign T_285 = T_284 & xact_is_builtin_type;
  assign T_294_0 = 3'h4;
  assign T_294_1 = 3'h5;
  assign T_294_2 = 3'h6;
  assign T_296 = T_294_0 == xact_a_type;
  assign T_297 = T_294_1 == xact_a_type;
  assign T_298 = T_294_2 == xact_a_type;
  assign T_301 = T_296 | T_297;
  assign T_302 = T_301 | T_298;
  assign T_303 = T_285 & T_302;
  assign T_305 = T_303 == 1'h0;
  assign T_306 = T_305 | reset;
  assign T_308 = T_306 == 1'h0;
  assign GEN_229 = $signed(1'h1);
  assign T_313 = $unsigned(GEN_229);
  assign GEN_230 = {{3'd0}, 1'h1};
  assign T_316 = GEN_230 << io_inner_acquire_bits_client_id;
  assign T_318 = ~ T_313;
  assign GEN_232 = {{3'd0}, T_318};
  assign T_319 = GEN_232 | T_316;
  assign T_320 = ~ T_319;
  assign T_321 = ~ io_incoherent_0;
  assign GEN_233 = {{3'd0}, T_321};
  assign mask_incoherent = T_320 & GEN_233;
  assign T_324 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_334_0 = 3'h3;
  assign T_336 = T_334_0 == io_inner_acquire_bits_a_type;
  assign T_339 = io_inner_acquire_bits_is_builtin_type & T_336;
  assign T_340 = T_324 & T_339;
  assign T_344 = T_342 == 3'h7;
  assign GEN_234 = {{2'd0}, 1'h1};
  assign T_346 = T_342 + GEN_234;
  assign T_347 = T_346[2:0];
  assign GEN_6 = T_340 ? T_347 : T_342;
  assign T_348 = T_340 & T_344;
  assign iacq_data_done = T_339 ? T_348 : T_324;
  assign T_350 = io_inner_release_ready & io_inner_release_valid;
  assign T_358_0 = 3'h0;
  assign T_358_1 = 3'h1;
  assign T_358_2 = 3'h2;
  assign T_360 = T_358_0 == io_inner_release_bits_r_type;
  assign T_361 = T_358_1 == io_inner_release_bits_r_type;
  assign T_362 = T_358_2 == io_inner_release_bits_r_type;
  assign T_365 = T_360 | T_361;
  assign T_366 = T_365 | T_362;
  assign T_368 = T_350 & T_366;
  assign T_374 = T_370 + GEN_234;
  assign T_375 = T_374[2:0];
  assign GEN_7 = T_368 ? T_375 : T_370;
  assign T_379 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_387_0 = 3'h5;
  assign GEN_236 = {{1'd0}, T_387_0};
  assign T_389 = GEN_236 == io_inner_grant_bits_g_type;
  assign T_397_0 = 2'h0;
  assign T_397_1 = 2'h1;
  assign GEN_237 = {{2'd0}, T_397_0};
  assign T_399 = GEN_237 == io_inner_grant_bits_g_type;
  assign GEN_238 = {{2'd0}, T_397_1};
  assign T_400 = GEN_238 == io_inner_grant_bits_g_type;
  assign T_403 = T_399 | T_400;
  assign T_404 = io_inner_grant_bits_is_builtin_type ? T_389 : T_403;
  assign T_406 = T_379 & T_404;
  assign T_410 = T_408 == 3'h7;
  assign T_412 = T_408 + GEN_234;
  assign T_413 = T_412[2:0];
  assign GEN_8 = T_406 ? T_413 : T_408;
  assign T_414 = T_406 & T_410;
  assign ignt_data_done = T_404 ? T_414 : T_379;
  assign T_416 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_425_0 = 3'h3;
  assign T_427 = T_425_0 == io_outer_acquire_bits_a_type;
  assign T_430 = io_outer_acquire_bits_is_builtin_type & T_427;
  assign T_431 = T_416 & T_430;
  assign T_435 = T_433 == 3'h7;
  assign T_437 = T_433 + GEN_234;
  assign T_438 = T_437[2:0];
  assign GEN_9 = T_431 ? T_438 : T_433;
  assign T_439 = T_431 & T_435;
  assign oacq_data_cnt = T_430 ? T_433 : {{2'd0}, 1'h0};
  assign oacq_data_done = T_430 ? T_439 : T_416;
  assign T_440 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_449_0 = 3'h5;
  assign GEN_241 = {{1'd0}, T_449_0};
  assign T_451 = GEN_241 == io_outer_grant_bits_g_type;
  assign T_459_0 = 1'h0;
  assign GEN_242 = {{3'd0}, T_459_0};
  assign T_461 = GEN_242 == io_outer_grant_bits_g_type;
  assign T_464 = io_outer_grant_bits_is_builtin_type ? T_451 : T_461;
  assign T_466 = T_440 & T_464;
  assign T_472 = T_468 + GEN_234;
  assign T_473 = T_472[2:0];
  assign GEN_10 = T_466 ? T_473 : T_468;
  assign T_485_0 = 3'h2;
  assign T_485_1 = 3'h3;
  assign T_485_2 = 3'h4;
  assign T_487 = T_485_0 == xact_a_type;
  assign T_488 = T_485_1 == xact_a_type;
  assign T_489 = T_485_2 == xact_a_type;
  assign T_492 = T_487 | T_488;
  assign T_493 = T_492 | T_489;
  assign pending_outer_write = xact_is_builtin_type & T_493;
  assign T_502_0 = 3'h2;
  assign T_502_1 = 3'h3;
  assign T_502_2 = 3'h4;
  assign T_504 = T_502_0 == io_inner_acquire_bits_a_type;
  assign T_505 = T_502_1 == io_inner_acquire_bits_a_type;
  assign T_506 = T_502_2 == io_inner_acquire_bits_a_type;
  assign T_509 = T_504 | T_505;
  assign T_510 = T_509 | T_506;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T_510;
  assign T_518_0 = 3'h5;
  assign T_518_1 = 3'h4;
  assign GEN_244 = {{1'd0}, T_518_0};
  assign T_520 = GEN_244 == io_inner_grant_bits_g_type;
  assign GEN_245 = {{1'd0}, T_518_1};
  assign T_521 = GEN_245 == io_inner_grant_bits_g_type;
  assign T_524 = T_520 | T_521;
  assign T_530_0 = 2'h0;
  assign T_530_1 = 2'h1;
  assign GEN_246 = {{2'd0}, T_530_0};
  assign T_532 = GEN_246 == io_inner_grant_bits_g_type;
  assign GEN_247 = {{2'd0}, T_530_1};
  assign T_533 = GEN_247 == io_inner_grant_bits_g_type;
  assign T_536 = T_532 | T_533;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T_524 : T_536;
  assign T_555 = 3'h6 == io_inner_acquire_bits_a_type;
  assign T_556 = T_555 ? 3'h1 : 3'h3;
  assign T_557 = 3'h5 == io_inner_acquire_bits_a_type;
  assign T_558 = T_557 ? 3'h1 : T_556;
  assign T_559 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T_560 = T_559 ? 3'h4 : T_558;
  assign T_561 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T_562 = T_561 ? 3'h3 : T_560;
  assign T_563 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T_564 = T_563 ? 3'h3 : T_562;
  assign T_565 = 3'h1 == io_inner_acquire_bits_a_type;
  assign T_566 = T_565 ? 3'h5 : T_564;
  assign T_567 = 3'h0 == io_inner_acquire_bits_a_type;
  assign T_568 = T_567 ? 3'h4 : T_566;
  assign GEN_248 = {{2'd0}, 1'h0};
  assign T_569 = io_inner_acquire_bits_a_type == GEN_248;
  assign T_574 = T_569 ? 2'h0 : 2'h1;
  assign T_575 = io_inner_acquire_bits_is_builtin_type ? T_568 : {{1'd0}, T_574};
  assign T_584_addr_beat = {{2'd0}, 1'h0};
  assign T_584_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign T_584_manager_xact_id = {{1'd0}, 2'h2};
  assign T_584_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign T_584_g_type = {{1'd0}, T_575};
  assign T_584_data = {{4'd0}, 1'h0};
  assign T_584_client_id = io_inner_acquire_bits_client_id;
  assign T_599_0 = 3'h5;
  assign T_599_1 = 3'h4;
  assign GEN_249 = {{1'd0}, T_599_0};
  assign T_601 = GEN_249 == T_584_g_type;
  assign GEN_250 = {{1'd0}, T_599_1};
  assign T_602 = GEN_250 == T_584_g_type;
  assign T_605 = T_601 | T_602;
  assign T_611_0 = 2'h0;
  assign T_611_1 = 2'h1;
  assign GEN_251 = {{2'd0}, T_611_0};
  assign T_613 = GEN_251 == T_584_g_type;
  assign GEN_252 = {{2'd0}, T_611_1};
  assign T_614 = GEN_252 == T_584_g_type;
  assign T_617 = T_613 | T_614;
  assign pending_outer_read_ = T_584_is_builtin_type ? T_605 : T_617;
  assign T_626_0 = 3'h2;
  assign T_626_1 = 3'h0;
  assign T_626_2 = 3'h4;
  assign T_628 = T_626_0 == xact_a_type;
  assign T_629 = T_626_1 == xact_a_type;
  assign T_630 = T_626_2 == xact_a_type;
  assign T_633 = T_628 | T_629;
  assign T_634 = T_633 | T_630;
  assign subblock_type = xact_is_builtin_type & T_634;
  assign T_636 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign T_637 = T_284 & T_636;
  assign T_639 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T_640 = T_284 & T_639;
  assign T_642 = io_inner_release_bits_voluntary == 1'h0;
  assign T_643 = T_640 & T_642;
  assign GEN_253 = $signed(8'hff);
  assign T_649 = $unsigned(GEN_253);
  assign T_674 = {T_649,1'h1};
  assign T_692 = 1'h1 ? {{3'd0}, T_674} : 12'h0;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign oacq_probe_client_xact_id = {{1'd0}, 2'h2};
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign oacq_probe_a_type = 3'h3;
  assign oacq_probe_union = T_692;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T_716 = xact_a_type == 3'h4;
  assign T_717 = xact_is_builtin_type & T_716;
  assign GEN_254 = {{7'd0}, 1'h1};
  assign T_721 = 8'h0 - GEN_254;
  assign T_722 = T_721[7:0];
  assign T_728_0 = T_722;
  assign T_731 = xact_a_type == 3'h3;
  assign T_732 = xact_is_builtin_type & T_731;
  assign T_734 = xact_a_type == 3'h2;
  assign T_735 = xact_is_builtin_type & T_734;
  assign T_736 = T_732 | T_735;
  assign T_737 = xact_union[8:1];
  assign T_739 = T_736 ? T_737 : {{7'd0}, 1'h0};
  assign T_740 = T_717 ? T_728_0 : T_739;
  assign T_767 = {T_740,1'h1};
  assign T_787 = 1'h1 ? {{3'd0}, T_767} : 12'h0;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_write_beat_client_xact_id = {{1'd0}, 2'h2};
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_write_beat_union = T_787;
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign GEN_0 = GEN_17;
  assign GEN_11 = GEN_234 == oacq_data_cnt ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign GEN_256 = {{1'd0}, 2'h2};
  assign GEN_12 = GEN_256 == oacq_data_cnt ? xact_wmask_buffer_2 : GEN_11;
  assign GEN_257 = {{1'd0}, 2'h3};
  assign GEN_13 = GEN_257 == oacq_data_cnt ? xact_wmask_buffer_3 : GEN_12;
  assign GEN_14 = 3'h4 == oacq_data_cnt ? xact_wmask_buffer_4 : GEN_13;
  assign GEN_15 = 3'h5 == oacq_data_cnt ? xact_wmask_buffer_5 : GEN_14;
  assign GEN_16 = 3'h6 == oacq_data_cnt ? xact_wmask_buffer_6 : GEN_15;
  assign GEN_17 = 3'h7 == oacq_data_cnt ? xact_wmask_buffer_7 : GEN_16;
  assign T_834 = {GEN_0,1'h1};
  assign T_852 = 1'h1 ? {{3'd0}, T_834} : 12'h0;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_block_client_xact_id = {{1'd0}, 2'h2};
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_block_union = T_852;
  assign oacq_write_block_data = GEN_1;
  assign GEN_1 = GEN_24;
  assign GEN_18 = GEN_234 == oacq_data_cnt ? xact_data_buffer_1 : xact_data_buffer_0;
  assign GEN_19 = GEN_256 == oacq_data_cnt ? xact_data_buffer_2 : GEN_18;
  assign GEN_20 = GEN_257 == oacq_data_cnt ? xact_data_buffer_3 : GEN_19;
  assign GEN_21 = 3'h4 == oacq_data_cnt ? xact_data_buffer_4 : GEN_20;
  assign GEN_22 = 3'h5 == oacq_data_cnt ? xact_data_buffer_5 : GEN_21;
  assign GEN_23 = 3'h6 == oacq_data_cnt ? xact_data_buffer_6 : GEN_22;
  assign GEN_24 = 3'h7 == oacq_data_cnt ? xact_data_buffer_7 : GEN_23;
  assign T_875 = xact_union[11:9];
  assign T_876 = xact_union[8:6];
  assign T_897 = {T_875,T_876};
  assign T_898 = {T_897,6'h0};
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign oacq_read_beat_client_xact_id = {{1'd0}, 2'h2};
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign oacq_read_beat_union = T_898;
  assign oacq_read_beat_data = {{4'd0}, 1'h0};
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_block_client_xact_id = {{1'd0}, 2'h2};
  assign oacq_read_block_addr_beat = {{2'd0}, 1'h0};
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_block_union = 12'h1c1;
  assign oacq_read_block_data = {{4'd0}, 1'h0};
  assign T_1013 = state == 3'h1;
  assign T_1014 = state == 3'h3;
  assign T_1015_addr_block = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign T_1015_client_xact_id = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign T_1015_addr_beat = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign T_1015_is_builtin_type = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign T_1015_a_type = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign T_1015_union = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign T_1015_data = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign T_1023_addr_block = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign T_1023_client_xact_id = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign T_1023_addr_beat = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign T_1023_is_builtin_type = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign T_1023_a_type = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign T_1023_union = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign T_1023_data = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign T_1031_addr_block = T_1014 ? T_1015_addr_block : T_1023_addr_block;
  assign T_1031_client_xact_id = T_1014 ? T_1015_client_xact_id : T_1023_client_xact_id;
  assign T_1031_addr_beat = T_1014 ? T_1015_addr_beat : T_1023_addr_beat;
  assign T_1031_is_builtin_type = T_1014 ? T_1015_is_builtin_type : T_1023_is_builtin_type;
  assign T_1031_a_type = T_1014 ? T_1015_a_type : T_1023_a_type;
  assign T_1031_union = T_1014 ? T_1015_union : T_1023_union;
  assign T_1031_data = T_1014 ? T_1015_data : T_1023_data;
  assign T_1039_addr_block = T_1013 ? oacq_probe_addr_block : T_1031_addr_block;
  assign T_1039_client_xact_id = T_1013 ? oacq_probe_client_xact_id : T_1031_client_xact_id;
  assign T_1039_addr_beat = T_1013 ? oacq_probe_addr_beat : T_1031_addr_beat;
  assign T_1039_is_builtin_type = T_1013 ? oacq_probe_is_builtin_type : T_1031_is_builtin_type;
  assign T_1039_a_type = T_1013 ? oacq_probe_a_type : T_1031_a_type;
  assign T_1039_union = T_1013 ? oacq_probe_union : T_1031_union;
  assign T_1039_data = T_1013 ? oacq_probe_data : T_1031_data;
  assign T_1056 = 3'h4 == xact_a_type;
  assign T_1057 = T_1056 ? 2'h0 : 2'h2;
  assign T_1058 = 3'h6 == xact_a_type;
  assign T_1059 = T_1058 ? 2'h0 : T_1057;
  assign T_1060 = 3'h5 == xact_a_type;
  assign T_1061 = T_1060 ? 2'h2 : T_1059;
  assign T_1062 = 3'h2 == xact_a_type;
  assign T_1063 = T_1062 ? 2'h0 : T_1061;
  assign T_1064 = 3'h0 == xact_a_type;
  assign T_1065 = T_1064 ? 2'h2 : T_1063;
  assign T_1066 = 3'h3 == xact_a_type;
  assign T_1067 = T_1066 ? 2'h0 : T_1065;
  assign T_1068 = 3'h1 == xact_a_type;
  assign T_1069 = T_1068 ? 2'h2 : T_1067;
  assign T_1070 = GEN_234 == xact_a_type;
  assign T_1071 = T_1070 ? 2'h0 : 2'h2;
  assign T_1072 = GEN_248 == xact_a_type;
  assign T_1073 = T_1072 ? 2'h1 : T_1071;
  assign T_1074 = xact_is_builtin_type ? T_1069 : T_1073;
  assign T_1079_addr_block = xact_addr_block;
  assign T_1079_p_type = T_1074;
  assign T_1079_client_id = {{1'd0}, 1'h0};
  assign T_1103 = T_1058 ? 3'h1 : 3'h3;
  assign T_1105 = T_1060 ? 3'h1 : T_1103;
  assign T_1107 = T_1056 ? 3'h4 : T_1105;
  assign T_1109 = T_1066 ? 3'h3 : T_1107;
  assign T_1111 = T_1062 ? 3'h3 : T_1109;
  assign T_1113 = T_1068 ? 3'h5 : T_1111;
  assign T_1115 = T_1064 ? 3'h4 : T_1113;
  assign T_1116 = xact_a_type == GEN_248;
  assign T_1121 = T_1116 ? 2'h0 : 2'h1;
  assign T_1122 = xact_is_builtin_type ? T_1115 : {{1'd0}, T_1121};
  assign T_1131_addr_beat = {{2'd0}, 1'h0};
  assign T_1131_client_xact_id = xact_client_xact_id;
  assign T_1131_manager_xact_id = {{1'd0}, 2'h2};
  assign T_1131_is_builtin_type = xact_is_builtin_type;
  assign T_1131_g_type = {{1'd0}, T_1122};
  assign T_1131_data = {{4'd0}, 1'h0};
  assign T_1131_client_id = xact_client_id;
  assign T_1143 = T_284 & collect_iacq_data;
  assign T_1145 = T_1143 & T_324;
  assign T_1146 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T_1147 = T_1145 & T_1146;
  assign T_1149 = T_1147 == 1'h0;
  assign T_1150 = T_1149 | reset;
  assign T_1152 = T_1150 == 1'h0;
  assign T_1157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T_1158 = T_1145 & T_1157;
  assign T_1160 = T_1158 == 1'h0;
  assign T_1161 = T_1160 | reset;
  assign T_1163 = T_1161 == 1'h0;
  assign T_1164 = state == 3'h0;
  assign T_1166 = T_1164 & T_324;
  assign T_1167 = T_1166 & io_alloc_iacq;
  assign T_1176_0 = 3'h3;
  assign T_1178 = T_1176_0 == io_inner_acquire_bits_a_type;
  assign T_1181 = io_inner_acquire_bits_is_builtin_type & T_1178;
  assign T_1182 = T_1167 & T_1181;
  assign T_1184 = io_inner_acquire_bits_addr_beat != GEN_248;
  assign T_1185 = T_1182 & T_1184;
  assign T_1187 = T_1185 == 1'h0;
  assign T_1188 = T_1187 | reset;
  assign T_1190 = T_1188 == 1'h0;
  assign GEN_2 = io_inner_acquire_bits_data;
  assign GEN_25 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_0;
  assign GEN_26 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_1;
  assign GEN_27 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_2;
  assign GEN_28 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_3;
  assign GEN_29 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_4;
  assign GEN_30 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_5;
  assign GEN_31 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_6;
  assign GEN_32 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_7;
  assign T_1193 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_1194 = io_inner_acquire_bits_is_builtin_type & T_1193;
  assign T_1205_0 = T_722;
  assign T_1208 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1209 = io_inner_acquire_bits_is_builtin_type & T_1208;
  assign T_1211 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1212 = io_inner_acquire_bits_is_builtin_type & T_1211;
  assign T_1213 = T_1209 | T_1212;
  assign T_1214 = io_inner_acquire_bits_union[8:1];
  assign T_1216 = T_1213 ? T_1214 : {{7'd0}, 1'h0};
  assign T_1217 = T_1194 ? T_1205_0 : T_1216;
  assign GEN_3 = T_1217;
  assign GEN_33 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_0;
  assign GEN_34 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_1;
  assign GEN_35 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_2;
  assign GEN_36 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_3;
  assign GEN_37 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_4;
  assign GEN_38 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_5;
  assign GEN_39 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_6;
  assign GEN_40 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_7;
  assign T_1220 = GEN_254 << io_inner_acquire_bits_addr_beat;
  assign T_1221 = iacq_data_valid | T_1220;
  assign GEN_42 = io_inner_acquire_valid ? GEN_25 : xact_data_buffer_0;
  assign GEN_43 = io_inner_acquire_valid ? GEN_26 : xact_data_buffer_1;
  assign GEN_44 = io_inner_acquire_valid ? GEN_27 : xact_data_buffer_2;
  assign GEN_45 = io_inner_acquire_valid ? GEN_28 : xact_data_buffer_3;
  assign GEN_46 = io_inner_acquire_valid ? GEN_29 : xact_data_buffer_4;
  assign GEN_47 = io_inner_acquire_valid ? GEN_30 : xact_data_buffer_5;
  assign GEN_48 = io_inner_acquire_valid ? GEN_31 : xact_data_buffer_6;
  assign GEN_49 = io_inner_acquire_valid ? GEN_32 : xact_data_buffer_7;
  assign GEN_52 = io_inner_acquire_valid ? GEN_33 : xact_wmask_buffer_0;
  assign GEN_53 = io_inner_acquire_valid ? GEN_34 : xact_wmask_buffer_1;
  assign GEN_54 = io_inner_acquire_valid ? GEN_35 : xact_wmask_buffer_2;
  assign GEN_55 = io_inner_acquire_valid ? GEN_36 : xact_wmask_buffer_3;
  assign GEN_56 = io_inner_acquire_valid ? GEN_37 : xact_wmask_buffer_4;
  assign GEN_57 = io_inner_acquire_valid ? GEN_38 : xact_wmask_buffer_5;
  assign GEN_58 = io_inner_acquire_valid ? GEN_39 : xact_wmask_buffer_6;
  assign GEN_59 = io_inner_acquire_valid ? GEN_40 : xact_wmask_buffer_7;
  assign GEN_60 = io_inner_acquire_valid ? T_1221 : iacq_data_valid;
  assign GEN_61 = iacq_data_done ? 1'h0 : collect_iacq_data;
  assign GEN_64 = collect_iacq_data ? GEN_42 : xact_data_buffer_0;
  assign GEN_65 = collect_iacq_data ? GEN_43 : xact_data_buffer_1;
  assign GEN_66 = collect_iacq_data ? GEN_44 : xact_data_buffer_2;
  assign GEN_67 = collect_iacq_data ? GEN_45 : xact_data_buffer_3;
  assign GEN_68 = collect_iacq_data ? GEN_46 : xact_data_buffer_4;
  assign GEN_69 = collect_iacq_data ? GEN_47 : xact_data_buffer_5;
  assign GEN_70 = collect_iacq_data ? GEN_48 : xact_data_buffer_6;
  assign GEN_71 = collect_iacq_data ? GEN_49 : xact_data_buffer_7;
  assign GEN_74 = collect_iacq_data ? GEN_52 : xact_wmask_buffer_0;
  assign GEN_75 = collect_iacq_data ? GEN_53 : xact_wmask_buffer_1;
  assign GEN_76 = collect_iacq_data ? GEN_54 : xact_wmask_buffer_2;
  assign GEN_77 = collect_iacq_data ? GEN_55 : xact_wmask_buffer_3;
  assign GEN_78 = collect_iacq_data ? GEN_56 : xact_wmask_buffer_4;
  assign GEN_79 = collect_iacq_data ? GEN_57 : xact_wmask_buffer_5;
  assign GEN_80 = collect_iacq_data ? GEN_58 : xact_wmask_buffer_6;
  assign GEN_81 = collect_iacq_data ? GEN_59 : xact_wmask_buffer_7;
  assign GEN_82 = collect_iacq_data ? GEN_60 : iacq_data_valid;
  assign GEN_83 = collect_iacq_data ? GEN_61 : collect_iacq_data;
  assign GEN_84 = io_outer_grant_valid ? 1'h0 : pending_ognt_ack;
  assign GEN_86 = pending_ognt_ack ? GEN_84 : pending_ognt_ack;
  assign T_1229 = 3'h0 == state;
  assign T_1231 = io_inner_acquire_valid & io_alloc_iacq;
  assign GEN_4 = io_inner_acquire_bits_data;
  assign T_1247_0 = T_722;
  assign T_1259 = T_1194 ? T_1247_0 : T_1216;
  assign GEN_5 = T_1259;
  assign T_1268_0 = 3'h3;
  assign T_1270 = T_1268_0 == io_inner_acquire_bits_a_type;
  assign T_1273 = io_inner_acquire_bits_is_builtin_type & T_1270;
  assign T_1282_0 = 3'h2;
  assign T_1282_1 = 3'h3;
  assign T_1282_2 = 3'h4;
  assign T_1284 = T_1282_0 == io_inner_acquire_bits_a_type;
  assign T_1285 = T_1282_1 == io_inner_acquire_bits_a_type;
  assign T_1286 = T_1282_2 == io_inner_acquire_bits_a_type;
  assign T_1289 = T_1284 | T_1285;
  assign T_1290 = T_1289 | T_1286;
  assign T_1291 = io_inner_acquire_bits_is_builtin_type & T_1290;
  assign GEN_276 = {{7'd0}, T_1291};
  assign T_1292 = GEN_276 << io_inner_acquire_bits_addr_beat;
  assign GEN_277 = {{3'd0}, 1'h0};
  assign T_1294 = mask_incoherent != GEN_277;
  assign T_1295 = mask_incoherent[0];
  assign T_1296 = mask_incoherent[1];
  assign T_1297 = mask_incoherent[2];
  assign T_1298 = mask_incoherent[3];
  assign T_1300 = {1'h0,T_1296};
  assign GEN_278 = {{1'd0}, T_1295};
  assign T_1301 = GEN_278 + T_1300;
  assign T_1302 = T_1301[1:0];
  assign T_1305 = {1'h0,T_1298};
  assign GEN_279 = {{1'd0}, T_1297};
  assign T_1306 = GEN_279 + T_1305;
  assign T_1307 = T_1306[1:0];
  assign T_1308 = {1'h0,T_1307};
  assign GEN_280 = {{1'd0}, T_1302};
  assign T_1309 = GEN_280 + T_1308;
  assign T_1310 = T_1309[2:0];
  assign GEN_103 = T_1294 ? mask_incoherent : {{3'd0}, pending_probes};
  assign GEN_104 = T_1294 ? T_1310 : {{2'd0}, release_count};
  assign T_1311 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign T_1312 = pending_outer_write_ ? 3'h3 : T_1311;
  assign T_1313 = T_1294 ? 3'h1 : T_1312;
  assign GEN_105 = T_1231 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_106 = T_1231 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign GEN_107 = T_1231 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign GEN_108 = T_1231 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign GEN_109 = T_1231 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign GEN_110 = T_1231 ? io_inner_acquire_bits_union : xact_union;
  assign GEN_111 = T_1231 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign GEN_113 = T_1231 ? GEN_4 : GEN_64;
  assign GEN_123 = T_1231 ? GEN_5 : GEN_74;
  assign GEN_132 = T_1231 ? T_1273 : GEN_83;
  assign GEN_136 = T_1231 ? T_1292 : GEN_82;
  assign GEN_137 = T_1231 ? GEN_103 : {{3'd0}, pending_probes};
  assign GEN_138 = T_1231 ? GEN_104 : {{2'd0}, release_count};
  assign GEN_139 = T_1231 ? T_1313 : state;
  assign GEN_140 = T_1229 ? 1'h1 : collect_iacq_data;
  assign GEN_141 = T_1229 ? GEN_105 : xact_addr_block;
  assign GEN_142 = T_1229 ? GEN_106 : xact_client_xact_id;
  assign GEN_143 = T_1229 ? GEN_107 : xact_addr_beat;
  assign GEN_144 = T_1229 ? GEN_108 : xact_is_builtin_type;
  assign GEN_145 = T_1229 ? GEN_109 : xact_a_type;
  assign GEN_146 = T_1229 ? GEN_110 : xact_union;
  assign GEN_147 = T_1229 ? GEN_111 : xact_client_id;
  assign GEN_149 = T_1229 ? GEN_113 : GEN_64;
  assign GEN_159 = T_1229 ? GEN_123 : GEN_74;
  assign GEN_168 = T_1229 ? GEN_132 : GEN_83;
  assign GEN_172 = T_1229 ? GEN_136 : GEN_82;
  assign GEN_173 = T_1229 ? GEN_137 : {{3'd0}, pending_probes};
  assign GEN_174 = T_1229 ? GEN_138 : {{2'd0}, release_count};
  assign GEN_175 = T_1229 ? GEN_139 : state;
  assign T_1314 = 3'h1 == state;
  assign GEN_281 = {{1'd0}, 1'h1};
  assign T_1318 = GEN_281 << 1'h0;
  assign T_1319 = ~ T_1318;
  assign GEN_282 = {{1'd0}, pending_probes};
  assign T_1320 = GEN_282 & T_1319;
  assign GEN_176 = io_inner_probe_ready ? {{2'd0}, T_1320} : GEN_173;
  assign T_1326_0 = 3'h0;
  assign T_1326_1 = 3'h1;
  assign T_1326_2 = 3'h2;
  assign T_1328 = T_1326_0 == io_inner_release_bits_r_type;
  assign T_1329 = T_1326_1 == io_inner_release_bits_r_type;
  assign T_1330 = T_1326_2 == io_inner_release_bits_r_type;
  assign T_1333 = T_1328 | T_1329;
  assign T_1334 = T_1333 | T_1330;
  assign T_1336 = T_1334 == 1'h0;
  assign T_1337 = T_1336 | io_outer_acquire_ready;
  assign T_1338 = T_1337 & io_matches_irel;
  assign T_1339 = io_inner_release_valid & io_matches_irel;
  assign T_1345_0 = 3'h0;
  assign T_1345_1 = 3'h1;
  assign T_1345_2 = 3'h2;
  assign T_1347 = T_1345_0 == io_inner_release_bits_r_type;
  assign T_1348 = T_1345_1 == io_inner_release_bits_r_type;
  assign T_1349 = T_1345_2 == io_inner_release_bits_r_type;
  assign T_1352 = T_1347 | T_1348;
  assign T_1353 = T_1352 | T_1349;
  assign T_1357 = release_count - 1'h1;
  assign T_1358 = T_1357[0:0];
  assign T_1361 = pending_outer_read ? 3'h2 : 3'h4;
  assign T_1362 = pending_outer_write ? 3'h3 : T_1361;
  assign GEN_177 = release_count ? T_1362 : GEN_175;
  assign GEN_178 = oacq_data_done ? 1'h1 : GEN_86;
  assign GEN_179 = oacq_data_done ? {{2'd0}, T_1358} : GEN_174;
  assign GEN_180 = oacq_data_done ? GEN_177 : GEN_175;
  assign GEN_181 = io_outer_acquire_ready ? GEN_178 : GEN_86;
  assign GEN_182 = io_outer_acquire_ready ? GEN_179 : GEN_174;
  assign GEN_183 = io_outer_acquire_ready ? GEN_180 : GEN_175;
  assign GEN_185 = T_1353 ? GEN_181 : GEN_86;
  assign GEN_186 = T_1353 ? GEN_182 : GEN_174;
  assign GEN_187 = T_1353 ? GEN_183 : GEN_175;
  assign T_1364 = T_1353 == 1'h0;
  assign GEN_188 = release_count ? T_1362 : GEN_187;
  assign GEN_189 = T_1364 ? {{2'd0}, T_1358} : GEN_186;
  assign GEN_190 = T_1364 ? GEN_188 : GEN_187;
  assign GEN_194 = T_1339 ? T_1353 : 1'h0;
  assign GEN_195 = T_1339 ? GEN_185 : GEN_86;
  assign GEN_196 = T_1339 ? GEN_189 : GEN_174;
  assign GEN_197 = T_1339 ? GEN_190 : GEN_175;
  assign GEN_198 = T_1314 ? pending_probes : 1'h0;
  assign GEN_199 = T_1314 ? GEN_176 : GEN_173;
  assign GEN_203 = T_1314 ? T_1338 : 1'h0;
  assign GEN_207 = T_1314 ? GEN_194 : 1'h0;
  assign GEN_208 = T_1314 ? GEN_195 : GEN_86;
  assign GEN_209 = T_1314 ? GEN_196 : GEN_174;
  assign GEN_210 = T_1314 ? GEN_197 : GEN_175;
  assign T_1372 = 3'h3 == state;
  assign T_1374 = pending_ognt_ack == 1'h0;
  assign T_1376 = collect_iacq_data == 1'h0;
  assign T_1377 = iacq_data_valid >> oacq_data_cnt;
  assign T_1378 = T_1377[0];
  assign T_1379 = T_1376 | T_1378;
  assign T_1380 = T_1374 & T_1379;
  assign T_1382 = pending_outer_read ? 3'h2 : 3'h5;
  assign GEN_211 = oacq_data_done ? 1'h1 : GEN_208;
  assign GEN_212 = oacq_data_done ? T_1382 : GEN_210;
  assign GEN_213 = T_1372 ? T_1380 : GEN_207;
  assign GEN_214 = T_1372 ? GEN_211 : GEN_208;
  assign GEN_215 = T_1372 ? GEN_212 : GEN_210;
  assign T_1383 = 3'h2 == state;
  assign GEN_216 = T_416 ? 3'h5 : GEN_215;
  assign GEN_217 = T_1383 ? T_1374 : GEN_213;
  assign GEN_218 = T_1383 ? GEN_216 : GEN_215;
  assign T_1387 = 3'h5 == state;
  assign GEN_283 = {{1'd0}, 3'h0};
  assign T_1392 = io_inner_grant_bits_g_type == GEN_283;
  assign T_1393 = io_inner_grant_bits_is_builtin_type & T_1392;
  assign T_1395 = T_1393 == 1'h0;
  assign T_1397 = T_1395 ? 3'h6 : 3'h0;
  assign GEN_219 = ignt_data_done ? T_1397 : GEN_218;
  assign GEN_220 = T_1387 ? io_inner_grant_ready : pending_ognt_ack;
  assign GEN_221 = T_1387 ? io_outer_grant_valid : 1'h0;
  assign GEN_222 = T_1387 ? GEN_219 : GEN_218;
  assign T_1398 = 3'h4 == state;
  assign GEN_223 = io_inner_grant_ready ? T_1397 : GEN_222;
  assign GEN_224 = T_1398 ? 1'h1 : GEN_221;
  assign GEN_225 = T_1398 ? GEN_223 : GEN_222;
  assign T_1410 = 3'h6 == state;
  assign GEN_226 = io_inner_finish_valid ? 3'h0 : GEN_225;
  assign GEN_228 = T_1410 ? GEN_226 : GEN_225;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_41 = {1{$random}};
  state = GEN_41[2:0];
  GEN_50 = {1{$random}};
  xact_addr_block = GEN_50[25:0];
  GEN_51 = {1{$random}};
  xact_client_xact_id = GEN_51[1:0];
  GEN_62 = {1{$random}};
  xact_addr_beat = GEN_62[2:0];
  GEN_63 = {1{$random}};
  xact_is_builtin_type = GEN_63[0:0];
  GEN_72 = {1{$random}};
  xact_a_type = GEN_72[2:0];
  GEN_73 = {1{$random}};
  xact_union = GEN_73[11:0];
  GEN_85 = {1{$random}};
  xact_data_buffer_0 = GEN_85[4:0];
  GEN_87 = {1{$random}};
  xact_data_buffer_1 = GEN_87[4:0];
  GEN_88 = {1{$random}};
  xact_data_buffer_2 = GEN_88[4:0];
  GEN_89 = {1{$random}};
  xact_data_buffer_3 = GEN_89[4:0];
  GEN_90 = {1{$random}};
  xact_data_buffer_4 = GEN_90[4:0];
  GEN_91 = {1{$random}};
  xact_data_buffer_5 = GEN_91[4:0];
  GEN_92 = {1{$random}};
  xact_data_buffer_6 = GEN_92[4:0];
  GEN_93 = {1{$random}};
  xact_data_buffer_7 = GEN_93[4:0];
  GEN_94 = {1{$random}};
  xact_wmask_buffer_0 = GEN_94[7:0];
  GEN_95 = {1{$random}};
  xact_wmask_buffer_1 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  xact_wmask_buffer_2 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  xact_wmask_buffer_3 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  xact_wmask_buffer_4 = GEN_98[7:0];
  GEN_99 = {1{$random}};
  xact_wmask_buffer_5 = GEN_99[7:0];
  GEN_100 = {1{$random}};
  xact_wmask_buffer_6 = GEN_100[7:0];
  GEN_101 = {1{$random}};
  xact_wmask_buffer_7 = GEN_101[7:0];
  GEN_102 = {1{$random}};
  xact_client_id = GEN_102[1:0];
  GEN_112 = {1{$random}};
  release_count = GEN_112[0:0];
  GEN_114 = {1{$random}};
  pending_probes = GEN_114[0:0];
  GEN_115 = {1{$random}};
  collect_iacq_data = GEN_115[0:0];
  GEN_116 = {1{$random}};
  iacq_data_valid = GEN_116[7:0];
  GEN_117 = {1{$random}};
  T_342 = GEN_117[2:0];
  GEN_118 = {1{$random}};
  T_370 = GEN_118[2:0];
  GEN_119 = {1{$random}};
  T_408 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  T_433 = GEN_120[2:0];
  GEN_121 = {1{$random}};
  T_468 = GEN_121[2:0];
  GEN_122 = {1{$random}};
  pending_ognt_ack = GEN_122[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_228;
    end
    if(1'h0) begin
    end else begin
      xact_addr_block <= GEN_141;
    end
    if(1'h0) begin
    end else begin
      xact_client_xact_id <= GEN_142;
    end
    if(1'h0) begin
    end else begin
      xact_addr_beat <= GEN_143;
    end
    if(1'h0) begin
    end else begin
      xact_is_builtin_type <= GEN_144;
    end
    if(1'h0) begin
    end else begin
      xact_a_type <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      xact_union <= GEN_146;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_0 <= GEN_149;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_1 <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_2 <= GEN_66;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_3 <= GEN_67;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_4 <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_5 <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_6 <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_7 <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_0 <= GEN_159;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_1 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_2 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_3 <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_4 <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_5 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_6 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_7 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      xact_client_id <= GEN_147;
    end
    if(reset) begin
      release_count <= 1'h0;
    end else begin
      release_count <= GEN_209[0];
    end
    if(reset) begin
      pending_probes <= 1'h0;
    end else begin
      pending_probes <= GEN_199[0];
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else begin
      collect_iacq_data <= GEN_168;
    end
    if(reset) begin
      iacq_data_valid <= 8'h0;
    end else begin
      iacq_data_valid <= GEN_172;
    end
    if(reset) begin
      T_342 <= 3'h0;
    end else begin
      T_342 <= GEN_6;
    end
    if(reset) begin
      T_370 <= 3'h0;
    end else begin
      T_370 <= GEN_7;
    end
    if(reset) begin
      T_408 <= 3'h0;
    end else begin
      T_408 <= GEN_8;
    end
    if(reset) begin
      T_433 <= 3'h0;
    end else begin
      T_433 <= GEN_9;
    end
    if(reset) begin
      T_468 <= 3'h0;
    end else begin
      T_468 <= GEN_10;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else begin
      pending_ognt_ack <= GEN_214;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics or prefetches\n    at broadcast.scala:203 assert(!(state =/= s_idle && xact.isBuiltInType() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different network source than initial request.\n    at broadcast.scala:285 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different client transaction than initial request.\n    at broadcast.scala:289 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at broadcast.scala:293 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module BroadcastAcquireTracker_29(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [4:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [4:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [4:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [4:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [4:0] io_outer_grant_bits_data,
  output  io_matches_iacq,
  output  io_matches_irel,
  output  io_matches_oprb,
  input   io_alloc_iacq,
  input   io_alloc_irel,
  input   io_alloc_oprb
);
  reg [2:0] state;
  reg [31:0] GEN_41;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_50;
  reg [1:0] xact_client_xact_id;
  reg [31:0] GEN_51;
  reg [2:0] xact_addr_beat;
  reg [31:0] GEN_62;
  reg  xact_is_builtin_type;
  reg [31:0] GEN_63;
  reg [2:0] xact_a_type;
  reg [31:0] GEN_72;
  reg [11:0] xact_union;
  reg [31:0] GEN_73;
  reg [4:0] xact_data_buffer_0;
  reg [31:0] GEN_85;
  reg [4:0] xact_data_buffer_1;
  reg [31:0] GEN_87;
  reg [4:0] xact_data_buffer_2;
  reg [31:0] GEN_88;
  reg [4:0] xact_data_buffer_3;
  reg [31:0] GEN_89;
  reg [4:0] xact_data_buffer_4;
  reg [31:0] GEN_90;
  reg [4:0] xact_data_buffer_5;
  reg [31:0] GEN_91;
  reg [4:0] xact_data_buffer_6;
  reg [31:0] GEN_92;
  reg [4:0] xact_data_buffer_7;
  reg [31:0] GEN_93;
  reg [7:0] xact_wmask_buffer_0;
  reg [31:0] GEN_94;
  reg [7:0] xact_wmask_buffer_1;
  reg [31:0] GEN_95;
  reg [7:0] xact_wmask_buffer_2;
  reg [31:0] GEN_96;
  reg [7:0] xact_wmask_buffer_3;
  reg [31:0] GEN_97;
  reg [7:0] xact_wmask_buffer_4;
  reg [31:0] GEN_98;
  reg [7:0] xact_wmask_buffer_5;
  reg [31:0] GEN_99;
  reg [7:0] xact_wmask_buffer_6;
  reg [31:0] GEN_100;
  reg [7:0] xact_wmask_buffer_7;
  reg [31:0] GEN_101;
  reg [1:0] xact_client_id;
  reg [31:0] GEN_102;
  wire  coh_sharers;
  wire  T_284;
  wire  T_285;
  wire [2:0] T_294_0;
  wire [2:0] T_294_1;
  wire [2:0] T_294_2;
  wire  T_296;
  wire  T_297;
  wire  T_298;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_305;
  wire  T_306;
  wire  T_308;
  reg  release_count;
  reg [31:0] GEN_112;
  reg  pending_probes;
  reg [31:0] GEN_114;
  wire  GEN_229;
  wire  T_313;
  wire [3:0] GEN_230;
  wire [3:0] T_316;
  wire  T_318;
  wire [3:0] GEN_232;
  wire [3:0] T_319;
  wire [3:0] T_320;
  wire  T_321;
  wire [3:0] GEN_233;
  wire [3:0] mask_incoherent;
  reg  collect_iacq_data;
  reg [31:0] GEN_115;
  reg [7:0] iacq_data_valid;
  reg [31:0] GEN_116;
  wire  T_324;
  wire [2:0] T_334_0;
  wire  T_336;
  wire  T_339;
  wire  T_340;
  reg [2:0] T_342;
  reg [31:0] GEN_117;
  wire  T_344;
  wire [2:0] GEN_234;
  wire [3:0] T_346;
  wire [2:0] T_347;
  wire [2:0] GEN_6;
  wire  T_348;
  wire  iacq_data_done;
  wire  T_350;
  wire [2:0] T_358_0;
  wire [2:0] T_358_1;
  wire [2:0] T_358_2;
  wire  T_360;
  wire  T_361;
  wire  T_362;
  wire  T_365;
  wire  T_366;
  wire  T_368;
  reg [2:0] T_370;
  reg [31:0] GEN_118;
  wire [3:0] T_374;
  wire [2:0] T_375;
  wire [2:0] GEN_7;
  wire  T_379;
  wire [2:0] T_387_0;
  wire [3:0] GEN_236;
  wire  T_389;
  wire [1:0] T_397_0;
  wire [1:0] T_397_1;
  wire [3:0] GEN_237;
  wire  T_399;
  wire [3:0] GEN_238;
  wire  T_400;
  wire  T_403;
  wire  T_404;
  wire  T_406;
  reg [2:0] T_408;
  reg [31:0] GEN_119;
  wire  T_410;
  wire [3:0] T_412;
  wire [2:0] T_413;
  wire [2:0] GEN_8;
  wire  T_414;
  wire  ignt_data_done;
  wire  T_416;
  wire [2:0] T_425_0;
  wire  T_427;
  wire  T_430;
  wire  T_431;
  reg [2:0] T_433;
  reg [31:0] GEN_120;
  wire  T_435;
  wire [3:0] T_437;
  wire [2:0] T_438;
  wire [2:0] GEN_9;
  wire  T_439;
  wire [2:0] oacq_data_cnt;
  wire  oacq_data_done;
  wire  T_440;
  wire [2:0] T_449_0;
  wire [3:0] GEN_241;
  wire  T_451;
  wire  T_459_0;
  wire [3:0] GEN_242;
  wire  T_461;
  wire  T_464;
  wire  T_466;
  reg [2:0] T_468;
  reg [31:0] GEN_121;
  wire [3:0] T_472;
  wire [2:0] T_473;
  wire [2:0] GEN_10;
  reg  pending_ognt_ack;
  reg [31:0] GEN_122;
  wire [2:0] T_485_0;
  wire [2:0] T_485_1;
  wire [2:0] T_485_2;
  wire  T_487;
  wire  T_488;
  wire  T_489;
  wire  T_492;
  wire  T_493;
  wire  pending_outer_write;
  wire [2:0] T_502_0;
  wire [2:0] T_502_1;
  wire [2:0] T_502_2;
  wire  T_504;
  wire  T_505;
  wire  T_506;
  wire  T_509;
  wire  T_510;
  wire  pending_outer_write_;
  wire [2:0] T_518_0;
  wire [2:0] T_518_1;
  wire [3:0] GEN_244;
  wire  T_520;
  wire [3:0] GEN_245;
  wire  T_521;
  wire  T_524;
  wire [1:0] T_530_0;
  wire [1:0] T_530_1;
  wire [3:0] GEN_246;
  wire  T_532;
  wire [3:0] GEN_247;
  wire  T_533;
  wire  T_536;
  wire  pending_outer_read;
  wire  T_555;
  wire [2:0] T_556;
  wire  T_557;
  wire [2:0] T_558;
  wire  T_559;
  wire [2:0] T_560;
  wire  T_561;
  wire [2:0] T_562;
  wire  T_563;
  wire [2:0] T_564;
  wire  T_565;
  wire [2:0] T_566;
  wire  T_567;
  wire [2:0] T_568;
  wire [2:0] GEN_248;
  wire  T_569;
  wire [1:0] T_574;
  wire [2:0] T_575;
  wire [2:0] T_584_addr_beat;
  wire [1:0] T_584_client_xact_id;
  wire [2:0] T_584_manager_xact_id;
  wire  T_584_is_builtin_type;
  wire [3:0] T_584_g_type;
  wire [4:0] T_584_data;
  wire [1:0] T_584_client_id;
  wire [2:0] T_599_0;
  wire [2:0] T_599_1;
  wire [3:0] GEN_249;
  wire  T_601;
  wire [3:0] GEN_250;
  wire  T_602;
  wire  T_605;
  wire [1:0] T_611_0;
  wire [1:0] T_611_1;
  wire [3:0] GEN_251;
  wire  T_613;
  wire [3:0] GEN_252;
  wire  T_614;
  wire  T_617;
  wire  pending_outer_read_;
  wire [2:0] T_626_0;
  wire [2:0] T_626_1;
  wire [2:0] T_626_2;
  wire  T_628;
  wire  T_629;
  wire  T_630;
  wire  T_633;
  wire  T_634;
  wire  subblock_type;
  wire  T_636;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire  T_642;
  wire  T_643;
  wire [7:0] GEN_253;
  wire [7:0] T_649;
  wire [8:0] T_674;
  wire [11:0] T_692;
  wire [25:0] oacq_probe_addr_block;
  wire [2:0] oacq_probe_client_xact_id;
  wire [2:0] oacq_probe_addr_beat;
  wire  oacq_probe_is_builtin_type;
  wire [2:0] oacq_probe_a_type;
  wire [11:0] oacq_probe_union;
  wire [4:0] oacq_probe_data;
  wire  T_716;
  wire  T_717;
  wire [7:0] GEN_254;
  wire [8:0] T_721;
  wire [7:0] T_722;
  wire [7:0] T_728_0;
  wire  T_731;
  wire  T_732;
  wire  T_734;
  wire  T_735;
  wire  T_736;
  wire [7:0] T_737;
  wire [7:0] T_739;
  wire [7:0] T_740;
  wire [8:0] T_767;
  wire [11:0] T_787;
  wire [25:0] oacq_write_beat_addr_block;
  wire [2:0] oacq_write_beat_client_xact_id;
  wire [2:0] oacq_write_beat_addr_beat;
  wire  oacq_write_beat_is_builtin_type;
  wire [2:0] oacq_write_beat_a_type;
  wire [11:0] oacq_write_beat_union;
  wire [4:0] oacq_write_beat_data;
  wire [7:0] GEN_0;
  wire [7:0] GEN_11;
  wire [2:0] GEN_256;
  wire [7:0] GEN_12;
  wire [2:0] GEN_257;
  wire [7:0] GEN_13;
  wire [7:0] GEN_14;
  wire [7:0] GEN_15;
  wire [7:0] GEN_16;
  wire [7:0] GEN_17;
  wire [8:0] T_834;
  wire [11:0] T_852;
  wire [25:0] oacq_write_block_addr_block;
  wire [2:0] oacq_write_block_client_xact_id;
  wire [2:0] oacq_write_block_addr_beat;
  wire  oacq_write_block_is_builtin_type;
  wire [2:0] oacq_write_block_a_type;
  wire [11:0] oacq_write_block_union;
  wire [4:0] oacq_write_block_data;
  wire [4:0] GEN_1;
  wire [4:0] GEN_18;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [2:0] T_875;
  wire [2:0] T_876;
  wire [5:0] T_897;
  wire [11:0] T_898;
  wire [25:0] oacq_read_beat_addr_block;
  wire [2:0] oacq_read_beat_client_xact_id;
  wire [2:0] oacq_read_beat_addr_beat;
  wire  oacq_read_beat_is_builtin_type;
  wire [2:0] oacq_read_beat_a_type;
  wire [11:0] oacq_read_beat_union;
  wire [4:0] oacq_read_beat_data;
  wire [25:0] oacq_read_block_addr_block;
  wire [2:0] oacq_read_block_client_xact_id;
  wire [2:0] oacq_read_block_addr_beat;
  wire  oacq_read_block_is_builtin_type;
  wire [2:0] oacq_read_block_a_type;
  wire [11:0] oacq_read_block_union;
  wire [4:0] oacq_read_block_data;
  wire  T_1013;
  wire  T_1014;
  wire [25:0] T_1015_addr_block;
  wire [2:0] T_1015_client_xact_id;
  wire [2:0] T_1015_addr_beat;
  wire  T_1015_is_builtin_type;
  wire [2:0] T_1015_a_type;
  wire [11:0] T_1015_union;
  wire [4:0] T_1015_data;
  wire [25:0] T_1023_addr_block;
  wire [2:0] T_1023_client_xact_id;
  wire [2:0] T_1023_addr_beat;
  wire  T_1023_is_builtin_type;
  wire [2:0] T_1023_a_type;
  wire [11:0] T_1023_union;
  wire [4:0] T_1023_data;
  wire [25:0] T_1031_addr_block;
  wire [2:0] T_1031_client_xact_id;
  wire [2:0] T_1031_addr_beat;
  wire  T_1031_is_builtin_type;
  wire [2:0] T_1031_a_type;
  wire [11:0] T_1031_union;
  wire [4:0] T_1031_data;
  wire [25:0] T_1039_addr_block;
  wire [2:0] T_1039_client_xact_id;
  wire [2:0] T_1039_addr_beat;
  wire  T_1039_is_builtin_type;
  wire [2:0] T_1039_a_type;
  wire [11:0] T_1039_union;
  wire [4:0] T_1039_data;
  wire  T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire  T_1060;
  wire [1:0] T_1061;
  wire  T_1062;
  wire [1:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire  T_1066;
  wire [1:0] T_1067;
  wire  T_1068;
  wire [1:0] T_1069;
  wire  T_1070;
  wire [1:0] T_1071;
  wire  T_1072;
  wire [1:0] T_1073;
  wire [1:0] T_1074;
  wire [25:0] T_1079_addr_block;
  wire [1:0] T_1079_p_type;
  wire [1:0] T_1079_client_id;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1107;
  wire [2:0] T_1109;
  wire [2:0] T_1111;
  wire [2:0] T_1113;
  wire [2:0] T_1115;
  wire  T_1116;
  wire [1:0] T_1121;
  wire [2:0] T_1122;
  wire [2:0] T_1131_addr_beat;
  wire [1:0] T_1131_client_xact_id;
  wire [2:0] T_1131_manager_xact_id;
  wire  T_1131_is_builtin_type;
  wire [3:0] T_1131_g_type;
  wire [4:0] T_1131_data;
  wire [1:0] T_1131_client_id;
  wire  T_1143;
  wire  T_1145;
  wire  T_1146;
  wire  T_1147;
  wire  T_1149;
  wire  T_1150;
  wire  T_1152;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire [2:0] T_1176_0;
  wire  T_1178;
  wire  T_1181;
  wire  T_1182;
  wire  T_1184;
  wire  T_1185;
  wire  T_1187;
  wire  T_1188;
  wire  T_1190;
  wire [4:0] GEN_2;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire [4:0] GEN_29;
  wire [4:0] GEN_30;
  wire [4:0] GEN_31;
  wire [4:0] GEN_32;
  wire  T_1193;
  wire  T_1194;
  wire [7:0] T_1205_0;
  wire  T_1208;
  wire  T_1209;
  wire  T_1211;
  wire  T_1212;
  wire  T_1213;
  wire [7:0] T_1214;
  wire [7:0] T_1216;
  wire [7:0] T_1217;
  wire [7:0] GEN_3;
  wire [7:0] GEN_33;
  wire [7:0] GEN_34;
  wire [7:0] GEN_35;
  wire [7:0] GEN_36;
  wire [7:0] GEN_37;
  wire [7:0] GEN_38;
  wire [7:0] GEN_39;
  wire [7:0] GEN_40;
  wire [7:0] T_1220;
  wire [7:0] T_1221;
  wire [4:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [4:0] GEN_45;
  wire [4:0] GEN_46;
  wire [4:0] GEN_47;
  wire [4:0] GEN_48;
  wire [4:0] GEN_49;
  wire [7:0] GEN_52;
  wire [7:0] GEN_53;
  wire [7:0] GEN_54;
  wire [7:0] GEN_55;
  wire [7:0] GEN_56;
  wire [7:0] GEN_57;
  wire [7:0] GEN_58;
  wire [7:0] GEN_59;
  wire [7:0] GEN_60;
  wire  GEN_61;
  wire [4:0] GEN_64;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] GEN_71;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire [7:0] GEN_78;
  wire [7:0] GEN_79;
  wire [7:0] GEN_80;
  wire [7:0] GEN_81;
  wire [7:0] GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_86;
  wire  T_1229;
  wire  T_1231;
  wire [4:0] GEN_4;
  wire [7:0] T_1247_0;
  wire [7:0] T_1259;
  wire [7:0] GEN_5;
  wire [2:0] T_1268_0;
  wire  T_1270;
  wire  T_1273;
  wire [2:0] T_1282_0;
  wire [2:0] T_1282_1;
  wire [2:0] T_1282_2;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1289;
  wire  T_1290;
  wire  T_1291;
  wire [7:0] GEN_276;
  wire [7:0] T_1292;
  wire [3:0] GEN_277;
  wire  T_1294;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire  T_1298;
  wire [1:0] T_1300;
  wire [1:0] GEN_278;
  wire [2:0] T_1301;
  wire [1:0] T_1302;
  wire [1:0] T_1305;
  wire [1:0] GEN_279;
  wire [2:0] T_1306;
  wire [1:0] T_1307;
  wire [2:0] T_1308;
  wire [2:0] GEN_280;
  wire [3:0] T_1309;
  wire [2:0] T_1310;
  wire [3:0] GEN_103;
  wire [2:0] GEN_104;
  wire [2:0] T_1311;
  wire [2:0] T_1312;
  wire [2:0] T_1313;
  wire [25:0] GEN_105;
  wire [1:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire [2:0] GEN_109;
  wire [11:0] GEN_110;
  wire [1:0] GEN_111;
  wire [4:0] GEN_113;
  wire [7:0] GEN_123;
  wire  GEN_132;
  wire [7:0] GEN_136;
  wire [3:0] GEN_137;
  wire [2:0] GEN_138;
  wire [2:0] GEN_139;
  wire  GEN_140;
  wire [25:0] GEN_141;
  wire [1:0] GEN_142;
  wire [2:0] GEN_143;
  wire  GEN_144;
  wire [2:0] GEN_145;
  wire [11:0] GEN_146;
  wire [1:0] GEN_147;
  wire [4:0] GEN_149;
  wire [7:0] GEN_159;
  wire  GEN_168;
  wire [7:0] GEN_172;
  wire [3:0] GEN_173;
  wire [2:0] GEN_174;
  wire [2:0] GEN_175;
  wire  T_1314;
  wire [1:0] GEN_281;
  wire [1:0] T_1318;
  wire [1:0] T_1319;
  wire [1:0] GEN_282;
  wire [1:0] T_1320;
  wire [3:0] GEN_176;
  wire [2:0] T_1326_0;
  wire [2:0] T_1326_1;
  wire [2:0] T_1326_2;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire  T_1339;
  wire [2:0] T_1345_0;
  wire [2:0] T_1345_1;
  wire [2:0] T_1345_2;
  wire  T_1347;
  wire  T_1348;
  wire  T_1349;
  wire  T_1352;
  wire  T_1353;
  wire [1:0] T_1357;
  wire  T_1358;
  wire [2:0] T_1361;
  wire [2:0] T_1362;
  wire [2:0] GEN_177;
  wire  GEN_178;
  wire [2:0] GEN_179;
  wire [2:0] GEN_180;
  wire  GEN_181;
  wire [2:0] GEN_182;
  wire [2:0] GEN_183;
  wire  GEN_185;
  wire [2:0] GEN_186;
  wire [2:0] GEN_187;
  wire  T_1364;
  wire [2:0] GEN_188;
  wire [2:0] GEN_189;
  wire [2:0] GEN_190;
  wire  GEN_194;
  wire  GEN_195;
  wire [2:0] GEN_196;
  wire [2:0] GEN_197;
  wire  GEN_198;
  wire [3:0] GEN_199;
  wire  GEN_203;
  wire  GEN_207;
  wire  GEN_208;
  wire [2:0] GEN_209;
  wire [2:0] GEN_210;
  wire  T_1372;
  wire  T_1374;
  wire  T_1376;
  wire [7:0] T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1380;
  wire [2:0] T_1382;
  wire  GEN_211;
  wire [2:0] GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire [2:0] GEN_215;
  wire  T_1383;
  wire [2:0] GEN_216;
  wire  GEN_217;
  wire [2:0] GEN_218;
  wire  T_1387;
  wire [3:0] GEN_283;
  wire  T_1392;
  wire  T_1393;
  wire  T_1395;
  wire [2:0] T_1397;
  wire [2:0] GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire [2:0] GEN_222;
  wire  T_1398;
  wire [2:0] GEN_223;
  wire  GEN_224;
  wire [2:0] GEN_225;
  wire  T_1410;
  wire [2:0] GEN_226;
  wire [2:0] GEN_228;
  assign io_inner_acquire_ready = GEN_140;
  assign io_inner_grant_valid = GEN_224;
  assign io_inner_grant_bits_addr_beat = T_1131_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1131_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1131_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1131_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1131_g_type;
  assign io_inner_grant_bits_data = T_1131_data;
  assign io_inner_grant_bits_client_id = T_1131_client_id;
  assign io_inner_finish_ready = T_1410;
  assign io_inner_probe_valid = GEN_198;
  assign io_inner_probe_bits_addr_block = T_1079_addr_block;
  assign io_inner_probe_bits_p_type = T_1079_p_type;
  assign io_inner_probe_bits_client_id = T_1079_client_id;
  assign io_inner_release_ready = GEN_203;
  assign io_outer_acquire_valid = GEN_217;
  assign io_outer_acquire_bits_addr_block = T_1039_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_1039_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_1039_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_1039_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_1039_a_type;
  assign io_outer_acquire_bits_union = T_1039_union;
  assign io_outer_acquire_bits_data = T_1039_data;
  assign io_outer_grant_ready = GEN_220;
  assign io_matches_iacq = T_637;
  assign io_matches_irel = T_643;
  assign io_matches_oprb = 1'h0;
  assign coh_sharers = 1'h0;
  assign T_284 = state != 3'h0;
  assign T_285 = T_284 & xact_is_builtin_type;
  assign T_294_0 = 3'h4;
  assign T_294_1 = 3'h5;
  assign T_294_2 = 3'h6;
  assign T_296 = T_294_0 == xact_a_type;
  assign T_297 = T_294_1 == xact_a_type;
  assign T_298 = T_294_2 == xact_a_type;
  assign T_301 = T_296 | T_297;
  assign T_302 = T_301 | T_298;
  assign T_303 = T_285 & T_302;
  assign T_305 = T_303 == 1'h0;
  assign T_306 = T_305 | reset;
  assign T_308 = T_306 == 1'h0;
  assign GEN_229 = $signed(1'h1);
  assign T_313 = $unsigned(GEN_229);
  assign GEN_230 = {{3'd0}, 1'h1};
  assign T_316 = GEN_230 << io_inner_acquire_bits_client_id;
  assign T_318 = ~ T_313;
  assign GEN_232 = {{3'd0}, T_318};
  assign T_319 = GEN_232 | T_316;
  assign T_320 = ~ T_319;
  assign T_321 = ~ io_incoherent_0;
  assign GEN_233 = {{3'd0}, T_321};
  assign mask_incoherent = T_320 & GEN_233;
  assign T_324 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_334_0 = 3'h3;
  assign T_336 = T_334_0 == io_inner_acquire_bits_a_type;
  assign T_339 = io_inner_acquire_bits_is_builtin_type & T_336;
  assign T_340 = T_324 & T_339;
  assign T_344 = T_342 == 3'h7;
  assign GEN_234 = {{2'd0}, 1'h1};
  assign T_346 = T_342 + GEN_234;
  assign T_347 = T_346[2:0];
  assign GEN_6 = T_340 ? T_347 : T_342;
  assign T_348 = T_340 & T_344;
  assign iacq_data_done = T_339 ? T_348 : T_324;
  assign T_350 = io_inner_release_ready & io_inner_release_valid;
  assign T_358_0 = 3'h0;
  assign T_358_1 = 3'h1;
  assign T_358_2 = 3'h2;
  assign T_360 = T_358_0 == io_inner_release_bits_r_type;
  assign T_361 = T_358_1 == io_inner_release_bits_r_type;
  assign T_362 = T_358_2 == io_inner_release_bits_r_type;
  assign T_365 = T_360 | T_361;
  assign T_366 = T_365 | T_362;
  assign T_368 = T_350 & T_366;
  assign T_374 = T_370 + GEN_234;
  assign T_375 = T_374[2:0];
  assign GEN_7 = T_368 ? T_375 : T_370;
  assign T_379 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_387_0 = 3'h5;
  assign GEN_236 = {{1'd0}, T_387_0};
  assign T_389 = GEN_236 == io_inner_grant_bits_g_type;
  assign T_397_0 = 2'h0;
  assign T_397_1 = 2'h1;
  assign GEN_237 = {{2'd0}, T_397_0};
  assign T_399 = GEN_237 == io_inner_grant_bits_g_type;
  assign GEN_238 = {{2'd0}, T_397_1};
  assign T_400 = GEN_238 == io_inner_grant_bits_g_type;
  assign T_403 = T_399 | T_400;
  assign T_404 = io_inner_grant_bits_is_builtin_type ? T_389 : T_403;
  assign T_406 = T_379 & T_404;
  assign T_410 = T_408 == 3'h7;
  assign T_412 = T_408 + GEN_234;
  assign T_413 = T_412[2:0];
  assign GEN_8 = T_406 ? T_413 : T_408;
  assign T_414 = T_406 & T_410;
  assign ignt_data_done = T_404 ? T_414 : T_379;
  assign T_416 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_425_0 = 3'h3;
  assign T_427 = T_425_0 == io_outer_acquire_bits_a_type;
  assign T_430 = io_outer_acquire_bits_is_builtin_type & T_427;
  assign T_431 = T_416 & T_430;
  assign T_435 = T_433 == 3'h7;
  assign T_437 = T_433 + GEN_234;
  assign T_438 = T_437[2:0];
  assign GEN_9 = T_431 ? T_438 : T_433;
  assign T_439 = T_431 & T_435;
  assign oacq_data_cnt = T_430 ? T_433 : {{2'd0}, 1'h0};
  assign oacq_data_done = T_430 ? T_439 : T_416;
  assign T_440 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_449_0 = 3'h5;
  assign GEN_241 = {{1'd0}, T_449_0};
  assign T_451 = GEN_241 == io_outer_grant_bits_g_type;
  assign T_459_0 = 1'h0;
  assign GEN_242 = {{3'd0}, T_459_0};
  assign T_461 = GEN_242 == io_outer_grant_bits_g_type;
  assign T_464 = io_outer_grant_bits_is_builtin_type ? T_451 : T_461;
  assign T_466 = T_440 & T_464;
  assign T_472 = T_468 + GEN_234;
  assign T_473 = T_472[2:0];
  assign GEN_10 = T_466 ? T_473 : T_468;
  assign T_485_0 = 3'h2;
  assign T_485_1 = 3'h3;
  assign T_485_2 = 3'h4;
  assign T_487 = T_485_0 == xact_a_type;
  assign T_488 = T_485_1 == xact_a_type;
  assign T_489 = T_485_2 == xact_a_type;
  assign T_492 = T_487 | T_488;
  assign T_493 = T_492 | T_489;
  assign pending_outer_write = xact_is_builtin_type & T_493;
  assign T_502_0 = 3'h2;
  assign T_502_1 = 3'h3;
  assign T_502_2 = 3'h4;
  assign T_504 = T_502_0 == io_inner_acquire_bits_a_type;
  assign T_505 = T_502_1 == io_inner_acquire_bits_a_type;
  assign T_506 = T_502_2 == io_inner_acquire_bits_a_type;
  assign T_509 = T_504 | T_505;
  assign T_510 = T_509 | T_506;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T_510;
  assign T_518_0 = 3'h5;
  assign T_518_1 = 3'h4;
  assign GEN_244 = {{1'd0}, T_518_0};
  assign T_520 = GEN_244 == io_inner_grant_bits_g_type;
  assign GEN_245 = {{1'd0}, T_518_1};
  assign T_521 = GEN_245 == io_inner_grant_bits_g_type;
  assign T_524 = T_520 | T_521;
  assign T_530_0 = 2'h0;
  assign T_530_1 = 2'h1;
  assign GEN_246 = {{2'd0}, T_530_0};
  assign T_532 = GEN_246 == io_inner_grant_bits_g_type;
  assign GEN_247 = {{2'd0}, T_530_1};
  assign T_533 = GEN_247 == io_inner_grant_bits_g_type;
  assign T_536 = T_532 | T_533;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T_524 : T_536;
  assign T_555 = 3'h6 == io_inner_acquire_bits_a_type;
  assign T_556 = T_555 ? 3'h1 : 3'h3;
  assign T_557 = 3'h5 == io_inner_acquire_bits_a_type;
  assign T_558 = T_557 ? 3'h1 : T_556;
  assign T_559 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T_560 = T_559 ? 3'h4 : T_558;
  assign T_561 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T_562 = T_561 ? 3'h3 : T_560;
  assign T_563 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T_564 = T_563 ? 3'h3 : T_562;
  assign T_565 = 3'h1 == io_inner_acquire_bits_a_type;
  assign T_566 = T_565 ? 3'h5 : T_564;
  assign T_567 = 3'h0 == io_inner_acquire_bits_a_type;
  assign T_568 = T_567 ? 3'h4 : T_566;
  assign GEN_248 = {{2'd0}, 1'h0};
  assign T_569 = io_inner_acquire_bits_a_type == GEN_248;
  assign T_574 = T_569 ? 2'h0 : 2'h1;
  assign T_575 = io_inner_acquire_bits_is_builtin_type ? T_568 : {{1'd0}, T_574};
  assign T_584_addr_beat = {{2'd0}, 1'h0};
  assign T_584_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign T_584_manager_xact_id = {{1'd0}, 2'h3};
  assign T_584_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign T_584_g_type = {{1'd0}, T_575};
  assign T_584_data = {{4'd0}, 1'h0};
  assign T_584_client_id = io_inner_acquire_bits_client_id;
  assign T_599_0 = 3'h5;
  assign T_599_1 = 3'h4;
  assign GEN_249 = {{1'd0}, T_599_0};
  assign T_601 = GEN_249 == T_584_g_type;
  assign GEN_250 = {{1'd0}, T_599_1};
  assign T_602 = GEN_250 == T_584_g_type;
  assign T_605 = T_601 | T_602;
  assign T_611_0 = 2'h0;
  assign T_611_1 = 2'h1;
  assign GEN_251 = {{2'd0}, T_611_0};
  assign T_613 = GEN_251 == T_584_g_type;
  assign GEN_252 = {{2'd0}, T_611_1};
  assign T_614 = GEN_252 == T_584_g_type;
  assign T_617 = T_613 | T_614;
  assign pending_outer_read_ = T_584_is_builtin_type ? T_605 : T_617;
  assign T_626_0 = 3'h2;
  assign T_626_1 = 3'h0;
  assign T_626_2 = 3'h4;
  assign T_628 = T_626_0 == xact_a_type;
  assign T_629 = T_626_1 == xact_a_type;
  assign T_630 = T_626_2 == xact_a_type;
  assign T_633 = T_628 | T_629;
  assign T_634 = T_633 | T_630;
  assign subblock_type = xact_is_builtin_type & T_634;
  assign T_636 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign T_637 = T_284 & T_636;
  assign T_639 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T_640 = T_284 & T_639;
  assign T_642 = io_inner_release_bits_voluntary == 1'h0;
  assign T_643 = T_640 & T_642;
  assign GEN_253 = $signed(8'hff);
  assign T_649 = $unsigned(GEN_253);
  assign T_674 = {T_649,1'h1};
  assign T_692 = 1'h1 ? {{3'd0}, T_674} : 12'h0;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign oacq_probe_client_xact_id = {{1'd0}, 2'h3};
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign oacq_probe_a_type = 3'h3;
  assign oacq_probe_union = T_692;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T_716 = xact_a_type == 3'h4;
  assign T_717 = xact_is_builtin_type & T_716;
  assign GEN_254 = {{7'd0}, 1'h1};
  assign T_721 = 8'h0 - GEN_254;
  assign T_722 = T_721[7:0];
  assign T_728_0 = T_722;
  assign T_731 = xact_a_type == 3'h3;
  assign T_732 = xact_is_builtin_type & T_731;
  assign T_734 = xact_a_type == 3'h2;
  assign T_735 = xact_is_builtin_type & T_734;
  assign T_736 = T_732 | T_735;
  assign T_737 = xact_union[8:1];
  assign T_739 = T_736 ? T_737 : {{7'd0}, 1'h0};
  assign T_740 = T_717 ? T_728_0 : T_739;
  assign T_767 = {T_740,1'h1};
  assign T_787 = 1'h1 ? {{3'd0}, T_767} : 12'h0;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_write_beat_client_xact_id = {{1'd0}, 2'h3};
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_write_beat_union = T_787;
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign GEN_0 = GEN_17;
  assign GEN_11 = GEN_234 == oacq_data_cnt ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign GEN_256 = {{1'd0}, 2'h2};
  assign GEN_12 = GEN_256 == oacq_data_cnt ? xact_wmask_buffer_2 : GEN_11;
  assign GEN_257 = {{1'd0}, 2'h3};
  assign GEN_13 = GEN_257 == oacq_data_cnt ? xact_wmask_buffer_3 : GEN_12;
  assign GEN_14 = 3'h4 == oacq_data_cnt ? xact_wmask_buffer_4 : GEN_13;
  assign GEN_15 = 3'h5 == oacq_data_cnt ? xact_wmask_buffer_5 : GEN_14;
  assign GEN_16 = 3'h6 == oacq_data_cnt ? xact_wmask_buffer_6 : GEN_15;
  assign GEN_17 = 3'h7 == oacq_data_cnt ? xact_wmask_buffer_7 : GEN_16;
  assign T_834 = {GEN_0,1'h1};
  assign T_852 = 1'h1 ? {{3'd0}, T_834} : 12'h0;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_block_client_xact_id = {{1'd0}, 2'h3};
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_block_union = T_852;
  assign oacq_write_block_data = GEN_1;
  assign GEN_1 = GEN_24;
  assign GEN_18 = GEN_234 == oacq_data_cnt ? xact_data_buffer_1 : xact_data_buffer_0;
  assign GEN_19 = GEN_256 == oacq_data_cnt ? xact_data_buffer_2 : GEN_18;
  assign GEN_20 = GEN_257 == oacq_data_cnt ? xact_data_buffer_3 : GEN_19;
  assign GEN_21 = 3'h4 == oacq_data_cnt ? xact_data_buffer_4 : GEN_20;
  assign GEN_22 = 3'h5 == oacq_data_cnt ? xact_data_buffer_5 : GEN_21;
  assign GEN_23 = 3'h6 == oacq_data_cnt ? xact_data_buffer_6 : GEN_22;
  assign GEN_24 = 3'h7 == oacq_data_cnt ? xact_data_buffer_7 : GEN_23;
  assign T_875 = xact_union[11:9];
  assign T_876 = xact_union[8:6];
  assign T_897 = {T_875,T_876};
  assign T_898 = {T_897,6'h0};
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign oacq_read_beat_client_xact_id = {{1'd0}, 2'h3};
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign oacq_read_beat_union = T_898;
  assign oacq_read_beat_data = {{4'd0}, 1'h0};
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_block_client_xact_id = {{1'd0}, 2'h3};
  assign oacq_read_block_addr_beat = {{2'd0}, 1'h0};
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_block_union = 12'h1c1;
  assign oacq_read_block_data = {{4'd0}, 1'h0};
  assign T_1013 = state == 3'h1;
  assign T_1014 = state == 3'h3;
  assign T_1015_addr_block = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign T_1015_client_xact_id = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign T_1015_addr_beat = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign T_1015_is_builtin_type = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign T_1015_a_type = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign T_1015_union = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign T_1015_data = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign T_1023_addr_block = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign T_1023_client_xact_id = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign T_1023_addr_beat = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign T_1023_is_builtin_type = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign T_1023_a_type = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign T_1023_union = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign T_1023_data = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign T_1031_addr_block = T_1014 ? T_1015_addr_block : T_1023_addr_block;
  assign T_1031_client_xact_id = T_1014 ? T_1015_client_xact_id : T_1023_client_xact_id;
  assign T_1031_addr_beat = T_1014 ? T_1015_addr_beat : T_1023_addr_beat;
  assign T_1031_is_builtin_type = T_1014 ? T_1015_is_builtin_type : T_1023_is_builtin_type;
  assign T_1031_a_type = T_1014 ? T_1015_a_type : T_1023_a_type;
  assign T_1031_union = T_1014 ? T_1015_union : T_1023_union;
  assign T_1031_data = T_1014 ? T_1015_data : T_1023_data;
  assign T_1039_addr_block = T_1013 ? oacq_probe_addr_block : T_1031_addr_block;
  assign T_1039_client_xact_id = T_1013 ? oacq_probe_client_xact_id : T_1031_client_xact_id;
  assign T_1039_addr_beat = T_1013 ? oacq_probe_addr_beat : T_1031_addr_beat;
  assign T_1039_is_builtin_type = T_1013 ? oacq_probe_is_builtin_type : T_1031_is_builtin_type;
  assign T_1039_a_type = T_1013 ? oacq_probe_a_type : T_1031_a_type;
  assign T_1039_union = T_1013 ? oacq_probe_union : T_1031_union;
  assign T_1039_data = T_1013 ? oacq_probe_data : T_1031_data;
  assign T_1056 = 3'h4 == xact_a_type;
  assign T_1057 = T_1056 ? 2'h0 : 2'h2;
  assign T_1058 = 3'h6 == xact_a_type;
  assign T_1059 = T_1058 ? 2'h0 : T_1057;
  assign T_1060 = 3'h5 == xact_a_type;
  assign T_1061 = T_1060 ? 2'h2 : T_1059;
  assign T_1062 = 3'h2 == xact_a_type;
  assign T_1063 = T_1062 ? 2'h0 : T_1061;
  assign T_1064 = 3'h0 == xact_a_type;
  assign T_1065 = T_1064 ? 2'h2 : T_1063;
  assign T_1066 = 3'h3 == xact_a_type;
  assign T_1067 = T_1066 ? 2'h0 : T_1065;
  assign T_1068 = 3'h1 == xact_a_type;
  assign T_1069 = T_1068 ? 2'h2 : T_1067;
  assign T_1070 = GEN_234 == xact_a_type;
  assign T_1071 = T_1070 ? 2'h0 : 2'h2;
  assign T_1072 = GEN_248 == xact_a_type;
  assign T_1073 = T_1072 ? 2'h1 : T_1071;
  assign T_1074 = xact_is_builtin_type ? T_1069 : T_1073;
  assign T_1079_addr_block = xact_addr_block;
  assign T_1079_p_type = T_1074;
  assign T_1079_client_id = {{1'd0}, 1'h0};
  assign T_1103 = T_1058 ? 3'h1 : 3'h3;
  assign T_1105 = T_1060 ? 3'h1 : T_1103;
  assign T_1107 = T_1056 ? 3'h4 : T_1105;
  assign T_1109 = T_1066 ? 3'h3 : T_1107;
  assign T_1111 = T_1062 ? 3'h3 : T_1109;
  assign T_1113 = T_1068 ? 3'h5 : T_1111;
  assign T_1115 = T_1064 ? 3'h4 : T_1113;
  assign T_1116 = xact_a_type == GEN_248;
  assign T_1121 = T_1116 ? 2'h0 : 2'h1;
  assign T_1122 = xact_is_builtin_type ? T_1115 : {{1'd0}, T_1121};
  assign T_1131_addr_beat = {{2'd0}, 1'h0};
  assign T_1131_client_xact_id = xact_client_xact_id;
  assign T_1131_manager_xact_id = {{1'd0}, 2'h3};
  assign T_1131_is_builtin_type = xact_is_builtin_type;
  assign T_1131_g_type = {{1'd0}, T_1122};
  assign T_1131_data = {{4'd0}, 1'h0};
  assign T_1131_client_id = xact_client_id;
  assign T_1143 = T_284 & collect_iacq_data;
  assign T_1145 = T_1143 & T_324;
  assign T_1146 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T_1147 = T_1145 & T_1146;
  assign T_1149 = T_1147 == 1'h0;
  assign T_1150 = T_1149 | reset;
  assign T_1152 = T_1150 == 1'h0;
  assign T_1157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T_1158 = T_1145 & T_1157;
  assign T_1160 = T_1158 == 1'h0;
  assign T_1161 = T_1160 | reset;
  assign T_1163 = T_1161 == 1'h0;
  assign T_1164 = state == 3'h0;
  assign T_1166 = T_1164 & T_324;
  assign T_1167 = T_1166 & io_alloc_iacq;
  assign T_1176_0 = 3'h3;
  assign T_1178 = T_1176_0 == io_inner_acquire_bits_a_type;
  assign T_1181 = io_inner_acquire_bits_is_builtin_type & T_1178;
  assign T_1182 = T_1167 & T_1181;
  assign T_1184 = io_inner_acquire_bits_addr_beat != GEN_248;
  assign T_1185 = T_1182 & T_1184;
  assign T_1187 = T_1185 == 1'h0;
  assign T_1188 = T_1187 | reset;
  assign T_1190 = T_1188 == 1'h0;
  assign GEN_2 = io_inner_acquire_bits_data;
  assign GEN_25 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_0;
  assign GEN_26 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_1;
  assign GEN_27 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_2;
  assign GEN_28 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_3;
  assign GEN_29 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_4;
  assign GEN_30 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_5;
  assign GEN_31 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_6;
  assign GEN_32 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_7;
  assign T_1193 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_1194 = io_inner_acquire_bits_is_builtin_type & T_1193;
  assign T_1205_0 = T_722;
  assign T_1208 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1209 = io_inner_acquire_bits_is_builtin_type & T_1208;
  assign T_1211 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1212 = io_inner_acquire_bits_is_builtin_type & T_1211;
  assign T_1213 = T_1209 | T_1212;
  assign T_1214 = io_inner_acquire_bits_union[8:1];
  assign T_1216 = T_1213 ? T_1214 : {{7'd0}, 1'h0};
  assign T_1217 = T_1194 ? T_1205_0 : T_1216;
  assign GEN_3 = T_1217;
  assign GEN_33 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_0;
  assign GEN_34 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_1;
  assign GEN_35 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_2;
  assign GEN_36 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_3;
  assign GEN_37 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_4;
  assign GEN_38 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_5;
  assign GEN_39 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_6;
  assign GEN_40 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_7;
  assign T_1220 = GEN_254 << io_inner_acquire_bits_addr_beat;
  assign T_1221 = iacq_data_valid | T_1220;
  assign GEN_42 = io_inner_acquire_valid ? GEN_25 : xact_data_buffer_0;
  assign GEN_43 = io_inner_acquire_valid ? GEN_26 : xact_data_buffer_1;
  assign GEN_44 = io_inner_acquire_valid ? GEN_27 : xact_data_buffer_2;
  assign GEN_45 = io_inner_acquire_valid ? GEN_28 : xact_data_buffer_3;
  assign GEN_46 = io_inner_acquire_valid ? GEN_29 : xact_data_buffer_4;
  assign GEN_47 = io_inner_acquire_valid ? GEN_30 : xact_data_buffer_5;
  assign GEN_48 = io_inner_acquire_valid ? GEN_31 : xact_data_buffer_6;
  assign GEN_49 = io_inner_acquire_valid ? GEN_32 : xact_data_buffer_7;
  assign GEN_52 = io_inner_acquire_valid ? GEN_33 : xact_wmask_buffer_0;
  assign GEN_53 = io_inner_acquire_valid ? GEN_34 : xact_wmask_buffer_1;
  assign GEN_54 = io_inner_acquire_valid ? GEN_35 : xact_wmask_buffer_2;
  assign GEN_55 = io_inner_acquire_valid ? GEN_36 : xact_wmask_buffer_3;
  assign GEN_56 = io_inner_acquire_valid ? GEN_37 : xact_wmask_buffer_4;
  assign GEN_57 = io_inner_acquire_valid ? GEN_38 : xact_wmask_buffer_5;
  assign GEN_58 = io_inner_acquire_valid ? GEN_39 : xact_wmask_buffer_6;
  assign GEN_59 = io_inner_acquire_valid ? GEN_40 : xact_wmask_buffer_7;
  assign GEN_60 = io_inner_acquire_valid ? T_1221 : iacq_data_valid;
  assign GEN_61 = iacq_data_done ? 1'h0 : collect_iacq_data;
  assign GEN_64 = collect_iacq_data ? GEN_42 : xact_data_buffer_0;
  assign GEN_65 = collect_iacq_data ? GEN_43 : xact_data_buffer_1;
  assign GEN_66 = collect_iacq_data ? GEN_44 : xact_data_buffer_2;
  assign GEN_67 = collect_iacq_data ? GEN_45 : xact_data_buffer_3;
  assign GEN_68 = collect_iacq_data ? GEN_46 : xact_data_buffer_4;
  assign GEN_69 = collect_iacq_data ? GEN_47 : xact_data_buffer_5;
  assign GEN_70 = collect_iacq_data ? GEN_48 : xact_data_buffer_6;
  assign GEN_71 = collect_iacq_data ? GEN_49 : xact_data_buffer_7;
  assign GEN_74 = collect_iacq_data ? GEN_52 : xact_wmask_buffer_0;
  assign GEN_75 = collect_iacq_data ? GEN_53 : xact_wmask_buffer_1;
  assign GEN_76 = collect_iacq_data ? GEN_54 : xact_wmask_buffer_2;
  assign GEN_77 = collect_iacq_data ? GEN_55 : xact_wmask_buffer_3;
  assign GEN_78 = collect_iacq_data ? GEN_56 : xact_wmask_buffer_4;
  assign GEN_79 = collect_iacq_data ? GEN_57 : xact_wmask_buffer_5;
  assign GEN_80 = collect_iacq_data ? GEN_58 : xact_wmask_buffer_6;
  assign GEN_81 = collect_iacq_data ? GEN_59 : xact_wmask_buffer_7;
  assign GEN_82 = collect_iacq_data ? GEN_60 : iacq_data_valid;
  assign GEN_83 = collect_iacq_data ? GEN_61 : collect_iacq_data;
  assign GEN_84 = io_outer_grant_valid ? 1'h0 : pending_ognt_ack;
  assign GEN_86 = pending_ognt_ack ? GEN_84 : pending_ognt_ack;
  assign T_1229 = 3'h0 == state;
  assign T_1231 = io_inner_acquire_valid & io_alloc_iacq;
  assign GEN_4 = io_inner_acquire_bits_data;
  assign T_1247_0 = T_722;
  assign T_1259 = T_1194 ? T_1247_0 : T_1216;
  assign GEN_5 = T_1259;
  assign T_1268_0 = 3'h3;
  assign T_1270 = T_1268_0 == io_inner_acquire_bits_a_type;
  assign T_1273 = io_inner_acquire_bits_is_builtin_type & T_1270;
  assign T_1282_0 = 3'h2;
  assign T_1282_1 = 3'h3;
  assign T_1282_2 = 3'h4;
  assign T_1284 = T_1282_0 == io_inner_acquire_bits_a_type;
  assign T_1285 = T_1282_1 == io_inner_acquire_bits_a_type;
  assign T_1286 = T_1282_2 == io_inner_acquire_bits_a_type;
  assign T_1289 = T_1284 | T_1285;
  assign T_1290 = T_1289 | T_1286;
  assign T_1291 = io_inner_acquire_bits_is_builtin_type & T_1290;
  assign GEN_276 = {{7'd0}, T_1291};
  assign T_1292 = GEN_276 << io_inner_acquire_bits_addr_beat;
  assign GEN_277 = {{3'd0}, 1'h0};
  assign T_1294 = mask_incoherent != GEN_277;
  assign T_1295 = mask_incoherent[0];
  assign T_1296 = mask_incoherent[1];
  assign T_1297 = mask_incoherent[2];
  assign T_1298 = mask_incoherent[3];
  assign T_1300 = {1'h0,T_1296};
  assign GEN_278 = {{1'd0}, T_1295};
  assign T_1301 = GEN_278 + T_1300;
  assign T_1302 = T_1301[1:0];
  assign T_1305 = {1'h0,T_1298};
  assign GEN_279 = {{1'd0}, T_1297};
  assign T_1306 = GEN_279 + T_1305;
  assign T_1307 = T_1306[1:0];
  assign T_1308 = {1'h0,T_1307};
  assign GEN_280 = {{1'd0}, T_1302};
  assign T_1309 = GEN_280 + T_1308;
  assign T_1310 = T_1309[2:0];
  assign GEN_103 = T_1294 ? mask_incoherent : {{3'd0}, pending_probes};
  assign GEN_104 = T_1294 ? T_1310 : {{2'd0}, release_count};
  assign T_1311 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign T_1312 = pending_outer_write_ ? 3'h3 : T_1311;
  assign T_1313 = T_1294 ? 3'h1 : T_1312;
  assign GEN_105 = T_1231 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_106 = T_1231 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign GEN_107 = T_1231 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign GEN_108 = T_1231 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign GEN_109 = T_1231 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign GEN_110 = T_1231 ? io_inner_acquire_bits_union : xact_union;
  assign GEN_111 = T_1231 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign GEN_113 = T_1231 ? GEN_4 : GEN_64;
  assign GEN_123 = T_1231 ? GEN_5 : GEN_74;
  assign GEN_132 = T_1231 ? T_1273 : GEN_83;
  assign GEN_136 = T_1231 ? T_1292 : GEN_82;
  assign GEN_137 = T_1231 ? GEN_103 : {{3'd0}, pending_probes};
  assign GEN_138 = T_1231 ? GEN_104 : {{2'd0}, release_count};
  assign GEN_139 = T_1231 ? T_1313 : state;
  assign GEN_140 = T_1229 ? 1'h1 : collect_iacq_data;
  assign GEN_141 = T_1229 ? GEN_105 : xact_addr_block;
  assign GEN_142 = T_1229 ? GEN_106 : xact_client_xact_id;
  assign GEN_143 = T_1229 ? GEN_107 : xact_addr_beat;
  assign GEN_144 = T_1229 ? GEN_108 : xact_is_builtin_type;
  assign GEN_145 = T_1229 ? GEN_109 : xact_a_type;
  assign GEN_146 = T_1229 ? GEN_110 : xact_union;
  assign GEN_147 = T_1229 ? GEN_111 : xact_client_id;
  assign GEN_149 = T_1229 ? GEN_113 : GEN_64;
  assign GEN_159 = T_1229 ? GEN_123 : GEN_74;
  assign GEN_168 = T_1229 ? GEN_132 : GEN_83;
  assign GEN_172 = T_1229 ? GEN_136 : GEN_82;
  assign GEN_173 = T_1229 ? GEN_137 : {{3'd0}, pending_probes};
  assign GEN_174 = T_1229 ? GEN_138 : {{2'd0}, release_count};
  assign GEN_175 = T_1229 ? GEN_139 : state;
  assign T_1314 = 3'h1 == state;
  assign GEN_281 = {{1'd0}, 1'h1};
  assign T_1318 = GEN_281 << 1'h0;
  assign T_1319 = ~ T_1318;
  assign GEN_282 = {{1'd0}, pending_probes};
  assign T_1320 = GEN_282 & T_1319;
  assign GEN_176 = io_inner_probe_ready ? {{2'd0}, T_1320} : GEN_173;
  assign T_1326_0 = 3'h0;
  assign T_1326_1 = 3'h1;
  assign T_1326_2 = 3'h2;
  assign T_1328 = T_1326_0 == io_inner_release_bits_r_type;
  assign T_1329 = T_1326_1 == io_inner_release_bits_r_type;
  assign T_1330 = T_1326_2 == io_inner_release_bits_r_type;
  assign T_1333 = T_1328 | T_1329;
  assign T_1334 = T_1333 | T_1330;
  assign T_1336 = T_1334 == 1'h0;
  assign T_1337 = T_1336 | io_outer_acquire_ready;
  assign T_1338 = T_1337 & io_matches_irel;
  assign T_1339 = io_inner_release_valid & io_matches_irel;
  assign T_1345_0 = 3'h0;
  assign T_1345_1 = 3'h1;
  assign T_1345_2 = 3'h2;
  assign T_1347 = T_1345_0 == io_inner_release_bits_r_type;
  assign T_1348 = T_1345_1 == io_inner_release_bits_r_type;
  assign T_1349 = T_1345_2 == io_inner_release_bits_r_type;
  assign T_1352 = T_1347 | T_1348;
  assign T_1353 = T_1352 | T_1349;
  assign T_1357 = release_count - 1'h1;
  assign T_1358 = T_1357[0:0];
  assign T_1361 = pending_outer_read ? 3'h2 : 3'h4;
  assign T_1362 = pending_outer_write ? 3'h3 : T_1361;
  assign GEN_177 = release_count ? T_1362 : GEN_175;
  assign GEN_178 = oacq_data_done ? 1'h1 : GEN_86;
  assign GEN_179 = oacq_data_done ? {{2'd0}, T_1358} : GEN_174;
  assign GEN_180 = oacq_data_done ? GEN_177 : GEN_175;
  assign GEN_181 = io_outer_acquire_ready ? GEN_178 : GEN_86;
  assign GEN_182 = io_outer_acquire_ready ? GEN_179 : GEN_174;
  assign GEN_183 = io_outer_acquire_ready ? GEN_180 : GEN_175;
  assign GEN_185 = T_1353 ? GEN_181 : GEN_86;
  assign GEN_186 = T_1353 ? GEN_182 : GEN_174;
  assign GEN_187 = T_1353 ? GEN_183 : GEN_175;
  assign T_1364 = T_1353 == 1'h0;
  assign GEN_188 = release_count ? T_1362 : GEN_187;
  assign GEN_189 = T_1364 ? {{2'd0}, T_1358} : GEN_186;
  assign GEN_190 = T_1364 ? GEN_188 : GEN_187;
  assign GEN_194 = T_1339 ? T_1353 : 1'h0;
  assign GEN_195 = T_1339 ? GEN_185 : GEN_86;
  assign GEN_196 = T_1339 ? GEN_189 : GEN_174;
  assign GEN_197 = T_1339 ? GEN_190 : GEN_175;
  assign GEN_198 = T_1314 ? pending_probes : 1'h0;
  assign GEN_199 = T_1314 ? GEN_176 : GEN_173;
  assign GEN_203 = T_1314 ? T_1338 : 1'h0;
  assign GEN_207 = T_1314 ? GEN_194 : 1'h0;
  assign GEN_208 = T_1314 ? GEN_195 : GEN_86;
  assign GEN_209 = T_1314 ? GEN_196 : GEN_174;
  assign GEN_210 = T_1314 ? GEN_197 : GEN_175;
  assign T_1372 = 3'h3 == state;
  assign T_1374 = pending_ognt_ack == 1'h0;
  assign T_1376 = collect_iacq_data == 1'h0;
  assign T_1377 = iacq_data_valid >> oacq_data_cnt;
  assign T_1378 = T_1377[0];
  assign T_1379 = T_1376 | T_1378;
  assign T_1380 = T_1374 & T_1379;
  assign T_1382 = pending_outer_read ? 3'h2 : 3'h5;
  assign GEN_211 = oacq_data_done ? 1'h1 : GEN_208;
  assign GEN_212 = oacq_data_done ? T_1382 : GEN_210;
  assign GEN_213 = T_1372 ? T_1380 : GEN_207;
  assign GEN_214 = T_1372 ? GEN_211 : GEN_208;
  assign GEN_215 = T_1372 ? GEN_212 : GEN_210;
  assign T_1383 = 3'h2 == state;
  assign GEN_216 = T_416 ? 3'h5 : GEN_215;
  assign GEN_217 = T_1383 ? T_1374 : GEN_213;
  assign GEN_218 = T_1383 ? GEN_216 : GEN_215;
  assign T_1387 = 3'h5 == state;
  assign GEN_283 = {{1'd0}, 3'h0};
  assign T_1392 = io_inner_grant_bits_g_type == GEN_283;
  assign T_1393 = io_inner_grant_bits_is_builtin_type & T_1392;
  assign T_1395 = T_1393 == 1'h0;
  assign T_1397 = T_1395 ? 3'h6 : 3'h0;
  assign GEN_219 = ignt_data_done ? T_1397 : GEN_218;
  assign GEN_220 = T_1387 ? io_inner_grant_ready : pending_ognt_ack;
  assign GEN_221 = T_1387 ? io_outer_grant_valid : 1'h0;
  assign GEN_222 = T_1387 ? GEN_219 : GEN_218;
  assign T_1398 = 3'h4 == state;
  assign GEN_223 = io_inner_grant_ready ? T_1397 : GEN_222;
  assign GEN_224 = T_1398 ? 1'h1 : GEN_221;
  assign GEN_225 = T_1398 ? GEN_223 : GEN_222;
  assign T_1410 = 3'h6 == state;
  assign GEN_226 = io_inner_finish_valid ? 3'h0 : GEN_225;
  assign GEN_228 = T_1410 ? GEN_226 : GEN_225;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_41 = {1{$random}};
  state = GEN_41[2:0];
  GEN_50 = {1{$random}};
  xact_addr_block = GEN_50[25:0];
  GEN_51 = {1{$random}};
  xact_client_xact_id = GEN_51[1:0];
  GEN_62 = {1{$random}};
  xact_addr_beat = GEN_62[2:0];
  GEN_63 = {1{$random}};
  xact_is_builtin_type = GEN_63[0:0];
  GEN_72 = {1{$random}};
  xact_a_type = GEN_72[2:0];
  GEN_73 = {1{$random}};
  xact_union = GEN_73[11:0];
  GEN_85 = {1{$random}};
  xact_data_buffer_0 = GEN_85[4:0];
  GEN_87 = {1{$random}};
  xact_data_buffer_1 = GEN_87[4:0];
  GEN_88 = {1{$random}};
  xact_data_buffer_2 = GEN_88[4:0];
  GEN_89 = {1{$random}};
  xact_data_buffer_3 = GEN_89[4:0];
  GEN_90 = {1{$random}};
  xact_data_buffer_4 = GEN_90[4:0];
  GEN_91 = {1{$random}};
  xact_data_buffer_5 = GEN_91[4:0];
  GEN_92 = {1{$random}};
  xact_data_buffer_6 = GEN_92[4:0];
  GEN_93 = {1{$random}};
  xact_data_buffer_7 = GEN_93[4:0];
  GEN_94 = {1{$random}};
  xact_wmask_buffer_0 = GEN_94[7:0];
  GEN_95 = {1{$random}};
  xact_wmask_buffer_1 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  xact_wmask_buffer_2 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  xact_wmask_buffer_3 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  xact_wmask_buffer_4 = GEN_98[7:0];
  GEN_99 = {1{$random}};
  xact_wmask_buffer_5 = GEN_99[7:0];
  GEN_100 = {1{$random}};
  xact_wmask_buffer_6 = GEN_100[7:0];
  GEN_101 = {1{$random}};
  xact_wmask_buffer_7 = GEN_101[7:0];
  GEN_102 = {1{$random}};
  xact_client_id = GEN_102[1:0];
  GEN_112 = {1{$random}};
  release_count = GEN_112[0:0];
  GEN_114 = {1{$random}};
  pending_probes = GEN_114[0:0];
  GEN_115 = {1{$random}};
  collect_iacq_data = GEN_115[0:0];
  GEN_116 = {1{$random}};
  iacq_data_valid = GEN_116[7:0];
  GEN_117 = {1{$random}};
  T_342 = GEN_117[2:0];
  GEN_118 = {1{$random}};
  T_370 = GEN_118[2:0];
  GEN_119 = {1{$random}};
  T_408 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  T_433 = GEN_120[2:0];
  GEN_121 = {1{$random}};
  T_468 = GEN_121[2:0];
  GEN_122 = {1{$random}};
  pending_ognt_ack = GEN_122[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_228;
    end
    if(1'h0) begin
    end else begin
      xact_addr_block <= GEN_141;
    end
    if(1'h0) begin
    end else begin
      xact_client_xact_id <= GEN_142;
    end
    if(1'h0) begin
    end else begin
      xact_addr_beat <= GEN_143;
    end
    if(1'h0) begin
    end else begin
      xact_is_builtin_type <= GEN_144;
    end
    if(1'h0) begin
    end else begin
      xact_a_type <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      xact_union <= GEN_146;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_0 <= GEN_149;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_1 <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_2 <= GEN_66;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_3 <= GEN_67;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_4 <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_5 <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_6 <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_7 <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_0 <= GEN_159;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_1 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_2 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_3 <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_4 <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_5 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_6 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_7 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      xact_client_id <= GEN_147;
    end
    if(reset) begin
      release_count <= 1'h0;
    end else begin
      release_count <= GEN_209[0];
    end
    if(reset) begin
      pending_probes <= 1'h0;
    end else begin
      pending_probes <= GEN_199[0];
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else begin
      collect_iacq_data <= GEN_168;
    end
    if(reset) begin
      iacq_data_valid <= 8'h0;
    end else begin
      iacq_data_valid <= GEN_172;
    end
    if(reset) begin
      T_342 <= 3'h0;
    end else begin
      T_342 <= GEN_6;
    end
    if(reset) begin
      T_370 <= 3'h0;
    end else begin
      T_370 <= GEN_7;
    end
    if(reset) begin
      T_408 <= 3'h0;
    end else begin
      T_408 <= GEN_8;
    end
    if(reset) begin
      T_433 <= 3'h0;
    end else begin
      T_433 <= GEN_9;
    end
    if(reset) begin
      T_468 <= 3'h0;
    end else begin
      T_468 <= GEN_10;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else begin
      pending_ognt_ack <= GEN_214;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics or prefetches\n    at broadcast.scala:203 assert(!(state =/= s_idle && xact.isBuiltInType() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different network source than initial request.\n    at broadcast.scala:285 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different client transaction than initial request.\n    at broadcast.scala:289 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at broadcast.scala:293 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module BroadcastAcquireTracker_30(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [4:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [4:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [4:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [4:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [4:0] io_outer_grant_bits_data,
  output  io_matches_iacq,
  output  io_matches_irel,
  output  io_matches_oprb,
  input   io_alloc_iacq,
  input   io_alloc_irel,
  input   io_alloc_oprb
);
  reg [2:0] state;
  reg [31:0] GEN_41;
  reg [25:0] xact_addr_block;
  reg [31:0] GEN_50;
  reg [1:0] xact_client_xact_id;
  reg [31:0] GEN_51;
  reg [2:0] xact_addr_beat;
  reg [31:0] GEN_62;
  reg  xact_is_builtin_type;
  reg [31:0] GEN_63;
  reg [2:0] xact_a_type;
  reg [31:0] GEN_72;
  reg [11:0] xact_union;
  reg [31:0] GEN_73;
  reg [4:0] xact_data_buffer_0;
  reg [31:0] GEN_85;
  reg [4:0] xact_data_buffer_1;
  reg [31:0] GEN_87;
  reg [4:0] xact_data_buffer_2;
  reg [31:0] GEN_88;
  reg [4:0] xact_data_buffer_3;
  reg [31:0] GEN_89;
  reg [4:0] xact_data_buffer_4;
  reg [31:0] GEN_90;
  reg [4:0] xact_data_buffer_5;
  reg [31:0] GEN_91;
  reg [4:0] xact_data_buffer_6;
  reg [31:0] GEN_92;
  reg [4:0] xact_data_buffer_7;
  reg [31:0] GEN_93;
  reg [7:0] xact_wmask_buffer_0;
  reg [31:0] GEN_94;
  reg [7:0] xact_wmask_buffer_1;
  reg [31:0] GEN_95;
  reg [7:0] xact_wmask_buffer_2;
  reg [31:0] GEN_96;
  reg [7:0] xact_wmask_buffer_3;
  reg [31:0] GEN_97;
  reg [7:0] xact_wmask_buffer_4;
  reg [31:0] GEN_98;
  reg [7:0] xact_wmask_buffer_5;
  reg [31:0] GEN_99;
  reg [7:0] xact_wmask_buffer_6;
  reg [31:0] GEN_100;
  reg [7:0] xact_wmask_buffer_7;
  reg [31:0] GEN_101;
  reg [1:0] xact_client_id;
  reg [31:0] GEN_102;
  wire  coh_sharers;
  wire  T_284;
  wire  T_285;
  wire [2:0] T_294_0;
  wire [2:0] T_294_1;
  wire [2:0] T_294_2;
  wire  T_296;
  wire  T_297;
  wire  T_298;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_305;
  wire  T_306;
  wire  T_308;
  reg  release_count;
  reg [31:0] GEN_112;
  reg  pending_probes;
  reg [31:0] GEN_114;
  wire  GEN_229;
  wire  T_313;
  wire [3:0] GEN_230;
  wire [3:0] T_316;
  wire  T_318;
  wire [3:0] GEN_232;
  wire [3:0] T_319;
  wire [3:0] T_320;
  wire  T_321;
  wire [3:0] GEN_233;
  wire [3:0] mask_incoherent;
  reg  collect_iacq_data;
  reg [31:0] GEN_115;
  reg [7:0] iacq_data_valid;
  reg [31:0] GEN_116;
  wire  T_324;
  wire [2:0] T_334_0;
  wire  T_336;
  wire  T_339;
  wire  T_340;
  reg [2:0] T_342;
  reg [31:0] GEN_117;
  wire  T_344;
  wire [2:0] GEN_234;
  wire [3:0] T_346;
  wire [2:0] T_347;
  wire [2:0] GEN_6;
  wire  T_348;
  wire  iacq_data_done;
  wire  T_350;
  wire [2:0] T_358_0;
  wire [2:0] T_358_1;
  wire [2:0] T_358_2;
  wire  T_360;
  wire  T_361;
  wire  T_362;
  wire  T_365;
  wire  T_366;
  wire  T_368;
  reg [2:0] T_370;
  reg [31:0] GEN_118;
  wire [3:0] T_374;
  wire [2:0] T_375;
  wire [2:0] GEN_7;
  wire  T_379;
  wire [2:0] T_387_0;
  wire [3:0] GEN_236;
  wire  T_389;
  wire [1:0] T_397_0;
  wire [1:0] T_397_1;
  wire [3:0] GEN_237;
  wire  T_399;
  wire [3:0] GEN_238;
  wire  T_400;
  wire  T_403;
  wire  T_404;
  wire  T_406;
  reg [2:0] T_408;
  reg [31:0] GEN_119;
  wire  T_410;
  wire [3:0] T_412;
  wire [2:0] T_413;
  wire [2:0] GEN_8;
  wire  T_414;
  wire  ignt_data_done;
  wire  T_416;
  wire [2:0] T_425_0;
  wire  T_427;
  wire  T_430;
  wire  T_431;
  reg [2:0] T_433;
  reg [31:0] GEN_120;
  wire  T_435;
  wire [3:0] T_437;
  wire [2:0] T_438;
  wire [2:0] GEN_9;
  wire  T_439;
  wire [2:0] oacq_data_cnt;
  wire  oacq_data_done;
  wire  T_440;
  wire [2:0] T_449_0;
  wire [3:0] GEN_241;
  wire  T_451;
  wire  T_459_0;
  wire [3:0] GEN_242;
  wire  T_461;
  wire  T_464;
  wire  T_466;
  reg [2:0] T_468;
  reg [31:0] GEN_121;
  wire [3:0] T_472;
  wire [2:0] T_473;
  wire [2:0] GEN_10;
  reg  pending_ognt_ack;
  reg [31:0] GEN_122;
  wire [2:0] T_485_0;
  wire [2:0] T_485_1;
  wire [2:0] T_485_2;
  wire  T_487;
  wire  T_488;
  wire  T_489;
  wire  T_492;
  wire  T_493;
  wire  pending_outer_write;
  wire [2:0] T_502_0;
  wire [2:0] T_502_1;
  wire [2:0] T_502_2;
  wire  T_504;
  wire  T_505;
  wire  T_506;
  wire  T_509;
  wire  T_510;
  wire  pending_outer_write_;
  wire [2:0] T_518_0;
  wire [2:0] T_518_1;
  wire [3:0] GEN_244;
  wire  T_520;
  wire [3:0] GEN_245;
  wire  T_521;
  wire  T_524;
  wire [1:0] T_530_0;
  wire [1:0] T_530_1;
  wire [3:0] GEN_246;
  wire  T_532;
  wire [3:0] GEN_247;
  wire  T_533;
  wire  T_536;
  wire  pending_outer_read;
  wire  T_555;
  wire [2:0] T_556;
  wire  T_557;
  wire [2:0] T_558;
  wire  T_559;
  wire [2:0] T_560;
  wire  T_561;
  wire [2:0] T_562;
  wire  T_563;
  wire [2:0] T_564;
  wire  T_565;
  wire [2:0] T_566;
  wire  T_567;
  wire [2:0] T_568;
  wire [2:0] GEN_248;
  wire  T_569;
  wire [1:0] T_574;
  wire [2:0] T_575;
  wire [2:0] T_584_addr_beat;
  wire [1:0] T_584_client_xact_id;
  wire [2:0] T_584_manager_xact_id;
  wire  T_584_is_builtin_type;
  wire [3:0] T_584_g_type;
  wire [4:0] T_584_data;
  wire [1:0] T_584_client_id;
  wire [2:0] T_599_0;
  wire [2:0] T_599_1;
  wire [3:0] GEN_249;
  wire  T_601;
  wire [3:0] GEN_250;
  wire  T_602;
  wire  T_605;
  wire [1:0] T_611_0;
  wire [1:0] T_611_1;
  wire [3:0] GEN_251;
  wire  T_613;
  wire [3:0] GEN_252;
  wire  T_614;
  wire  T_617;
  wire  pending_outer_read_;
  wire [2:0] T_626_0;
  wire [2:0] T_626_1;
  wire [2:0] T_626_2;
  wire  T_628;
  wire  T_629;
  wire  T_630;
  wire  T_633;
  wire  T_634;
  wire  subblock_type;
  wire  T_636;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire  T_642;
  wire  T_643;
  wire [7:0] GEN_253;
  wire [7:0] T_649;
  wire [8:0] T_674;
  wire [11:0] T_692;
  wire [25:0] oacq_probe_addr_block;
  wire [2:0] oacq_probe_client_xact_id;
  wire [2:0] oacq_probe_addr_beat;
  wire  oacq_probe_is_builtin_type;
  wire [2:0] oacq_probe_a_type;
  wire [11:0] oacq_probe_union;
  wire [4:0] oacq_probe_data;
  wire  T_716;
  wire  T_717;
  wire [7:0] GEN_254;
  wire [8:0] T_721;
  wire [7:0] T_722;
  wire [7:0] T_728_0;
  wire  T_731;
  wire  T_732;
  wire  T_734;
  wire  T_735;
  wire  T_736;
  wire [7:0] T_737;
  wire [7:0] T_739;
  wire [7:0] T_740;
  wire [8:0] T_767;
  wire [11:0] T_787;
  wire [25:0] oacq_write_beat_addr_block;
  wire [2:0] oacq_write_beat_client_xact_id;
  wire [2:0] oacq_write_beat_addr_beat;
  wire  oacq_write_beat_is_builtin_type;
  wire [2:0] oacq_write_beat_a_type;
  wire [11:0] oacq_write_beat_union;
  wire [4:0] oacq_write_beat_data;
  wire [7:0] GEN_0;
  wire [7:0] GEN_11;
  wire [2:0] GEN_256;
  wire [7:0] GEN_12;
  wire [2:0] GEN_257;
  wire [7:0] GEN_13;
  wire [7:0] GEN_14;
  wire [7:0] GEN_15;
  wire [7:0] GEN_16;
  wire [7:0] GEN_17;
  wire [8:0] T_834;
  wire [11:0] T_852;
  wire [25:0] oacq_write_block_addr_block;
  wire [2:0] oacq_write_block_client_xact_id;
  wire [2:0] oacq_write_block_addr_beat;
  wire  oacq_write_block_is_builtin_type;
  wire [2:0] oacq_write_block_a_type;
  wire [11:0] oacq_write_block_union;
  wire [4:0] oacq_write_block_data;
  wire [4:0] GEN_1;
  wire [4:0] GEN_18;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [2:0] T_875;
  wire [2:0] T_876;
  wire [5:0] T_897;
  wire [11:0] T_898;
  wire [25:0] oacq_read_beat_addr_block;
  wire [2:0] oacq_read_beat_client_xact_id;
  wire [2:0] oacq_read_beat_addr_beat;
  wire  oacq_read_beat_is_builtin_type;
  wire [2:0] oacq_read_beat_a_type;
  wire [11:0] oacq_read_beat_union;
  wire [4:0] oacq_read_beat_data;
  wire [25:0] oacq_read_block_addr_block;
  wire [2:0] oacq_read_block_client_xact_id;
  wire [2:0] oacq_read_block_addr_beat;
  wire  oacq_read_block_is_builtin_type;
  wire [2:0] oacq_read_block_a_type;
  wire [11:0] oacq_read_block_union;
  wire [4:0] oacq_read_block_data;
  wire  T_1013;
  wire  T_1014;
  wire [25:0] T_1015_addr_block;
  wire [2:0] T_1015_client_xact_id;
  wire [2:0] T_1015_addr_beat;
  wire  T_1015_is_builtin_type;
  wire [2:0] T_1015_a_type;
  wire [11:0] T_1015_union;
  wire [4:0] T_1015_data;
  wire [25:0] T_1023_addr_block;
  wire [2:0] T_1023_client_xact_id;
  wire [2:0] T_1023_addr_beat;
  wire  T_1023_is_builtin_type;
  wire [2:0] T_1023_a_type;
  wire [11:0] T_1023_union;
  wire [4:0] T_1023_data;
  wire [25:0] T_1031_addr_block;
  wire [2:0] T_1031_client_xact_id;
  wire [2:0] T_1031_addr_beat;
  wire  T_1031_is_builtin_type;
  wire [2:0] T_1031_a_type;
  wire [11:0] T_1031_union;
  wire [4:0] T_1031_data;
  wire [25:0] T_1039_addr_block;
  wire [2:0] T_1039_client_xact_id;
  wire [2:0] T_1039_addr_beat;
  wire  T_1039_is_builtin_type;
  wire [2:0] T_1039_a_type;
  wire [11:0] T_1039_union;
  wire [4:0] T_1039_data;
  wire  T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire  T_1060;
  wire [1:0] T_1061;
  wire  T_1062;
  wire [1:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire  T_1066;
  wire [1:0] T_1067;
  wire  T_1068;
  wire [1:0] T_1069;
  wire  T_1070;
  wire [1:0] T_1071;
  wire  T_1072;
  wire [1:0] T_1073;
  wire [1:0] T_1074;
  wire [25:0] T_1079_addr_block;
  wire [1:0] T_1079_p_type;
  wire [1:0] T_1079_client_id;
  wire [2:0] T_1103;
  wire [2:0] T_1105;
  wire [2:0] T_1107;
  wire [2:0] T_1109;
  wire [2:0] T_1111;
  wire [2:0] T_1113;
  wire [2:0] T_1115;
  wire  T_1116;
  wire [1:0] T_1121;
  wire [2:0] T_1122;
  wire [2:0] T_1131_addr_beat;
  wire [1:0] T_1131_client_xact_id;
  wire [2:0] T_1131_manager_xact_id;
  wire  T_1131_is_builtin_type;
  wire [3:0] T_1131_g_type;
  wire [4:0] T_1131_data;
  wire [1:0] T_1131_client_id;
  wire  T_1143;
  wire  T_1145;
  wire  T_1146;
  wire  T_1147;
  wire  T_1149;
  wire  T_1150;
  wire  T_1152;
  wire  T_1157;
  wire  T_1158;
  wire  T_1160;
  wire  T_1161;
  wire  T_1163;
  wire  T_1164;
  wire  T_1166;
  wire  T_1167;
  wire [2:0] T_1176_0;
  wire  T_1178;
  wire  T_1181;
  wire  T_1182;
  wire  T_1184;
  wire  T_1185;
  wire  T_1187;
  wire  T_1188;
  wire  T_1190;
  wire [4:0] GEN_2;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire [4:0] GEN_29;
  wire [4:0] GEN_30;
  wire [4:0] GEN_31;
  wire [4:0] GEN_32;
  wire  T_1193;
  wire  T_1194;
  wire [7:0] T_1205_0;
  wire  T_1208;
  wire  T_1209;
  wire  T_1211;
  wire  T_1212;
  wire  T_1213;
  wire [7:0] T_1214;
  wire [7:0] T_1216;
  wire [7:0] T_1217;
  wire [7:0] GEN_3;
  wire [7:0] GEN_33;
  wire [7:0] GEN_34;
  wire [7:0] GEN_35;
  wire [7:0] GEN_36;
  wire [7:0] GEN_37;
  wire [7:0] GEN_38;
  wire [7:0] GEN_39;
  wire [7:0] GEN_40;
  wire [7:0] T_1220;
  wire [7:0] T_1221;
  wire [4:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [4:0] GEN_45;
  wire [4:0] GEN_46;
  wire [4:0] GEN_47;
  wire [4:0] GEN_48;
  wire [4:0] GEN_49;
  wire [7:0] GEN_52;
  wire [7:0] GEN_53;
  wire [7:0] GEN_54;
  wire [7:0] GEN_55;
  wire [7:0] GEN_56;
  wire [7:0] GEN_57;
  wire [7:0] GEN_58;
  wire [7:0] GEN_59;
  wire [7:0] GEN_60;
  wire  GEN_61;
  wire [4:0] GEN_64;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] GEN_71;
  wire [7:0] GEN_74;
  wire [7:0] GEN_75;
  wire [7:0] GEN_76;
  wire [7:0] GEN_77;
  wire [7:0] GEN_78;
  wire [7:0] GEN_79;
  wire [7:0] GEN_80;
  wire [7:0] GEN_81;
  wire [7:0] GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_86;
  wire  T_1229;
  wire  T_1231;
  wire [4:0] GEN_4;
  wire [7:0] T_1247_0;
  wire [7:0] T_1259;
  wire [7:0] GEN_5;
  wire [2:0] T_1268_0;
  wire  T_1270;
  wire  T_1273;
  wire [2:0] T_1282_0;
  wire [2:0] T_1282_1;
  wire [2:0] T_1282_2;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1289;
  wire  T_1290;
  wire  T_1291;
  wire [7:0] GEN_276;
  wire [7:0] T_1292;
  wire [3:0] GEN_277;
  wire  T_1294;
  wire  T_1295;
  wire  T_1296;
  wire  T_1297;
  wire  T_1298;
  wire [1:0] T_1300;
  wire [1:0] GEN_278;
  wire [2:0] T_1301;
  wire [1:0] T_1302;
  wire [1:0] T_1305;
  wire [1:0] GEN_279;
  wire [2:0] T_1306;
  wire [1:0] T_1307;
  wire [2:0] T_1308;
  wire [2:0] GEN_280;
  wire [3:0] T_1309;
  wire [2:0] T_1310;
  wire [3:0] GEN_103;
  wire [2:0] GEN_104;
  wire [2:0] T_1311;
  wire [2:0] T_1312;
  wire [2:0] T_1313;
  wire [25:0] GEN_105;
  wire [1:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire [2:0] GEN_109;
  wire [11:0] GEN_110;
  wire [1:0] GEN_111;
  wire [4:0] GEN_113;
  wire [7:0] GEN_123;
  wire  GEN_132;
  wire [7:0] GEN_136;
  wire [3:0] GEN_137;
  wire [2:0] GEN_138;
  wire [2:0] GEN_139;
  wire  GEN_140;
  wire [25:0] GEN_141;
  wire [1:0] GEN_142;
  wire [2:0] GEN_143;
  wire  GEN_144;
  wire [2:0] GEN_145;
  wire [11:0] GEN_146;
  wire [1:0] GEN_147;
  wire [4:0] GEN_149;
  wire [7:0] GEN_159;
  wire  GEN_168;
  wire [7:0] GEN_172;
  wire [3:0] GEN_173;
  wire [2:0] GEN_174;
  wire [2:0] GEN_175;
  wire  T_1314;
  wire [1:0] GEN_281;
  wire [1:0] T_1318;
  wire [1:0] T_1319;
  wire [1:0] GEN_282;
  wire [1:0] T_1320;
  wire [3:0] GEN_176;
  wire [2:0] T_1326_0;
  wire [2:0] T_1326_1;
  wire [2:0] T_1326_2;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire  T_1339;
  wire [2:0] T_1345_0;
  wire [2:0] T_1345_1;
  wire [2:0] T_1345_2;
  wire  T_1347;
  wire  T_1348;
  wire  T_1349;
  wire  T_1352;
  wire  T_1353;
  wire [1:0] T_1357;
  wire  T_1358;
  wire [2:0] T_1361;
  wire [2:0] T_1362;
  wire [2:0] GEN_177;
  wire  GEN_178;
  wire [2:0] GEN_179;
  wire [2:0] GEN_180;
  wire  GEN_181;
  wire [2:0] GEN_182;
  wire [2:0] GEN_183;
  wire  GEN_185;
  wire [2:0] GEN_186;
  wire [2:0] GEN_187;
  wire  T_1364;
  wire [2:0] GEN_188;
  wire [2:0] GEN_189;
  wire [2:0] GEN_190;
  wire  GEN_194;
  wire  GEN_195;
  wire [2:0] GEN_196;
  wire [2:0] GEN_197;
  wire  GEN_198;
  wire [3:0] GEN_199;
  wire  GEN_203;
  wire  GEN_207;
  wire  GEN_208;
  wire [2:0] GEN_209;
  wire [2:0] GEN_210;
  wire  T_1372;
  wire  T_1374;
  wire  T_1376;
  wire [7:0] T_1377;
  wire  T_1378;
  wire  T_1379;
  wire  T_1380;
  wire [2:0] T_1382;
  wire  GEN_211;
  wire [2:0] GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire [2:0] GEN_215;
  wire  T_1383;
  wire [2:0] GEN_216;
  wire  GEN_217;
  wire [2:0] GEN_218;
  wire  T_1387;
  wire [3:0] GEN_283;
  wire  T_1392;
  wire  T_1393;
  wire  T_1395;
  wire [2:0] T_1397;
  wire [2:0] GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire [2:0] GEN_222;
  wire  T_1398;
  wire [2:0] GEN_223;
  wire  GEN_224;
  wire [2:0] GEN_225;
  wire  T_1410;
  wire [2:0] GEN_226;
  wire [2:0] GEN_228;
  assign io_inner_acquire_ready = GEN_140;
  assign io_inner_grant_valid = GEN_224;
  assign io_inner_grant_bits_addr_beat = T_1131_addr_beat;
  assign io_inner_grant_bits_client_xact_id = T_1131_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = T_1131_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = T_1131_is_builtin_type;
  assign io_inner_grant_bits_g_type = T_1131_g_type;
  assign io_inner_grant_bits_data = T_1131_data;
  assign io_inner_grant_bits_client_id = T_1131_client_id;
  assign io_inner_finish_ready = T_1410;
  assign io_inner_probe_valid = GEN_198;
  assign io_inner_probe_bits_addr_block = T_1079_addr_block;
  assign io_inner_probe_bits_p_type = T_1079_p_type;
  assign io_inner_probe_bits_client_id = T_1079_client_id;
  assign io_inner_release_ready = GEN_203;
  assign io_outer_acquire_valid = GEN_217;
  assign io_outer_acquire_bits_addr_block = T_1039_addr_block;
  assign io_outer_acquire_bits_client_xact_id = T_1039_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = T_1039_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = T_1039_is_builtin_type;
  assign io_outer_acquire_bits_a_type = T_1039_a_type;
  assign io_outer_acquire_bits_union = T_1039_union;
  assign io_outer_acquire_bits_data = T_1039_data;
  assign io_outer_grant_ready = GEN_220;
  assign io_matches_iacq = T_637;
  assign io_matches_irel = T_643;
  assign io_matches_oprb = 1'h0;
  assign coh_sharers = 1'h0;
  assign T_284 = state != 3'h0;
  assign T_285 = T_284 & xact_is_builtin_type;
  assign T_294_0 = 3'h4;
  assign T_294_1 = 3'h5;
  assign T_294_2 = 3'h6;
  assign T_296 = T_294_0 == xact_a_type;
  assign T_297 = T_294_1 == xact_a_type;
  assign T_298 = T_294_2 == xact_a_type;
  assign T_301 = T_296 | T_297;
  assign T_302 = T_301 | T_298;
  assign T_303 = T_285 & T_302;
  assign T_305 = T_303 == 1'h0;
  assign T_306 = T_305 | reset;
  assign T_308 = T_306 == 1'h0;
  assign GEN_229 = $signed(1'h1);
  assign T_313 = $unsigned(GEN_229);
  assign GEN_230 = {{3'd0}, 1'h1};
  assign T_316 = GEN_230 << io_inner_acquire_bits_client_id;
  assign T_318 = ~ T_313;
  assign GEN_232 = {{3'd0}, T_318};
  assign T_319 = GEN_232 | T_316;
  assign T_320 = ~ T_319;
  assign T_321 = ~ io_incoherent_0;
  assign GEN_233 = {{3'd0}, T_321};
  assign mask_incoherent = T_320 & GEN_233;
  assign T_324 = io_inner_acquire_ready & io_inner_acquire_valid;
  assign T_334_0 = 3'h3;
  assign T_336 = T_334_0 == io_inner_acquire_bits_a_type;
  assign T_339 = io_inner_acquire_bits_is_builtin_type & T_336;
  assign T_340 = T_324 & T_339;
  assign T_344 = T_342 == 3'h7;
  assign GEN_234 = {{2'd0}, 1'h1};
  assign T_346 = T_342 + GEN_234;
  assign T_347 = T_346[2:0];
  assign GEN_6 = T_340 ? T_347 : T_342;
  assign T_348 = T_340 & T_344;
  assign iacq_data_done = T_339 ? T_348 : T_324;
  assign T_350 = io_inner_release_ready & io_inner_release_valid;
  assign T_358_0 = 3'h0;
  assign T_358_1 = 3'h1;
  assign T_358_2 = 3'h2;
  assign T_360 = T_358_0 == io_inner_release_bits_r_type;
  assign T_361 = T_358_1 == io_inner_release_bits_r_type;
  assign T_362 = T_358_2 == io_inner_release_bits_r_type;
  assign T_365 = T_360 | T_361;
  assign T_366 = T_365 | T_362;
  assign T_368 = T_350 & T_366;
  assign T_374 = T_370 + GEN_234;
  assign T_375 = T_374[2:0];
  assign GEN_7 = T_368 ? T_375 : T_370;
  assign T_379 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_387_0 = 3'h5;
  assign GEN_236 = {{1'd0}, T_387_0};
  assign T_389 = GEN_236 == io_inner_grant_bits_g_type;
  assign T_397_0 = 2'h0;
  assign T_397_1 = 2'h1;
  assign GEN_237 = {{2'd0}, T_397_0};
  assign T_399 = GEN_237 == io_inner_grant_bits_g_type;
  assign GEN_238 = {{2'd0}, T_397_1};
  assign T_400 = GEN_238 == io_inner_grant_bits_g_type;
  assign T_403 = T_399 | T_400;
  assign T_404 = io_inner_grant_bits_is_builtin_type ? T_389 : T_403;
  assign T_406 = T_379 & T_404;
  assign T_410 = T_408 == 3'h7;
  assign T_412 = T_408 + GEN_234;
  assign T_413 = T_412[2:0];
  assign GEN_8 = T_406 ? T_413 : T_408;
  assign T_414 = T_406 & T_410;
  assign ignt_data_done = T_404 ? T_414 : T_379;
  assign T_416 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_425_0 = 3'h3;
  assign T_427 = T_425_0 == io_outer_acquire_bits_a_type;
  assign T_430 = io_outer_acquire_bits_is_builtin_type & T_427;
  assign T_431 = T_416 & T_430;
  assign T_435 = T_433 == 3'h7;
  assign T_437 = T_433 + GEN_234;
  assign T_438 = T_437[2:0];
  assign GEN_9 = T_431 ? T_438 : T_433;
  assign T_439 = T_431 & T_435;
  assign oacq_data_cnt = T_430 ? T_433 : {{2'd0}, 1'h0};
  assign oacq_data_done = T_430 ? T_439 : T_416;
  assign T_440 = io_outer_grant_ready & io_outer_grant_valid;
  assign T_449_0 = 3'h5;
  assign GEN_241 = {{1'd0}, T_449_0};
  assign T_451 = GEN_241 == io_outer_grant_bits_g_type;
  assign T_459_0 = 1'h0;
  assign GEN_242 = {{3'd0}, T_459_0};
  assign T_461 = GEN_242 == io_outer_grant_bits_g_type;
  assign T_464 = io_outer_grant_bits_is_builtin_type ? T_451 : T_461;
  assign T_466 = T_440 & T_464;
  assign T_472 = T_468 + GEN_234;
  assign T_473 = T_472[2:0];
  assign GEN_10 = T_466 ? T_473 : T_468;
  assign T_485_0 = 3'h2;
  assign T_485_1 = 3'h3;
  assign T_485_2 = 3'h4;
  assign T_487 = T_485_0 == xact_a_type;
  assign T_488 = T_485_1 == xact_a_type;
  assign T_489 = T_485_2 == xact_a_type;
  assign T_492 = T_487 | T_488;
  assign T_493 = T_492 | T_489;
  assign pending_outer_write = xact_is_builtin_type & T_493;
  assign T_502_0 = 3'h2;
  assign T_502_1 = 3'h3;
  assign T_502_2 = 3'h4;
  assign T_504 = T_502_0 == io_inner_acquire_bits_a_type;
  assign T_505 = T_502_1 == io_inner_acquire_bits_a_type;
  assign T_506 = T_502_2 == io_inner_acquire_bits_a_type;
  assign T_509 = T_504 | T_505;
  assign T_510 = T_509 | T_506;
  assign pending_outer_write_ = io_inner_acquire_bits_is_builtin_type & T_510;
  assign T_518_0 = 3'h5;
  assign T_518_1 = 3'h4;
  assign GEN_244 = {{1'd0}, T_518_0};
  assign T_520 = GEN_244 == io_inner_grant_bits_g_type;
  assign GEN_245 = {{1'd0}, T_518_1};
  assign T_521 = GEN_245 == io_inner_grant_bits_g_type;
  assign T_524 = T_520 | T_521;
  assign T_530_0 = 2'h0;
  assign T_530_1 = 2'h1;
  assign GEN_246 = {{2'd0}, T_530_0};
  assign T_532 = GEN_246 == io_inner_grant_bits_g_type;
  assign GEN_247 = {{2'd0}, T_530_1};
  assign T_533 = GEN_247 == io_inner_grant_bits_g_type;
  assign T_536 = T_532 | T_533;
  assign pending_outer_read = io_inner_grant_bits_is_builtin_type ? T_524 : T_536;
  assign T_555 = 3'h6 == io_inner_acquire_bits_a_type;
  assign T_556 = T_555 ? 3'h1 : 3'h3;
  assign T_557 = 3'h5 == io_inner_acquire_bits_a_type;
  assign T_558 = T_557 ? 3'h1 : T_556;
  assign T_559 = 3'h4 == io_inner_acquire_bits_a_type;
  assign T_560 = T_559 ? 3'h4 : T_558;
  assign T_561 = 3'h3 == io_inner_acquire_bits_a_type;
  assign T_562 = T_561 ? 3'h3 : T_560;
  assign T_563 = 3'h2 == io_inner_acquire_bits_a_type;
  assign T_564 = T_563 ? 3'h3 : T_562;
  assign T_565 = 3'h1 == io_inner_acquire_bits_a_type;
  assign T_566 = T_565 ? 3'h5 : T_564;
  assign T_567 = 3'h0 == io_inner_acquire_bits_a_type;
  assign T_568 = T_567 ? 3'h4 : T_566;
  assign GEN_248 = {{2'd0}, 1'h0};
  assign T_569 = io_inner_acquire_bits_a_type == GEN_248;
  assign T_574 = T_569 ? 2'h0 : 2'h1;
  assign T_575 = io_inner_acquire_bits_is_builtin_type ? T_568 : {{1'd0}, T_574};
  assign T_584_addr_beat = {{2'd0}, 1'h0};
  assign T_584_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign T_584_manager_xact_id = 3'h4;
  assign T_584_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign T_584_g_type = {{1'd0}, T_575};
  assign T_584_data = {{4'd0}, 1'h0};
  assign T_584_client_id = io_inner_acquire_bits_client_id;
  assign T_599_0 = 3'h5;
  assign T_599_1 = 3'h4;
  assign GEN_249 = {{1'd0}, T_599_0};
  assign T_601 = GEN_249 == T_584_g_type;
  assign GEN_250 = {{1'd0}, T_599_1};
  assign T_602 = GEN_250 == T_584_g_type;
  assign T_605 = T_601 | T_602;
  assign T_611_0 = 2'h0;
  assign T_611_1 = 2'h1;
  assign GEN_251 = {{2'd0}, T_611_0};
  assign T_613 = GEN_251 == T_584_g_type;
  assign GEN_252 = {{2'd0}, T_611_1};
  assign T_614 = GEN_252 == T_584_g_type;
  assign T_617 = T_613 | T_614;
  assign pending_outer_read_ = T_584_is_builtin_type ? T_605 : T_617;
  assign T_626_0 = 3'h2;
  assign T_626_1 = 3'h0;
  assign T_626_2 = 3'h4;
  assign T_628 = T_626_0 == xact_a_type;
  assign T_629 = T_626_1 == xact_a_type;
  assign T_630 = T_626_2 == xact_a_type;
  assign T_633 = T_628 | T_629;
  assign T_634 = T_633 | T_630;
  assign subblock_type = xact_is_builtin_type & T_634;
  assign T_636 = xact_addr_block == io_inner_acquire_bits_addr_block;
  assign T_637 = T_284 & T_636;
  assign T_639 = xact_addr_block == io_inner_release_bits_addr_block;
  assign T_640 = T_284 & T_639;
  assign T_642 = io_inner_release_bits_voluntary == 1'h0;
  assign T_643 = T_640 & T_642;
  assign GEN_253 = $signed(8'hff);
  assign T_649 = $unsigned(GEN_253);
  assign T_674 = {T_649,1'h1};
  assign T_692 = 1'h1 ? {{3'd0}, T_674} : 12'h0;
  assign oacq_probe_addr_block = io_inner_release_bits_addr_block;
  assign oacq_probe_client_xact_id = 3'h4;
  assign oacq_probe_addr_beat = io_inner_release_bits_addr_beat;
  assign oacq_probe_is_builtin_type = 1'h1;
  assign oacq_probe_a_type = 3'h3;
  assign oacq_probe_union = T_692;
  assign oacq_probe_data = io_inner_release_bits_data;
  assign T_716 = xact_a_type == 3'h4;
  assign T_717 = xact_is_builtin_type & T_716;
  assign GEN_254 = {{7'd0}, 1'h1};
  assign T_721 = 8'h0 - GEN_254;
  assign T_722 = T_721[7:0];
  assign T_728_0 = T_722;
  assign T_731 = xact_a_type == 3'h3;
  assign T_732 = xact_is_builtin_type & T_731;
  assign T_734 = xact_a_type == 3'h2;
  assign T_735 = xact_is_builtin_type & T_734;
  assign T_736 = T_732 | T_735;
  assign T_737 = xact_union[8:1];
  assign T_739 = T_736 ? T_737 : {{7'd0}, 1'h0};
  assign T_740 = T_717 ? T_728_0 : T_739;
  assign T_767 = {T_740,1'h1};
  assign T_787 = 1'h1 ? {{3'd0}, T_767} : 12'h0;
  assign oacq_write_beat_addr_block = xact_addr_block;
  assign oacq_write_beat_client_xact_id = 3'h4;
  assign oacq_write_beat_addr_beat = xact_addr_beat;
  assign oacq_write_beat_is_builtin_type = 1'h1;
  assign oacq_write_beat_a_type = 3'h2;
  assign oacq_write_beat_union = T_787;
  assign oacq_write_beat_data = xact_data_buffer_0;
  assign GEN_0 = GEN_17;
  assign GEN_11 = GEN_234 == oacq_data_cnt ? xact_wmask_buffer_1 : xact_wmask_buffer_0;
  assign GEN_256 = {{1'd0}, 2'h2};
  assign GEN_12 = GEN_256 == oacq_data_cnt ? xact_wmask_buffer_2 : GEN_11;
  assign GEN_257 = {{1'd0}, 2'h3};
  assign GEN_13 = GEN_257 == oacq_data_cnt ? xact_wmask_buffer_3 : GEN_12;
  assign GEN_14 = 3'h4 == oacq_data_cnt ? xact_wmask_buffer_4 : GEN_13;
  assign GEN_15 = 3'h5 == oacq_data_cnt ? xact_wmask_buffer_5 : GEN_14;
  assign GEN_16 = 3'h6 == oacq_data_cnt ? xact_wmask_buffer_6 : GEN_15;
  assign GEN_17 = 3'h7 == oacq_data_cnt ? xact_wmask_buffer_7 : GEN_16;
  assign T_834 = {GEN_0,1'h1};
  assign T_852 = 1'h1 ? {{3'd0}, T_834} : 12'h0;
  assign oacq_write_block_addr_block = xact_addr_block;
  assign oacq_write_block_client_xact_id = 3'h4;
  assign oacq_write_block_addr_beat = oacq_data_cnt;
  assign oacq_write_block_is_builtin_type = 1'h1;
  assign oacq_write_block_a_type = 3'h3;
  assign oacq_write_block_union = T_852;
  assign oacq_write_block_data = GEN_1;
  assign GEN_1 = GEN_24;
  assign GEN_18 = GEN_234 == oacq_data_cnt ? xact_data_buffer_1 : xact_data_buffer_0;
  assign GEN_19 = GEN_256 == oacq_data_cnt ? xact_data_buffer_2 : GEN_18;
  assign GEN_20 = GEN_257 == oacq_data_cnt ? xact_data_buffer_3 : GEN_19;
  assign GEN_21 = 3'h4 == oacq_data_cnt ? xact_data_buffer_4 : GEN_20;
  assign GEN_22 = 3'h5 == oacq_data_cnt ? xact_data_buffer_5 : GEN_21;
  assign GEN_23 = 3'h6 == oacq_data_cnt ? xact_data_buffer_6 : GEN_22;
  assign GEN_24 = 3'h7 == oacq_data_cnt ? xact_data_buffer_7 : GEN_23;
  assign T_875 = xact_union[11:9];
  assign T_876 = xact_union[8:6];
  assign T_897 = {T_875,T_876};
  assign T_898 = {T_897,6'h0};
  assign oacq_read_beat_addr_block = xact_addr_block;
  assign oacq_read_beat_client_xact_id = 3'h4;
  assign oacq_read_beat_addr_beat = xact_addr_beat;
  assign oacq_read_beat_is_builtin_type = 1'h1;
  assign oacq_read_beat_a_type = 3'h0;
  assign oacq_read_beat_union = T_898;
  assign oacq_read_beat_data = {{4'd0}, 1'h0};
  assign oacq_read_block_addr_block = xact_addr_block;
  assign oacq_read_block_client_xact_id = 3'h4;
  assign oacq_read_block_addr_beat = {{2'd0}, 1'h0};
  assign oacq_read_block_is_builtin_type = 1'h1;
  assign oacq_read_block_a_type = 3'h1;
  assign oacq_read_block_union = 12'h1c1;
  assign oacq_read_block_data = {{4'd0}, 1'h0};
  assign T_1013 = state == 3'h1;
  assign T_1014 = state == 3'h3;
  assign T_1015_addr_block = subblock_type ? oacq_write_beat_addr_block : oacq_write_block_addr_block;
  assign T_1015_client_xact_id = subblock_type ? oacq_write_beat_client_xact_id : oacq_write_block_client_xact_id;
  assign T_1015_addr_beat = subblock_type ? oacq_write_beat_addr_beat : oacq_write_block_addr_beat;
  assign T_1015_is_builtin_type = subblock_type ? oacq_write_beat_is_builtin_type : oacq_write_block_is_builtin_type;
  assign T_1015_a_type = subblock_type ? oacq_write_beat_a_type : oacq_write_block_a_type;
  assign T_1015_union = subblock_type ? oacq_write_beat_union : oacq_write_block_union;
  assign T_1015_data = subblock_type ? oacq_write_beat_data : oacq_write_block_data;
  assign T_1023_addr_block = subblock_type ? oacq_read_beat_addr_block : oacq_read_block_addr_block;
  assign T_1023_client_xact_id = subblock_type ? oacq_read_beat_client_xact_id : oacq_read_block_client_xact_id;
  assign T_1023_addr_beat = subblock_type ? oacq_read_beat_addr_beat : oacq_read_block_addr_beat;
  assign T_1023_is_builtin_type = subblock_type ? oacq_read_beat_is_builtin_type : oacq_read_block_is_builtin_type;
  assign T_1023_a_type = subblock_type ? oacq_read_beat_a_type : oacq_read_block_a_type;
  assign T_1023_union = subblock_type ? oacq_read_beat_union : oacq_read_block_union;
  assign T_1023_data = subblock_type ? oacq_read_beat_data : oacq_read_block_data;
  assign T_1031_addr_block = T_1014 ? T_1015_addr_block : T_1023_addr_block;
  assign T_1031_client_xact_id = T_1014 ? T_1015_client_xact_id : T_1023_client_xact_id;
  assign T_1031_addr_beat = T_1014 ? T_1015_addr_beat : T_1023_addr_beat;
  assign T_1031_is_builtin_type = T_1014 ? T_1015_is_builtin_type : T_1023_is_builtin_type;
  assign T_1031_a_type = T_1014 ? T_1015_a_type : T_1023_a_type;
  assign T_1031_union = T_1014 ? T_1015_union : T_1023_union;
  assign T_1031_data = T_1014 ? T_1015_data : T_1023_data;
  assign T_1039_addr_block = T_1013 ? oacq_probe_addr_block : T_1031_addr_block;
  assign T_1039_client_xact_id = T_1013 ? oacq_probe_client_xact_id : T_1031_client_xact_id;
  assign T_1039_addr_beat = T_1013 ? oacq_probe_addr_beat : T_1031_addr_beat;
  assign T_1039_is_builtin_type = T_1013 ? oacq_probe_is_builtin_type : T_1031_is_builtin_type;
  assign T_1039_a_type = T_1013 ? oacq_probe_a_type : T_1031_a_type;
  assign T_1039_union = T_1013 ? oacq_probe_union : T_1031_union;
  assign T_1039_data = T_1013 ? oacq_probe_data : T_1031_data;
  assign T_1056 = 3'h4 == xact_a_type;
  assign T_1057 = T_1056 ? 2'h0 : 2'h2;
  assign T_1058 = 3'h6 == xact_a_type;
  assign T_1059 = T_1058 ? 2'h0 : T_1057;
  assign T_1060 = 3'h5 == xact_a_type;
  assign T_1061 = T_1060 ? 2'h2 : T_1059;
  assign T_1062 = 3'h2 == xact_a_type;
  assign T_1063 = T_1062 ? 2'h0 : T_1061;
  assign T_1064 = 3'h0 == xact_a_type;
  assign T_1065 = T_1064 ? 2'h2 : T_1063;
  assign T_1066 = 3'h3 == xact_a_type;
  assign T_1067 = T_1066 ? 2'h0 : T_1065;
  assign T_1068 = 3'h1 == xact_a_type;
  assign T_1069 = T_1068 ? 2'h2 : T_1067;
  assign T_1070 = GEN_234 == xact_a_type;
  assign T_1071 = T_1070 ? 2'h0 : 2'h2;
  assign T_1072 = GEN_248 == xact_a_type;
  assign T_1073 = T_1072 ? 2'h1 : T_1071;
  assign T_1074 = xact_is_builtin_type ? T_1069 : T_1073;
  assign T_1079_addr_block = xact_addr_block;
  assign T_1079_p_type = T_1074;
  assign T_1079_client_id = {{1'd0}, 1'h0};
  assign T_1103 = T_1058 ? 3'h1 : 3'h3;
  assign T_1105 = T_1060 ? 3'h1 : T_1103;
  assign T_1107 = T_1056 ? 3'h4 : T_1105;
  assign T_1109 = T_1066 ? 3'h3 : T_1107;
  assign T_1111 = T_1062 ? 3'h3 : T_1109;
  assign T_1113 = T_1068 ? 3'h5 : T_1111;
  assign T_1115 = T_1064 ? 3'h4 : T_1113;
  assign T_1116 = xact_a_type == GEN_248;
  assign T_1121 = T_1116 ? 2'h0 : 2'h1;
  assign T_1122 = xact_is_builtin_type ? T_1115 : {{1'd0}, T_1121};
  assign T_1131_addr_beat = {{2'd0}, 1'h0};
  assign T_1131_client_xact_id = xact_client_xact_id;
  assign T_1131_manager_xact_id = 3'h4;
  assign T_1131_is_builtin_type = xact_is_builtin_type;
  assign T_1131_g_type = {{1'd0}, T_1122};
  assign T_1131_data = {{4'd0}, 1'h0};
  assign T_1131_client_id = xact_client_id;
  assign T_1143 = T_284 & collect_iacq_data;
  assign T_1145 = T_1143 & T_324;
  assign T_1146 = io_inner_acquire_bits_client_id != xact_client_id;
  assign T_1147 = T_1145 & T_1146;
  assign T_1149 = T_1147 == 1'h0;
  assign T_1150 = T_1149 | reset;
  assign T_1152 = T_1150 == 1'h0;
  assign T_1157 = io_inner_acquire_bits_client_xact_id != xact_client_xact_id;
  assign T_1158 = T_1145 & T_1157;
  assign T_1160 = T_1158 == 1'h0;
  assign T_1161 = T_1160 | reset;
  assign T_1163 = T_1161 == 1'h0;
  assign T_1164 = state == 3'h0;
  assign T_1166 = T_1164 & T_324;
  assign T_1167 = T_1166 & io_alloc_iacq;
  assign T_1176_0 = 3'h3;
  assign T_1178 = T_1176_0 == io_inner_acquire_bits_a_type;
  assign T_1181 = io_inner_acquire_bits_is_builtin_type & T_1178;
  assign T_1182 = T_1167 & T_1181;
  assign T_1184 = io_inner_acquire_bits_addr_beat != GEN_248;
  assign T_1185 = T_1182 & T_1184;
  assign T_1187 = T_1185 == 1'h0;
  assign T_1188 = T_1187 | reset;
  assign T_1190 = T_1188 == 1'h0;
  assign GEN_2 = io_inner_acquire_bits_data;
  assign GEN_25 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_0;
  assign GEN_26 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_1;
  assign GEN_27 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_2;
  assign GEN_28 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_3;
  assign GEN_29 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_4;
  assign GEN_30 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_5;
  assign GEN_31 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_6;
  assign GEN_32 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_2 : xact_data_buffer_7;
  assign T_1193 = io_inner_acquire_bits_a_type == 3'h4;
  assign T_1194 = io_inner_acquire_bits_is_builtin_type & T_1193;
  assign T_1205_0 = T_722;
  assign T_1208 = io_inner_acquire_bits_a_type == 3'h3;
  assign T_1209 = io_inner_acquire_bits_is_builtin_type & T_1208;
  assign T_1211 = io_inner_acquire_bits_a_type == 3'h2;
  assign T_1212 = io_inner_acquire_bits_is_builtin_type & T_1211;
  assign T_1213 = T_1209 | T_1212;
  assign T_1214 = io_inner_acquire_bits_union[8:1];
  assign T_1216 = T_1213 ? T_1214 : {{7'd0}, 1'h0};
  assign T_1217 = T_1194 ? T_1205_0 : T_1216;
  assign GEN_3 = T_1217;
  assign GEN_33 = GEN_248 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_0;
  assign GEN_34 = GEN_234 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_1;
  assign GEN_35 = GEN_256 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_2;
  assign GEN_36 = GEN_257 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_3;
  assign GEN_37 = 3'h4 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_4;
  assign GEN_38 = 3'h5 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_5;
  assign GEN_39 = 3'h6 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_6;
  assign GEN_40 = 3'h7 == io_inner_acquire_bits_addr_beat ? GEN_3 : xact_wmask_buffer_7;
  assign T_1220 = GEN_254 << io_inner_acquire_bits_addr_beat;
  assign T_1221 = iacq_data_valid | T_1220;
  assign GEN_42 = io_inner_acquire_valid ? GEN_25 : xact_data_buffer_0;
  assign GEN_43 = io_inner_acquire_valid ? GEN_26 : xact_data_buffer_1;
  assign GEN_44 = io_inner_acquire_valid ? GEN_27 : xact_data_buffer_2;
  assign GEN_45 = io_inner_acquire_valid ? GEN_28 : xact_data_buffer_3;
  assign GEN_46 = io_inner_acquire_valid ? GEN_29 : xact_data_buffer_4;
  assign GEN_47 = io_inner_acquire_valid ? GEN_30 : xact_data_buffer_5;
  assign GEN_48 = io_inner_acquire_valid ? GEN_31 : xact_data_buffer_6;
  assign GEN_49 = io_inner_acquire_valid ? GEN_32 : xact_data_buffer_7;
  assign GEN_52 = io_inner_acquire_valid ? GEN_33 : xact_wmask_buffer_0;
  assign GEN_53 = io_inner_acquire_valid ? GEN_34 : xact_wmask_buffer_1;
  assign GEN_54 = io_inner_acquire_valid ? GEN_35 : xact_wmask_buffer_2;
  assign GEN_55 = io_inner_acquire_valid ? GEN_36 : xact_wmask_buffer_3;
  assign GEN_56 = io_inner_acquire_valid ? GEN_37 : xact_wmask_buffer_4;
  assign GEN_57 = io_inner_acquire_valid ? GEN_38 : xact_wmask_buffer_5;
  assign GEN_58 = io_inner_acquire_valid ? GEN_39 : xact_wmask_buffer_6;
  assign GEN_59 = io_inner_acquire_valid ? GEN_40 : xact_wmask_buffer_7;
  assign GEN_60 = io_inner_acquire_valid ? T_1221 : iacq_data_valid;
  assign GEN_61 = iacq_data_done ? 1'h0 : collect_iacq_data;
  assign GEN_64 = collect_iacq_data ? GEN_42 : xact_data_buffer_0;
  assign GEN_65 = collect_iacq_data ? GEN_43 : xact_data_buffer_1;
  assign GEN_66 = collect_iacq_data ? GEN_44 : xact_data_buffer_2;
  assign GEN_67 = collect_iacq_data ? GEN_45 : xact_data_buffer_3;
  assign GEN_68 = collect_iacq_data ? GEN_46 : xact_data_buffer_4;
  assign GEN_69 = collect_iacq_data ? GEN_47 : xact_data_buffer_5;
  assign GEN_70 = collect_iacq_data ? GEN_48 : xact_data_buffer_6;
  assign GEN_71 = collect_iacq_data ? GEN_49 : xact_data_buffer_7;
  assign GEN_74 = collect_iacq_data ? GEN_52 : xact_wmask_buffer_0;
  assign GEN_75 = collect_iacq_data ? GEN_53 : xact_wmask_buffer_1;
  assign GEN_76 = collect_iacq_data ? GEN_54 : xact_wmask_buffer_2;
  assign GEN_77 = collect_iacq_data ? GEN_55 : xact_wmask_buffer_3;
  assign GEN_78 = collect_iacq_data ? GEN_56 : xact_wmask_buffer_4;
  assign GEN_79 = collect_iacq_data ? GEN_57 : xact_wmask_buffer_5;
  assign GEN_80 = collect_iacq_data ? GEN_58 : xact_wmask_buffer_6;
  assign GEN_81 = collect_iacq_data ? GEN_59 : xact_wmask_buffer_7;
  assign GEN_82 = collect_iacq_data ? GEN_60 : iacq_data_valid;
  assign GEN_83 = collect_iacq_data ? GEN_61 : collect_iacq_data;
  assign GEN_84 = io_outer_grant_valid ? 1'h0 : pending_ognt_ack;
  assign GEN_86 = pending_ognt_ack ? GEN_84 : pending_ognt_ack;
  assign T_1229 = 3'h0 == state;
  assign T_1231 = io_inner_acquire_valid & io_alloc_iacq;
  assign GEN_4 = io_inner_acquire_bits_data;
  assign T_1247_0 = T_722;
  assign T_1259 = T_1194 ? T_1247_0 : T_1216;
  assign GEN_5 = T_1259;
  assign T_1268_0 = 3'h3;
  assign T_1270 = T_1268_0 == io_inner_acquire_bits_a_type;
  assign T_1273 = io_inner_acquire_bits_is_builtin_type & T_1270;
  assign T_1282_0 = 3'h2;
  assign T_1282_1 = 3'h3;
  assign T_1282_2 = 3'h4;
  assign T_1284 = T_1282_0 == io_inner_acquire_bits_a_type;
  assign T_1285 = T_1282_1 == io_inner_acquire_bits_a_type;
  assign T_1286 = T_1282_2 == io_inner_acquire_bits_a_type;
  assign T_1289 = T_1284 | T_1285;
  assign T_1290 = T_1289 | T_1286;
  assign T_1291 = io_inner_acquire_bits_is_builtin_type & T_1290;
  assign GEN_276 = {{7'd0}, T_1291};
  assign T_1292 = GEN_276 << io_inner_acquire_bits_addr_beat;
  assign GEN_277 = {{3'd0}, 1'h0};
  assign T_1294 = mask_incoherent != GEN_277;
  assign T_1295 = mask_incoherent[0];
  assign T_1296 = mask_incoherent[1];
  assign T_1297 = mask_incoherent[2];
  assign T_1298 = mask_incoherent[3];
  assign T_1300 = {1'h0,T_1296};
  assign GEN_278 = {{1'd0}, T_1295};
  assign T_1301 = GEN_278 + T_1300;
  assign T_1302 = T_1301[1:0];
  assign T_1305 = {1'h0,T_1298};
  assign GEN_279 = {{1'd0}, T_1297};
  assign T_1306 = GEN_279 + T_1305;
  assign T_1307 = T_1306[1:0];
  assign T_1308 = {1'h0,T_1307};
  assign GEN_280 = {{1'd0}, T_1302};
  assign T_1309 = GEN_280 + T_1308;
  assign T_1310 = T_1309[2:0];
  assign GEN_103 = T_1294 ? mask_incoherent : {{3'd0}, pending_probes};
  assign GEN_104 = T_1294 ? T_1310 : {{2'd0}, release_count};
  assign T_1311 = pending_outer_read_ ? 3'h2 : 3'h4;
  assign T_1312 = pending_outer_write_ ? 3'h3 : T_1311;
  assign T_1313 = T_1294 ? 3'h1 : T_1312;
  assign GEN_105 = T_1231 ? io_inner_acquire_bits_addr_block : xact_addr_block;
  assign GEN_106 = T_1231 ? io_inner_acquire_bits_client_xact_id : xact_client_xact_id;
  assign GEN_107 = T_1231 ? io_inner_acquire_bits_addr_beat : xact_addr_beat;
  assign GEN_108 = T_1231 ? io_inner_acquire_bits_is_builtin_type : xact_is_builtin_type;
  assign GEN_109 = T_1231 ? io_inner_acquire_bits_a_type : xact_a_type;
  assign GEN_110 = T_1231 ? io_inner_acquire_bits_union : xact_union;
  assign GEN_111 = T_1231 ? io_inner_acquire_bits_client_id : xact_client_id;
  assign GEN_113 = T_1231 ? GEN_4 : GEN_64;
  assign GEN_123 = T_1231 ? GEN_5 : GEN_74;
  assign GEN_132 = T_1231 ? T_1273 : GEN_83;
  assign GEN_136 = T_1231 ? T_1292 : GEN_82;
  assign GEN_137 = T_1231 ? GEN_103 : {{3'd0}, pending_probes};
  assign GEN_138 = T_1231 ? GEN_104 : {{2'd0}, release_count};
  assign GEN_139 = T_1231 ? T_1313 : state;
  assign GEN_140 = T_1229 ? 1'h1 : collect_iacq_data;
  assign GEN_141 = T_1229 ? GEN_105 : xact_addr_block;
  assign GEN_142 = T_1229 ? GEN_106 : xact_client_xact_id;
  assign GEN_143 = T_1229 ? GEN_107 : xact_addr_beat;
  assign GEN_144 = T_1229 ? GEN_108 : xact_is_builtin_type;
  assign GEN_145 = T_1229 ? GEN_109 : xact_a_type;
  assign GEN_146 = T_1229 ? GEN_110 : xact_union;
  assign GEN_147 = T_1229 ? GEN_111 : xact_client_id;
  assign GEN_149 = T_1229 ? GEN_113 : GEN_64;
  assign GEN_159 = T_1229 ? GEN_123 : GEN_74;
  assign GEN_168 = T_1229 ? GEN_132 : GEN_83;
  assign GEN_172 = T_1229 ? GEN_136 : GEN_82;
  assign GEN_173 = T_1229 ? GEN_137 : {{3'd0}, pending_probes};
  assign GEN_174 = T_1229 ? GEN_138 : {{2'd0}, release_count};
  assign GEN_175 = T_1229 ? GEN_139 : state;
  assign T_1314 = 3'h1 == state;
  assign GEN_281 = {{1'd0}, 1'h1};
  assign T_1318 = GEN_281 << 1'h0;
  assign T_1319 = ~ T_1318;
  assign GEN_282 = {{1'd0}, pending_probes};
  assign T_1320 = GEN_282 & T_1319;
  assign GEN_176 = io_inner_probe_ready ? {{2'd0}, T_1320} : GEN_173;
  assign T_1326_0 = 3'h0;
  assign T_1326_1 = 3'h1;
  assign T_1326_2 = 3'h2;
  assign T_1328 = T_1326_0 == io_inner_release_bits_r_type;
  assign T_1329 = T_1326_1 == io_inner_release_bits_r_type;
  assign T_1330 = T_1326_2 == io_inner_release_bits_r_type;
  assign T_1333 = T_1328 | T_1329;
  assign T_1334 = T_1333 | T_1330;
  assign T_1336 = T_1334 == 1'h0;
  assign T_1337 = T_1336 | io_outer_acquire_ready;
  assign T_1338 = T_1337 & io_matches_irel;
  assign T_1339 = io_inner_release_valid & io_matches_irel;
  assign T_1345_0 = 3'h0;
  assign T_1345_1 = 3'h1;
  assign T_1345_2 = 3'h2;
  assign T_1347 = T_1345_0 == io_inner_release_bits_r_type;
  assign T_1348 = T_1345_1 == io_inner_release_bits_r_type;
  assign T_1349 = T_1345_2 == io_inner_release_bits_r_type;
  assign T_1352 = T_1347 | T_1348;
  assign T_1353 = T_1352 | T_1349;
  assign T_1357 = release_count - 1'h1;
  assign T_1358 = T_1357[0:0];
  assign T_1361 = pending_outer_read ? 3'h2 : 3'h4;
  assign T_1362 = pending_outer_write ? 3'h3 : T_1361;
  assign GEN_177 = release_count ? T_1362 : GEN_175;
  assign GEN_178 = oacq_data_done ? 1'h1 : GEN_86;
  assign GEN_179 = oacq_data_done ? {{2'd0}, T_1358} : GEN_174;
  assign GEN_180 = oacq_data_done ? GEN_177 : GEN_175;
  assign GEN_181 = io_outer_acquire_ready ? GEN_178 : GEN_86;
  assign GEN_182 = io_outer_acquire_ready ? GEN_179 : GEN_174;
  assign GEN_183 = io_outer_acquire_ready ? GEN_180 : GEN_175;
  assign GEN_185 = T_1353 ? GEN_181 : GEN_86;
  assign GEN_186 = T_1353 ? GEN_182 : GEN_174;
  assign GEN_187 = T_1353 ? GEN_183 : GEN_175;
  assign T_1364 = T_1353 == 1'h0;
  assign GEN_188 = release_count ? T_1362 : GEN_187;
  assign GEN_189 = T_1364 ? {{2'd0}, T_1358} : GEN_186;
  assign GEN_190 = T_1364 ? GEN_188 : GEN_187;
  assign GEN_194 = T_1339 ? T_1353 : 1'h0;
  assign GEN_195 = T_1339 ? GEN_185 : GEN_86;
  assign GEN_196 = T_1339 ? GEN_189 : GEN_174;
  assign GEN_197 = T_1339 ? GEN_190 : GEN_175;
  assign GEN_198 = T_1314 ? pending_probes : 1'h0;
  assign GEN_199 = T_1314 ? GEN_176 : GEN_173;
  assign GEN_203 = T_1314 ? T_1338 : 1'h0;
  assign GEN_207 = T_1314 ? GEN_194 : 1'h0;
  assign GEN_208 = T_1314 ? GEN_195 : GEN_86;
  assign GEN_209 = T_1314 ? GEN_196 : GEN_174;
  assign GEN_210 = T_1314 ? GEN_197 : GEN_175;
  assign T_1372 = 3'h3 == state;
  assign T_1374 = pending_ognt_ack == 1'h0;
  assign T_1376 = collect_iacq_data == 1'h0;
  assign T_1377 = iacq_data_valid >> oacq_data_cnt;
  assign T_1378 = T_1377[0];
  assign T_1379 = T_1376 | T_1378;
  assign T_1380 = T_1374 & T_1379;
  assign T_1382 = pending_outer_read ? 3'h2 : 3'h5;
  assign GEN_211 = oacq_data_done ? 1'h1 : GEN_208;
  assign GEN_212 = oacq_data_done ? T_1382 : GEN_210;
  assign GEN_213 = T_1372 ? T_1380 : GEN_207;
  assign GEN_214 = T_1372 ? GEN_211 : GEN_208;
  assign GEN_215 = T_1372 ? GEN_212 : GEN_210;
  assign T_1383 = 3'h2 == state;
  assign GEN_216 = T_416 ? 3'h5 : GEN_215;
  assign GEN_217 = T_1383 ? T_1374 : GEN_213;
  assign GEN_218 = T_1383 ? GEN_216 : GEN_215;
  assign T_1387 = 3'h5 == state;
  assign GEN_283 = {{1'd0}, 3'h0};
  assign T_1392 = io_inner_grant_bits_g_type == GEN_283;
  assign T_1393 = io_inner_grant_bits_is_builtin_type & T_1392;
  assign T_1395 = T_1393 == 1'h0;
  assign T_1397 = T_1395 ? 3'h6 : 3'h0;
  assign GEN_219 = ignt_data_done ? T_1397 : GEN_218;
  assign GEN_220 = T_1387 ? io_inner_grant_ready : pending_ognt_ack;
  assign GEN_221 = T_1387 ? io_outer_grant_valid : 1'h0;
  assign GEN_222 = T_1387 ? GEN_219 : GEN_218;
  assign T_1398 = 3'h4 == state;
  assign GEN_223 = io_inner_grant_ready ? T_1397 : GEN_222;
  assign GEN_224 = T_1398 ? 1'h1 : GEN_221;
  assign GEN_225 = T_1398 ? GEN_223 : GEN_222;
  assign T_1410 = 3'h6 == state;
  assign GEN_226 = io_inner_finish_valid ? 3'h0 : GEN_225;
  assign GEN_228 = T_1410 ? GEN_226 : GEN_225;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_41 = {1{$random}};
  state = GEN_41[2:0];
  GEN_50 = {1{$random}};
  xact_addr_block = GEN_50[25:0];
  GEN_51 = {1{$random}};
  xact_client_xact_id = GEN_51[1:0];
  GEN_62 = {1{$random}};
  xact_addr_beat = GEN_62[2:0];
  GEN_63 = {1{$random}};
  xact_is_builtin_type = GEN_63[0:0];
  GEN_72 = {1{$random}};
  xact_a_type = GEN_72[2:0];
  GEN_73 = {1{$random}};
  xact_union = GEN_73[11:0];
  GEN_85 = {1{$random}};
  xact_data_buffer_0 = GEN_85[4:0];
  GEN_87 = {1{$random}};
  xact_data_buffer_1 = GEN_87[4:0];
  GEN_88 = {1{$random}};
  xact_data_buffer_2 = GEN_88[4:0];
  GEN_89 = {1{$random}};
  xact_data_buffer_3 = GEN_89[4:0];
  GEN_90 = {1{$random}};
  xact_data_buffer_4 = GEN_90[4:0];
  GEN_91 = {1{$random}};
  xact_data_buffer_5 = GEN_91[4:0];
  GEN_92 = {1{$random}};
  xact_data_buffer_6 = GEN_92[4:0];
  GEN_93 = {1{$random}};
  xact_data_buffer_7 = GEN_93[4:0];
  GEN_94 = {1{$random}};
  xact_wmask_buffer_0 = GEN_94[7:0];
  GEN_95 = {1{$random}};
  xact_wmask_buffer_1 = GEN_95[7:0];
  GEN_96 = {1{$random}};
  xact_wmask_buffer_2 = GEN_96[7:0];
  GEN_97 = {1{$random}};
  xact_wmask_buffer_3 = GEN_97[7:0];
  GEN_98 = {1{$random}};
  xact_wmask_buffer_4 = GEN_98[7:0];
  GEN_99 = {1{$random}};
  xact_wmask_buffer_5 = GEN_99[7:0];
  GEN_100 = {1{$random}};
  xact_wmask_buffer_6 = GEN_100[7:0];
  GEN_101 = {1{$random}};
  xact_wmask_buffer_7 = GEN_101[7:0];
  GEN_102 = {1{$random}};
  xact_client_id = GEN_102[1:0];
  GEN_112 = {1{$random}};
  release_count = GEN_112[0:0];
  GEN_114 = {1{$random}};
  pending_probes = GEN_114[0:0];
  GEN_115 = {1{$random}};
  collect_iacq_data = GEN_115[0:0];
  GEN_116 = {1{$random}};
  iacq_data_valid = GEN_116[7:0];
  GEN_117 = {1{$random}};
  T_342 = GEN_117[2:0];
  GEN_118 = {1{$random}};
  T_370 = GEN_118[2:0];
  GEN_119 = {1{$random}};
  T_408 = GEN_119[2:0];
  GEN_120 = {1{$random}};
  T_433 = GEN_120[2:0];
  GEN_121 = {1{$random}};
  T_468 = GEN_121[2:0];
  GEN_122 = {1{$random}};
  pending_ognt_ack = GEN_122[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_228;
    end
    if(1'h0) begin
    end else begin
      xact_addr_block <= GEN_141;
    end
    if(1'h0) begin
    end else begin
      xact_client_xact_id <= GEN_142;
    end
    if(1'h0) begin
    end else begin
      xact_addr_beat <= GEN_143;
    end
    if(1'h0) begin
    end else begin
      xact_is_builtin_type <= GEN_144;
    end
    if(1'h0) begin
    end else begin
      xact_a_type <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      xact_union <= GEN_146;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_0 <= GEN_149;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_1 <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_2 <= GEN_66;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_3 <= GEN_67;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_4 <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_5 <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_6 <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      xact_data_buffer_7 <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_0 <= GEN_159;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_1 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_2 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_3 <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_4 <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_5 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_6 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      xact_wmask_buffer_7 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      xact_client_id <= GEN_147;
    end
    if(reset) begin
      release_count <= 1'h0;
    end else begin
      release_count <= GEN_209[0];
    end
    if(reset) begin
      pending_probes <= 1'h0;
    end else begin
      pending_probes <= GEN_199[0];
    end
    if(reset) begin
      collect_iacq_data <= 1'h0;
    end else begin
      collect_iacq_data <= GEN_168;
    end
    if(reset) begin
      iacq_data_valid <= 8'h0;
    end else begin
      iacq_data_valid <= GEN_172;
    end
    if(reset) begin
      T_342 <= 3'h0;
    end else begin
      T_342 <= GEN_6;
    end
    if(reset) begin
      T_370 <= 3'h0;
    end else begin
      T_370 <= GEN_7;
    end
    if(reset) begin
      T_408 <= 3'h0;
    end else begin
      T_408 <= GEN_8;
    end
    if(reset) begin
      T_433 <= 3'h0;
    end else begin
      T_433 <= GEN_9;
    end
    if(reset) begin
      T_468 <= 3'h0;
    end else begin
      T_468 <= GEN_10;
    end
    if(reset) begin
      pending_ognt_ack <= 1'h0;
    end else begin
      pending_ognt_ack <= GEN_214;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fwrite(32'h80000002,"Assertion failed: Broadcast Hub does not support PutAtomics or prefetches\n    at broadcast.scala:203 assert(!(state =/= s_idle && xact.isBuiltInType() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_308) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different network source than initial request.\n    at broadcast.scala:285 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1152) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker accepted data beat from different client transaction than initial request.\n    at broadcast.scala:289 assert(!(state =/= s_idle && collect_iacq_data && io.inner.acquire.fire() &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1163) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fwrite(32'h80000002,"Assertion failed: AcquireTracker initialized with a tail data beat.\n    at broadcast.scala:293 assert(!(state === s_idle && io.inner.acquire.fire() && io.alloc.iacq &&\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1190) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module LockingRRArbiter_31(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input  [1:0] io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input  [1:0] io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  input  [1:0] io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  input  [1:0] io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [1:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_manager_xact_id,
  input   io_in_4_bits_is_builtin_type,
  input  [3:0] io_in_4_bits_g_type,
  input  [63:0] io_in_4_bits_data,
  input  [1:0] io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [1:0] io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_52;
  wire  GEN_8;
  wire [2:0] GEN_53;
  wire  GEN_9;
  wire [2:0] GEN_54;
  wire  GEN_10;
  wire  GEN_11;
  wire [2:0] GEN_1;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire [1:0] GEN_2;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire [2:0] GEN_3;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire  GEN_4;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [3:0] GEN_5;
  wire [3:0] GEN_28;
  wire [3:0] GEN_29;
  wire [3:0] GEN_30;
  wire [3:0] GEN_31;
  wire [63:0] GEN_6;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [1:0] GEN_7;
  wire [1:0] GEN_36;
  wire [1:0] GEN_37;
  wire [1:0] GEN_38;
  wire [1:0] GEN_39;
  reg [2:0] T_1228;
  reg [31:0] GEN_55;
  reg [2:0] T_1230;
  reg [31:0] GEN_56;
  wire [2:0] GEN_76;
  wire  T_1232;
  wire [2:0] T_1240_0;
  wire [3:0] GEN_77;
  wire  T_1242;
  wire [1:0] T_1250_0;
  wire [1:0] T_1250_1;
  wire [3:0] GEN_78;
  wire  T_1252;
  wire [3:0] GEN_79;
  wire  T_1253;
  wire  T_1256;
  wire  T_1257;
  wire  T_1259;
  wire  T_1260;
  wire [3:0] T_1264;
  wire [2:0] T_1265;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  reg [2:0] lastGrant;
  reg [31:0] GEN_57;
  wire [2:0] GEN_43;
  wire  T_1270;
  wire  T_1272;
  wire  T_1274;
  wire  T_1276;
  wire  T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire  T_1287;
  wire  T_1288;
  wire  T_1289;
  wire  T_1290;
  wire  T_1294;
  wire  T_1296;
  wire  T_1298;
  wire  T_1300;
  wire  T_1302;
  wire  T_1304;
  wire  T_1306;
  wire  T_1308;
  wire  T_1312;
  wire  T_1313;
  wire  T_1314;
  wire  T_1315;
  wire  T_1316;
  wire  T_1317;
  wire  T_1318;
  wire  T_1320;
  wire  T_1321;
  wire  T_1322;
  wire  T_1324;
  wire  T_1325;
  wire  T_1326;
  wire  T_1328;
  wire  T_1329;
  wire  T_1330;
  wire  T_1332;
  wire  T_1333;
  wire  T_1334;
  wire  T_1336;
  wire  T_1337;
  wire  T_1338;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  wire [2:0] GEN_48;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  assign io_in_0_ready = T_1322;
  assign io_in_1_ready = T_1326;
  assign io_in_2_ready = T_1330;
  assign io_in_3_ready = T_1334;
  assign io_in_4_ready = T_1338;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_42;
  assign choice = GEN_51;
  assign GEN_0 = GEN_11;
  assign GEN_52 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_52 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_53 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_53 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_54 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_54 == io_chosen ? io_in_3_valid : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_valid : GEN_10;
  assign GEN_1 = GEN_15;
  assign GEN_12 = GEN_52 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_13 = GEN_53 == io_chosen ? io_in_2_bits_addr_beat : GEN_12;
  assign GEN_14 = GEN_54 == io_chosen ? io_in_3_bits_addr_beat : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_14;
  assign GEN_2 = GEN_19;
  assign GEN_16 = GEN_52 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_17 = GEN_53 == io_chosen ? io_in_2_bits_client_xact_id : GEN_16;
  assign GEN_18 = GEN_54 == io_chosen ? io_in_3_bits_client_xact_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_18;
  assign GEN_3 = GEN_23;
  assign GEN_20 = GEN_52 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_21 = GEN_53 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_20;
  assign GEN_22 = GEN_54 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_21;
  assign GEN_23 = 3'h4 == io_chosen ? io_in_4_bits_manager_xact_id : GEN_22;
  assign GEN_4 = GEN_27;
  assign GEN_24 = GEN_52 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_25 = GEN_53 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_24;
  assign GEN_26 = GEN_54 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_25;
  assign GEN_27 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_26;
  assign GEN_5 = GEN_31;
  assign GEN_28 = GEN_52 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_29 = GEN_53 == io_chosen ? io_in_2_bits_g_type : GEN_28;
  assign GEN_30 = GEN_54 == io_chosen ? io_in_3_bits_g_type : GEN_29;
  assign GEN_31 = 3'h4 == io_chosen ? io_in_4_bits_g_type : GEN_30;
  assign GEN_6 = GEN_35;
  assign GEN_32 = GEN_52 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_33 = GEN_53 == io_chosen ? io_in_2_bits_data : GEN_32;
  assign GEN_34 = GEN_54 == io_chosen ? io_in_3_bits_data : GEN_33;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_34;
  assign GEN_7 = GEN_39;
  assign GEN_36 = GEN_52 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_37 = GEN_53 == io_chosen ? io_in_2_bits_client_id : GEN_36;
  assign GEN_38 = GEN_54 == io_chosen ? io_in_3_bits_client_id : GEN_37;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_38;
  assign GEN_76 = {{2'd0}, 1'h0};
  assign T_1232 = T_1228 != GEN_76;
  assign T_1240_0 = 3'h5;
  assign GEN_77 = {{1'd0}, T_1240_0};
  assign T_1242 = GEN_77 == io_out_bits_g_type;
  assign T_1250_0 = 2'h0;
  assign T_1250_1 = 2'h1;
  assign GEN_78 = {{2'd0}, T_1250_0};
  assign T_1252 = GEN_78 == io_out_bits_g_type;
  assign GEN_79 = {{2'd0}, T_1250_1};
  assign T_1253 = GEN_79 == io_out_bits_g_type;
  assign T_1256 = T_1252 | T_1253;
  assign T_1257 = io_out_bits_is_builtin_type ? T_1242 : T_1256;
  assign T_1259 = io_out_ready & io_out_valid;
  assign T_1260 = T_1259 & T_1257;
  assign T_1264 = T_1228 + GEN_52;
  assign T_1265 = T_1264[2:0];
  assign GEN_40 = T_1260 ? io_chosen : T_1230;
  assign GEN_41 = T_1260 ? T_1265 : T_1228;
  assign GEN_42 = T_1232 ? T_1230 : choice;
  assign GEN_43 = T_1259 ? io_chosen : lastGrant;
  assign T_1270 = GEN_52 > lastGrant;
  assign T_1272 = GEN_53 > lastGrant;
  assign T_1274 = GEN_54 > lastGrant;
  assign T_1276 = 3'h4 > lastGrant;
  assign T_1278 = io_in_1_valid & T_1270;
  assign T_1279 = io_in_2_valid & T_1272;
  assign T_1280 = io_in_3_valid & T_1274;
  assign T_1281 = io_in_4_valid & T_1276;
  assign T_1284 = T_1278 | T_1279;
  assign T_1285 = T_1284 | T_1280;
  assign T_1286 = T_1285 | T_1281;
  assign T_1287 = T_1286 | io_in_0_valid;
  assign T_1288 = T_1287 | io_in_1_valid;
  assign T_1289 = T_1288 | io_in_2_valid;
  assign T_1290 = T_1289 | io_in_3_valid;
  assign T_1294 = T_1278 == 1'h0;
  assign T_1296 = T_1284 == 1'h0;
  assign T_1298 = T_1285 == 1'h0;
  assign T_1300 = T_1286 == 1'h0;
  assign T_1302 = T_1287 == 1'h0;
  assign T_1304 = T_1288 == 1'h0;
  assign T_1306 = T_1289 == 1'h0;
  assign T_1308 = T_1290 == 1'h0;
  assign T_1312 = T_1270 | T_1302;
  assign T_1313 = T_1294 & T_1272;
  assign T_1314 = T_1313 | T_1304;
  assign T_1315 = T_1296 & T_1274;
  assign T_1316 = T_1315 | T_1306;
  assign T_1317 = T_1298 & T_1276;
  assign T_1318 = T_1317 | T_1308;
  assign T_1320 = T_1230 == GEN_76;
  assign T_1321 = T_1232 ? T_1320 : T_1300;
  assign T_1322 = T_1321 & io_out_ready;
  assign T_1324 = T_1230 == GEN_52;
  assign T_1325 = T_1232 ? T_1324 : T_1312;
  assign T_1326 = T_1325 & io_out_ready;
  assign T_1328 = T_1230 == GEN_53;
  assign T_1329 = T_1232 ? T_1328 : T_1314;
  assign T_1330 = T_1329 & io_out_ready;
  assign T_1332 = T_1230 == GEN_54;
  assign T_1333 = T_1232 ? T_1332 : T_1316;
  assign T_1334 = T_1333 & io_out_ready;
  assign T_1336 = T_1230 == 3'h4;
  assign T_1337 = T_1232 ? T_1336 : T_1318;
  assign T_1338 = T_1337 & io_out_ready;
  assign GEN_44 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_45 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_45;
  assign GEN_47 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_46;
  assign GEN_48 = T_1281 ? 3'h4 : GEN_47;
  assign GEN_49 = T_1280 ? {{1'd0}, 2'h3} : GEN_48;
  assign GEN_50 = T_1279 ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = T_1278 ? {{2'd0}, 1'h1} : GEN_50;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_55 = {1{$random}};
  T_1228 = GEN_55[2:0];
  GEN_56 = {1{$random}};
  T_1230 = GEN_56[2:0];
  GEN_57 = {1{$random}};
  lastGrant = GEN_57[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1228 <= 3'h0;
    end else begin
      T_1228 <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      T_1230 <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_43;
    end
  end
endmodule
module LockingRRArbiter_32(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_p_type,
  input  [1:0] io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_p_type,
  input  [1:0] io_in_1_bits_client_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_p_type,
  input  [1:0] io_in_2_bits_client_id,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [1:0] io_in_3_bits_p_type,
  input  [1:0] io_in_3_bits_client_id,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [1:0] io_in_4_bits_p_type,
  input  [1:0] io_in_4_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_p_type,
  output [1:0] io_out_bits_client_id,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_32;
  wire  GEN_4;
  wire [2:0] GEN_33;
  wire  GEN_5;
  wire [2:0] GEN_34;
  wire  GEN_6;
  wire  GEN_7;
  wire [25:0] GEN_1;
  wire [25:0] GEN_8;
  wire [25:0] GEN_9;
  wire [25:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_2;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_3;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  reg [2:0] T_1076;
  reg [31:0] GEN_20;
  reg [2:0] T_1078;
  reg [31:0] GEN_21;
  wire [2:0] GEN_44;
  wire  T_1080;
  wire  T_1082;
  wire [2:0] GEN_22;
  reg [2:0] lastGrant;
  reg [31:0] GEN_35;
  wire [2:0] GEN_23;
  wire  T_1093;
  wire  T_1095;
  wire  T_1097;
  wire  T_1099;
  wire  T_1101;
  wire  T_1102;
  wire  T_1103;
  wire  T_1104;
  wire  T_1107;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire  T_1112;
  wire  T_1113;
  wire  T_1117;
  wire  T_1119;
  wire  T_1121;
  wire  T_1123;
  wire  T_1125;
  wire  T_1127;
  wire  T_1129;
  wire  T_1131;
  wire  T_1135;
  wire  T_1136;
  wire  T_1137;
  wire  T_1138;
  wire  T_1139;
  wire  T_1140;
  wire  T_1141;
  wire  T_1143;
  wire  T_1144;
  wire  T_1145;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1151;
  wire  T_1152;
  wire  T_1153;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1159;
  wire  T_1160;
  wire  T_1161;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire [2:0] GEN_27;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  assign io_in_0_ready = T_1145;
  assign io_in_1_ready = T_1149;
  assign io_in_2_ready = T_1153;
  assign io_in_3_ready = T_1157;
  assign io_in_4_ready = T_1161;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_p_type = GEN_2;
  assign io_out_bits_client_id = GEN_3;
  assign io_chosen = GEN_22;
  assign choice = GEN_31;
  assign GEN_0 = GEN_7;
  assign GEN_32 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_32 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_33 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_33 == io_chosen ? io_in_2_valid : GEN_4;
  assign GEN_34 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_34 == io_chosen ? io_in_3_valid : GEN_5;
  assign GEN_7 = 3'h4 == io_chosen ? io_in_4_valid : GEN_6;
  assign GEN_1 = GEN_11;
  assign GEN_8 = GEN_32 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_9 = GEN_33 == io_chosen ? io_in_2_bits_addr_block : GEN_8;
  assign GEN_10 = GEN_34 == io_chosen ? io_in_3_bits_addr_block : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_10;
  assign GEN_2 = GEN_15;
  assign GEN_12 = GEN_32 == io_chosen ? io_in_1_bits_p_type : io_in_0_bits_p_type;
  assign GEN_13 = GEN_33 == io_chosen ? io_in_2_bits_p_type : GEN_12;
  assign GEN_14 = GEN_34 == io_chosen ? io_in_3_bits_p_type : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_p_type : GEN_14;
  assign GEN_3 = GEN_19;
  assign GEN_16 = GEN_32 == io_chosen ? io_in_1_bits_client_id : io_in_0_bits_client_id;
  assign GEN_17 = GEN_33 == io_chosen ? io_in_2_bits_client_id : GEN_16;
  assign GEN_18 = GEN_34 == io_chosen ? io_in_3_bits_client_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_id : GEN_18;
  assign GEN_44 = {{2'd0}, 1'h0};
  assign T_1080 = T_1076 != GEN_44;
  assign T_1082 = io_out_ready & io_out_valid;
  assign GEN_22 = T_1080 ? T_1078 : choice;
  assign GEN_23 = T_1082 ? io_chosen : lastGrant;
  assign T_1093 = GEN_32 > lastGrant;
  assign T_1095 = GEN_33 > lastGrant;
  assign T_1097 = GEN_34 > lastGrant;
  assign T_1099 = 3'h4 > lastGrant;
  assign T_1101 = io_in_1_valid & T_1093;
  assign T_1102 = io_in_2_valid & T_1095;
  assign T_1103 = io_in_3_valid & T_1097;
  assign T_1104 = io_in_4_valid & T_1099;
  assign T_1107 = T_1101 | T_1102;
  assign T_1108 = T_1107 | T_1103;
  assign T_1109 = T_1108 | T_1104;
  assign T_1110 = T_1109 | io_in_0_valid;
  assign T_1111 = T_1110 | io_in_1_valid;
  assign T_1112 = T_1111 | io_in_2_valid;
  assign T_1113 = T_1112 | io_in_3_valid;
  assign T_1117 = T_1101 == 1'h0;
  assign T_1119 = T_1107 == 1'h0;
  assign T_1121 = T_1108 == 1'h0;
  assign T_1123 = T_1109 == 1'h0;
  assign T_1125 = T_1110 == 1'h0;
  assign T_1127 = T_1111 == 1'h0;
  assign T_1129 = T_1112 == 1'h0;
  assign T_1131 = T_1113 == 1'h0;
  assign T_1135 = T_1093 | T_1125;
  assign T_1136 = T_1117 & T_1095;
  assign T_1137 = T_1136 | T_1127;
  assign T_1138 = T_1119 & T_1097;
  assign T_1139 = T_1138 | T_1129;
  assign T_1140 = T_1121 & T_1099;
  assign T_1141 = T_1140 | T_1131;
  assign T_1143 = T_1078 == GEN_44;
  assign T_1144 = T_1080 ? T_1143 : T_1123;
  assign T_1145 = T_1144 & io_out_ready;
  assign T_1147 = T_1078 == GEN_32;
  assign T_1148 = T_1080 ? T_1147 : T_1135;
  assign T_1149 = T_1148 & io_out_ready;
  assign T_1151 = T_1078 == GEN_33;
  assign T_1152 = T_1080 ? T_1151 : T_1137;
  assign T_1153 = T_1152 & io_out_ready;
  assign T_1155 = T_1078 == GEN_34;
  assign T_1156 = T_1080 ? T_1155 : T_1139;
  assign T_1157 = T_1156 & io_out_ready;
  assign T_1159 = T_1078 == 3'h4;
  assign T_1160 = T_1080 ? T_1159 : T_1141;
  assign T_1161 = T_1160 & io_out_ready;
  assign GEN_24 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_25 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_24;
  assign GEN_26 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_25;
  assign GEN_27 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_26;
  assign GEN_28 = T_1104 ? 3'h4 : GEN_27;
  assign GEN_29 = T_1103 ? {{1'd0}, 2'h3} : GEN_28;
  assign GEN_30 = T_1102 ? {{1'd0}, 2'h2} : GEN_29;
  assign GEN_31 = T_1101 ? {{2'd0}, 1'h1} : GEN_30;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  T_1076 = GEN_20[2:0];
  GEN_21 = {1{$random}};
  T_1078 = GEN_21[2:0];
  GEN_35 = {1{$random}};
  lastGrant = GEN_35[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_1076 <= 3'h0;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_23;
    end
  end
endmodule
module LockingRRArbiter_33(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [4:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [4:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [2:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [11:0] io_in_2_bits_union,
  input  [4:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [25:0] io_in_3_bits_addr_block,
  input  [2:0] io_in_3_bits_client_xact_id,
  input  [2:0] io_in_3_bits_addr_beat,
  input   io_in_3_bits_is_builtin_type,
  input  [2:0] io_in_3_bits_a_type,
  input  [11:0] io_in_3_bits_union,
  input  [4:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [25:0] io_in_4_bits_addr_block,
  input  [2:0] io_in_4_bits_client_xact_id,
  input  [2:0] io_in_4_bits_addr_beat,
  input   io_in_4_bits_is_builtin_type,
  input  [2:0] io_in_4_bits_a_type,
  input  [11:0] io_in_4_bits_union,
  input  [4:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [4:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_52;
  wire  GEN_8;
  wire [2:0] GEN_53;
  wire  GEN_9;
  wire [2:0] GEN_54;
  wire  GEN_10;
  wire  GEN_11;
  wire [25:0] GEN_1;
  wire [25:0] GEN_12;
  wire [25:0] GEN_13;
  wire [25:0] GEN_14;
  wire [25:0] GEN_15;
  wire [2:0] GEN_2;
  wire [2:0] GEN_16;
  wire [2:0] GEN_17;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [2:0] GEN_3;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire  GEN_4;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [2:0] GEN_5;
  wire [2:0] GEN_28;
  wire [2:0] GEN_29;
  wire [2:0] GEN_30;
  wire [2:0] GEN_31;
  wire [11:0] GEN_6;
  wire [11:0] GEN_32;
  wire [11:0] GEN_33;
  wire [11:0] GEN_34;
  wire [11:0] GEN_35;
  wire [4:0] GEN_7;
  wire [4:0] GEN_36;
  wire [4:0] GEN_37;
  wire [4:0] GEN_38;
  wire [4:0] GEN_39;
  reg [2:0] T_354;
  reg [31:0] GEN_55;
  reg [2:0] T_356;
  reg [31:0] GEN_56;
  wire [2:0] GEN_76;
  wire  T_358;
  wire [2:0] T_367_0;
  wire  T_369;
  wire  T_372;
  wire  T_373;
  wire  T_374;
  wire [3:0] T_378;
  wire [2:0] T_379;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  reg [2:0] lastGrant;
  reg [31:0] GEN_57;
  wire [2:0] GEN_43;
  wire  T_384;
  wire  T_386;
  wire  T_388;
  wire  T_390;
  wire  T_392;
  wire  T_393;
  wire  T_394;
  wire  T_395;
  wire  T_398;
  wire  T_399;
  wire  T_400;
  wire  T_401;
  wire  T_402;
  wire  T_403;
  wire  T_404;
  wire  T_408;
  wire  T_410;
  wire  T_412;
  wire  T_414;
  wire  T_416;
  wire  T_418;
  wire  T_420;
  wire  T_422;
  wire  T_426;
  wire  T_427;
  wire  T_428;
  wire  T_429;
  wire  T_430;
  wire  T_431;
  wire  T_432;
  wire  T_434;
  wire  T_435;
  wire  T_436;
  wire  T_438;
  wire  T_439;
  wire  T_440;
  wire  T_442;
  wire  T_443;
  wire  T_444;
  wire  T_446;
  wire  T_447;
  wire  T_448;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  wire [2:0] GEN_48;
  wire [2:0] GEN_49;
  wire [2:0] GEN_50;
  wire [2:0] GEN_51;
  assign io_in_0_ready = T_436;
  assign io_in_1_ready = T_440;
  assign io_in_2_ready = T_444;
  assign io_in_3_ready = T_448;
  assign io_in_4_ready = T_452;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_42;
  assign choice = GEN_51;
  assign GEN_0 = GEN_11;
  assign GEN_52 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_52 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_53 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_53 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_54 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_54 == io_chosen ? io_in_3_valid : GEN_9;
  assign GEN_11 = 3'h4 == io_chosen ? io_in_4_valid : GEN_10;
  assign GEN_1 = GEN_15;
  assign GEN_12 = GEN_52 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_13 = GEN_53 == io_chosen ? io_in_2_bits_addr_block : GEN_12;
  assign GEN_14 = GEN_54 == io_chosen ? io_in_3_bits_addr_block : GEN_13;
  assign GEN_15 = 3'h4 == io_chosen ? io_in_4_bits_addr_block : GEN_14;
  assign GEN_2 = GEN_19;
  assign GEN_16 = GEN_52 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_17 = GEN_53 == io_chosen ? io_in_2_bits_client_xact_id : GEN_16;
  assign GEN_18 = GEN_54 == io_chosen ? io_in_3_bits_client_xact_id : GEN_17;
  assign GEN_19 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_18;
  assign GEN_3 = GEN_23;
  assign GEN_20 = GEN_52 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_21 = GEN_53 == io_chosen ? io_in_2_bits_addr_beat : GEN_20;
  assign GEN_22 = GEN_54 == io_chosen ? io_in_3_bits_addr_beat : GEN_21;
  assign GEN_23 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_22;
  assign GEN_4 = GEN_27;
  assign GEN_24 = GEN_52 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_25 = GEN_53 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_24;
  assign GEN_26 = GEN_54 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_25;
  assign GEN_27 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_26;
  assign GEN_5 = GEN_31;
  assign GEN_28 = GEN_52 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_29 = GEN_53 == io_chosen ? io_in_2_bits_a_type : GEN_28;
  assign GEN_30 = GEN_54 == io_chosen ? io_in_3_bits_a_type : GEN_29;
  assign GEN_31 = 3'h4 == io_chosen ? io_in_4_bits_a_type : GEN_30;
  assign GEN_6 = GEN_35;
  assign GEN_32 = GEN_52 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_33 = GEN_53 == io_chosen ? io_in_2_bits_union : GEN_32;
  assign GEN_34 = GEN_54 == io_chosen ? io_in_3_bits_union : GEN_33;
  assign GEN_35 = 3'h4 == io_chosen ? io_in_4_bits_union : GEN_34;
  assign GEN_7 = GEN_39;
  assign GEN_36 = GEN_52 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_37 = GEN_53 == io_chosen ? io_in_2_bits_data : GEN_36;
  assign GEN_38 = GEN_54 == io_chosen ? io_in_3_bits_data : GEN_37;
  assign GEN_39 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_38;
  assign GEN_76 = {{2'd0}, 1'h0};
  assign T_358 = T_354 != GEN_76;
  assign T_367_0 = 3'h3;
  assign T_369 = T_367_0 == io_out_bits_a_type;
  assign T_372 = io_out_bits_is_builtin_type & T_369;
  assign T_373 = io_out_ready & io_out_valid;
  assign T_374 = T_373 & T_372;
  assign T_378 = T_354 + GEN_52;
  assign T_379 = T_378[2:0];
  assign GEN_40 = T_374 ? io_chosen : T_356;
  assign GEN_41 = T_374 ? T_379 : T_354;
  assign GEN_42 = T_358 ? T_356 : choice;
  assign GEN_43 = T_373 ? io_chosen : lastGrant;
  assign T_384 = GEN_52 > lastGrant;
  assign T_386 = GEN_53 > lastGrant;
  assign T_388 = GEN_54 > lastGrant;
  assign T_390 = 3'h4 > lastGrant;
  assign T_392 = io_in_1_valid & T_384;
  assign T_393 = io_in_2_valid & T_386;
  assign T_394 = io_in_3_valid & T_388;
  assign T_395 = io_in_4_valid & T_390;
  assign T_398 = T_392 | T_393;
  assign T_399 = T_398 | T_394;
  assign T_400 = T_399 | T_395;
  assign T_401 = T_400 | io_in_0_valid;
  assign T_402 = T_401 | io_in_1_valid;
  assign T_403 = T_402 | io_in_2_valid;
  assign T_404 = T_403 | io_in_3_valid;
  assign T_408 = T_392 == 1'h0;
  assign T_410 = T_398 == 1'h0;
  assign T_412 = T_399 == 1'h0;
  assign T_414 = T_400 == 1'h0;
  assign T_416 = T_401 == 1'h0;
  assign T_418 = T_402 == 1'h0;
  assign T_420 = T_403 == 1'h0;
  assign T_422 = T_404 == 1'h0;
  assign T_426 = T_384 | T_416;
  assign T_427 = T_408 & T_386;
  assign T_428 = T_427 | T_418;
  assign T_429 = T_410 & T_388;
  assign T_430 = T_429 | T_420;
  assign T_431 = T_412 & T_390;
  assign T_432 = T_431 | T_422;
  assign T_434 = T_356 == GEN_76;
  assign T_435 = T_358 ? T_434 : T_414;
  assign T_436 = T_435 & io_out_ready;
  assign T_438 = T_356 == GEN_52;
  assign T_439 = T_358 ? T_438 : T_426;
  assign T_440 = T_439 & io_out_ready;
  assign T_442 = T_356 == GEN_53;
  assign T_443 = T_358 ? T_442 : T_428;
  assign T_444 = T_443 & io_out_ready;
  assign T_446 = T_356 == GEN_54;
  assign T_447 = T_358 ? T_446 : T_430;
  assign T_448 = T_447 & io_out_ready;
  assign T_450 = T_356 == 3'h4;
  assign T_451 = T_358 ? T_450 : T_432;
  assign T_452 = T_451 & io_out_ready;
  assign GEN_44 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_45 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_45;
  assign GEN_47 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_46;
  assign GEN_48 = T_395 ? 3'h4 : GEN_47;
  assign GEN_49 = T_394 ? {{1'd0}, 2'h3} : GEN_48;
  assign GEN_50 = T_393 ? {{1'd0}, 2'h2} : GEN_49;
  assign GEN_51 = T_392 ? {{2'd0}, 1'h1} : GEN_50;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_55 = {1{$random}};
  T_354 = GEN_55[2:0];
  GEN_56 = {1{$random}};
  T_356 = GEN_56[2:0];
  GEN_57 = {1{$random}};
  lastGrant = GEN_57[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_354 <= 3'h0;
    end else begin
      T_354 <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      T_356 <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_43;
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [4:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [4:0] io_in_0_grant_bits_data,
  output  io_in_1_acquire_ready,
  input   io_in_1_acquire_valid,
  input  [25:0] io_in_1_acquire_bits_addr_block,
  input  [2:0] io_in_1_acquire_bits_client_xact_id,
  input  [2:0] io_in_1_acquire_bits_addr_beat,
  input   io_in_1_acquire_bits_is_builtin_type,
  input  [2:0] io_in_1_acquire_bits_a_type,
  input  [11:0] io_in_1_acquire_bits_union,
  input  [4:0] io_in_1_acquire_bits_data,
  input   io_in_1_grant_ready,
  output  io_in_1_grant_valid,
  output [2:0] io_in_1_grant_bits_addr_beat,
  output [2:0] io_in_1_grant_bits_client_xact_id,
  output  io_in_1_grant_bits_manager_xact_id,
  output  io_in_1_grant_bits_is_builtin_type,
  output [3:0] io_in_1_grant_bits_g_type,
  output [4:0] io_in_1_grant_bits_data,
  output  io_in_2_acquire_ready,
  input   io_in_2_acquire_valid,
  input  [25:0] io_in_2_acquire_bits_addr_block,
  input  [2:0] io_in_2_acquire_bits_client_xact_id,
  input  [2:0] io_in_2_acquire_bits_addr_beat,
  input   io_in_2_acquire_bits_is_builtin_type,
  input  [2:0] io_in_2_acquire_bits_a_type,
  input  [11:0] io_in_2_acquire_bits_union,
  input  [4:0] io_in_2_acquire_bits_data,
  input   io_in_2_grant_ready,
  output  io_in_2_grant_valid,
  output [2:0] io_in_2_grant_bits_addr_beat,
  output [2:0] io_in_2_grant_bits_client_xact_id,
  output  io_in_2_grant_bits_manager_xact_id,
  output  io_in_2_grant_bits_is_builtin_type,
  output [3:0] io_in_2_grant_bits_g_type,
  output [4:0] io_in_2_grant_bits_data,
  output  io_in_3_acquire_ready,
  input   io_in_3_acquire_valid,
  input  [25:0] io_in_3_acquire_bits_addr_block,
  input  [2:0] io_in_3_acquire_bits_client_xact_id,
  input  [2:0] io_in_3_acquire_bits_addr_beat,
  input   io_in_3_acquire_bits_is_builtin_type,
  input  [2:0] io_in_3_acquire_bits_a_type,
  input  [11:0] io_in_3_acquire_bits_union,
  input  [4:0] io_in_3_acquire_bits_data,
  input   io_in_3_grant_ready,
  output  io_in_3_grant_valid,
  output [2:0] io_in_3_grant_bits_addr_beat,
  output [2:0] io_in_3_grant_bits_client_xact_id,
  output  io_in_3_grant_bits_manager_xact_id,
  output  io_in_3_grant_bits_is_builtin_type,
  output [3:0] io_in_3_grant_bits_g_type,
  output [4:0] io_in_3_grant_bits_data,
  output  io_in_4_acquire_ready,
  input   io_in_4_acquire_valid,
  input  [25:0] io_in_4_acquire_bits_addr_block,
  input  [2:0] io_in_4_acquire_bits_client_xact_id,
  input  [2:0] io_in_4_acquire_bits_addr_beat,
  input   io_in_4_acquire_bits_is_builtin_type,
  input  [2:0] io_in_4_acquire_bits_a_type,
  input  [11:0] io_in_4_acquire_bits_union,
  input  [4:0] io_in_4_acquire_bits_data,
  input   io_in_4_grant_ready,
  output  io_in_4_grant_valid,
  output [2:0] io_in_4_grant_bits_addr_beat,
  output [2:0] io_in_4_grant_bits_client_xact_id,
  output  io_in_4_grant_bits_manager_xact_id,
  output  io_in_4_grant_bits_is_builtin_type,
  output [3:0] io_in_4_grant_bits_g_type,
  output [4:0] io_in_4_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [4:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [4:0] io_out_grant_bits_data
);
  wire  LockingRRArbiter_33_1165_clk;
  wire  LockingRRArbiter_33_1165_reset;
  wire  LockingRRArbiter_33_1165_io_in_0_ready;
  wire  LockingRRArbiter_33_1165_io_in_0_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_in_0_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_in_0_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_in_0_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_in_0_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_in_0_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_in_0_bits_data;
  wire  LockingRRArbiter_33_1165_io_in_1_ready;
  wire  LockingRRArbiter_33_1165_io_in_1_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_in_1_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_in_1_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_in_1_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_in_1_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_in_1_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_in_1_bits_data;
  wire  LockingRRArbiter_33_1165_io_in_2_ready;
  wire  LockingRRArbiter_33_1165_io_in_2_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_in_2_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_in_2_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_in_2_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_in_2_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_in_2_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_in_2_bits_data;
  wire  LockingRRArbiter_33_1165_io_in_3_ready;
  wire  LockingRRArbiter_33_1165_io_in_3_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_in_3_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_in_3_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_in_3_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_in_3_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_in_3_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_in_3_bits_data;
  wire  LockingRRArbiter_33_1165_io_in_4_ready;
  wire  LockingRRArbiter_33_1165_io_in_4_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_in_4_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_in_4_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_in_4_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_in_4_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_in_4_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_in_4_bits_data;
  wire  LockingRRArbiter_33_1165_io_out_ready;
  wire  LockingRRArbiter_33_1165_io_out_valid;
  wire [25:0] LockingRRArbiter_33_1165_io_out_bits_addr_block;
  wire [2:0] LockingRRArbiter_33_1165_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_33_1165_io_out_bits_addr_beat;
  wire  LockingRRArbiter_33_1165_io_out_bits_is_builtin_type;
  wire [2:0] LockingRRArbiter_33_1165_io_out_bits_a_type;
  wire [11:0] LockingRRArbiter_33_1165_io_out_bits_union;
  wire [4:0] LockingRRArbiter_33_1165_io_out_bits_data;
  wire [2:0] LockingRRArbiter_33_1165_io_chosen;
  wire [5:0] T_1167;
  wire [5:0] T_1169;
  wire [5:0] T_1171;
  wire [5:0] T_1173;
  wire [5:0] T_1175;
  wire [2:0] GEN_10;
  wire  T_1180;
  wire  GEN_0;
  wire  GEN_1;
  wire [2:0] GEN_11;
  wire  T_1185;
  wire  GEN_2;
  wire  GEN_3;
  wire [2:0] GEN_12;
  wire  T_1190;
  wire  GEN_4;
  wire  GEN_5;
  wire [2:0] GEN_13;
  wire  T_1195;
  wire  GEN_6;
  wire  GEN_7;
  wire  T_1200;
  wire  GEN_8;
  wire  GEN_9;
  LockingRRArbiter_33 LockingRRArbiter_33_1165 (
    .clk(LockingRRArbiter_33_1165_clk),
    .reset(LockingRRArbiter_33_1165_reset),
    .io_in_0_ready(LockingRRArbiter_33_1165_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_33_1165_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_33_1165_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_33_1165_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(LockingRRArbiter_33_1165_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_33_1165_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(LockingRRArbiter_33_1165_io_in_0_bits_a_type),
    .io_in_0_bits_union(LockingRRArbiter_33_1165_io_in_0_bits_union),
    .io_in_0_bits_data(LockingRRArbiter_33_1165_io_in_0_bits_data),
    .io_in_1_ready(LockingRRArbiter_33_1165_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_33_1165_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_33_1165_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_33_1165_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(LockingRRArbiter_33_1165_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_33_1165_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(LockingRRArbiter_33_1165_io_in_1_bits_a_type),
    .io_in_1_bits_union(LockingRRArbiter_33_1165_io_in_1_bits_union),
    .io_in_1_bits_data(LockingRRArbiter_33_1165_io_in_1_bits_data),
    .io_in_2_ready(LockingRRArbiter_33_1165_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_33_1165_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_33_1165_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_33_1165_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(LockingRRArbiter_33_1165_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_33_1165_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(LockingRRArbiter_33_1165_io_in_2_bits_a_type),
    .io_in_2_bits_union(LockingRRArbiter_33_1165_io_in_2_bits_union),
    .io_in_2_bits_data(LockingRRArbiter_33_1165_io_in_2_bits_data),
    .io_in_3_ready(LockingRRArbiter_33_1165_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_33_1165_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_33_1165_io_in_3_bits_addr_block),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_33_1165_io_in_3_bits_client_xact_id),
    .io_in_3_bits_addr_beat(LockingRRArbiter_33_1165_io_in_3_bits_addr_beat),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_33_1165_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_a_type(LockingRRArbiter_33_1165_io_in_3_bits_a_type),
    .io_in_3_bits_union(LockingRRArbiter_33_1165_io_in_3_bits_union),
    .io_in_3_bits_data(LockingRRArbiter_33_1165_io_in_3_bits_data),
    .io_in_4_ready(LockingRRArbiter_33_1165_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_33_1165_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_33_1165_io_in_4_bits_addr_block),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_33_1165_io_in_4_bits_client_xact_id),
    .io_in_4_bits_addr_beat(LockingRRArbiter_33_1165_io_in_4_bits_addr_beat),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_33_1165_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_a_type(LockingRRArbiter_33_1165_io_in_4_bits_a_type),
    .io_in_4_bits_union(LockingRRArbiter_33_1165_io_in_4_bits_union),
    .io_in_4_bits_data(LockingRRArbiter_33_1165_io_in_4_bits_data),
    .io_out_ready(LockingRRArbiter_33_1165_io_out_ready),
    .io_out_valid(LockingRRArbiter_33_1165_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_33_1165_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(LockingRRArbiter_33_1165_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(LockingRRArbiter_33_1165_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(LockingRRArbiter_33_1165_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(LockingRRArbiter_33_1165_io_out_bits_a_type),
    .io_out_bits_union(LockingRRArbiter_33_1165_io_out_bits_union),
    .io_out_bits_data(LockingRRArbiter_33_1165_io_out_bits_data),
    .io_chosen(LockingRRArbiter_33_1165_io_chosen)
  );
  assign io_in_0_acquire_ready = LockingRRArbiter_33_1165_io_in_0_ready;
  assign io_in_0_grant_valid = GEN_0;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_in_1_acquire_ready = LockingRRArbiter_33_1165_io_in_1_ready;
  assign io_in_1_grant_valid = GEN_2;
  assign io_in_1_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_1_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_1_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_1_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_1_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_1_grant_bits_data = io_out_grant_bits_data;
  assign io_in_2_acquire_ready = LockingRRArbiter_33_1165_io_in_2_ready;
  assign io_in_2_grant_valid = GEN_4;
  assign io_in_2_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_2_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_2_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_2_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_2_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_2_grant_bits_data = io_out_grant_bits_data;
  assign io_in_3_acquire_ready = LockingRRArbiter_33_1165_io_in_3_ready;
  assign io_in_3_grant_valid = GEN_6;
  assign io_in_3_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_3_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_3_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_3_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_3_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_3_grant_bits_data = io_out_grant_bits_data;
  assign io_in_4_acquire_ready = LockingRRArbiter_33_1165_io_in_4_ready;
  assign io_in_4_grant_valid = GEN_8;
  assign io_in_4_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_4_grant_bits_client_xact_id = {{2'd0}, 1'h0};
  assign io_in_4_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_4_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_4_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_4_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = LockingRRArbiter_33_1165_io_out_valid;
  assign io_out_acquire_bits_addr_block = LockingRRArbiter_33_1165_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = LockingRRArbiter_33_1165_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = LockingRRArbiter_33_1165_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = LockingRRArbiter_33_1165_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = LockingRRArbiter_33_1165_io_out_bits_a_type;
  assign io_out_acquire_bits_union = LockingRRArbiter_33_1165_io_out_bits_union;
  assign io_out_acquire_bits_data = LockingRRArbiter_33_1165_io_out_bits_data;
  assign io_out_grant_ready = GEN_9;
  assign LockingRRArbiter_33_1165_clk = clk;
  assign LockingRRArbiter_33_1165_reset = reset;
  assign LockingRRArbiter_33_1165_io_in_0_valid = io_in_0_acquire_valid;
  assign LockingRRArbiter_33_1165_io_in_0_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign LockingRRArbiter_33_1165_io_in_0_bits_client_xact_id = T_1167[2:0];
  assign LockingRRArbiter_33_1165_io_in_0_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign LockingRRArbiter_33_1165_io_in_0_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_33_1165_io_in_0_bits_a_type = io_in_0_acquire_bits_a_type;
  assign LockingRRArbiter_33_1165_io_in_0_bits_union = io_in_0_acquire_bits_union;
  assign LockingRRArbiter_33_1165_io_in_0_bits_data = io_in_0_acquire_bits_data;
  assign LockingRRArbiter_33_1165_io_in_1_valid = io_in_1_acquire_valid;
  assign LockingRRArbiter_33_1165_io_in_1_bits_addr_block = io_in_1_acquire_bits_addr_block;
  assign LockingRRArbiter_33_1165_io_in_1_bits_client_xact_id = T_1169[2:0];
  assign LockingRRArbiter_33_1165_io_in_1_bits_addr_beat = io_in_1_acquire_bits_addr_beat;
  assign LockingRRArbiter_33_1165_io_in_1_bits_is_builtin_type = io_in_1_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_33_1165_io_in_1_bits_a_type = io_in_1_acquire_bits_a_type;
  assign LockingRRArbiter_33_1165_io_in_1_bits_union = io_in_1_acquire_bits_union;
  assign LockingRRArbiter_33_1165_io_in_1_bits_data = io_in_1_acquire_bits_data;
  assign LockingRRArbiter_33_1165_io_in_2_valid = io_in_2_acquire_valid;
  assign LockingRRArbiter_33_1165_io_in_2_bits_addr_block = io_in_2_acquire_bits_addr_block;
  assign LockingRRArbiter_33_1165_io_in_2_bits_client_xact_id = T_1171[2:0];
  assign LockingRRArbiter_33_1165_io_in_2_bits_addr_beat = io_in_2_acquire_bits_addr_beat;
  assign LockingRRArbiter_33_1165_io_in_2_bits_is_builtin_type = io_in_2_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_33_1165_io_in_2_bits_a_type = io_in_2_acquire_bits_a_type;
  assign LockingRRArbiter_33_1165_io_in_2_bits_union = io_in_2_acquire_bits_union;
  assign LockingRRArbiter_33_1165_io_in_2_bits_data = io_in_2_acquire_bits_data;
  assign LockingRRArbiter_33_1165_io_in_3_valid = io_in_3_acquire_valid;
  assign LockingRRArbiter_33_1165_io_in_3_bits_addr_block = io_in_3_acquire_bits_addr_block;
  assign LockingRRArbiter_33_1165_io_in_3_bits_client_xact_id = T_1173[2:0];
  assign LockingRRArbiter_33_1165_io_in_3_bits_addr_beat = io_in_3_acquire_bits_addr_beat;
  assign LockingRRArbiter_33_1165_io_in_3_bits_is_builtin_type = io_in_3_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_33_1165_io_in_3_bits_a_type = io_in_3_acquire_bits_a_type;
  assign LockingRRArbiter_33_1165_io_in_3_bits_union = io_in_3_acquire_bits_union;
  assign LockingRRArbiter_33_1165_io_in_3_bits_data = io_in_3_acquire_bits_data;
  assign LockingRRArbiter_33_1165_io_in_4_valid = io_in_4_acquire_valid;
  assign LockingRRArbiter_33_1165_io_in_4_bits_addr_block = io_in_4_acquire_bits_addr_block;
  assign LockingRRArbiter_33_1165_io_in_4_bits_client_xact_id = T_1175[2:0];
  assign LockingRRArbiter_33_1165_io_in_4_bits_addr_beat = io_in_4_acquire_bits_addr_beat;
  assign LockingRRArbiter_33_1165_io_in_4_bits_is_builtin_type = io_in_4_acquire_bits_is_builtin_type;
  assign LockingRRArbiter_33_1165_io_in_4_bits_a_type = io_in_4_acquire_bits_a_type;
  assign LockingRRArbiter_33_1165_io_in_4_bits_union = io_in_4_acquire_bits_union;
  assign LockingRRArbiter_33_1165_io_in_4_bits_data = io_in_4_acquire_bits_data;
  assign LockingRRArbiter_33_1165_io_out_ready = io_out_acquire_ready;
  assign T_1167 = {io_in_0_acquire_bits_client_xact_id,3'h0};
  assign T_1169 = {io_in_1_acquire_bits_client_xact_id,3'h1};
  assign T_1171 = {io_in_2_acquire_bits_client_xact_id,3'h2};
  assign T_1173 = {io_in_3_acquire_bits_client_xact_id,3'h3};
  assign T_1175 = {io_in_4_acquire_bits_client_xact_id,3'h4};
  assign GEN_10 = {{2'd0}, 1'h0};
  assign T_1180 = io_out_grant_bits_client_xact_id == GEN_10;
  assign GEN_0 = T_1180 ? io_out_grant_valid : 1'h0;
  assign GEN_1 = T_1180 ? io_in_0_grant_ready : 1'h0;
  assign GEN_11 = {{2'd0}, 1'h1};
  assign T_1185 = io_out_grant_bits_client_xact_id == GEN_11;
  assign GEN_2 = T_1185 ? io_out_grant_valid : 1'h0;
  assign GEN_3 = T_1185 ? io_in_1_grant_ready : GEN_1;
  assign GEN_12 = {{1'd0}, 2'h2};
  assign T_1190 = io_out_grant_bits_client_xact_id == GEN_12;
  assign GEN_4 = T_1190 ? io_out_grant_valid : 1'h0;
  assign GEN_5 = T_1190 ? io_in_2_grant_ready : GEN_3;
  assign GEN_13 = {{1'd0}, 2'h3};
  assign T_1195 = io_out_grant_bits_client_xact_id == GEN_13;
  assign GEN_6 = T_1195 ? io_out_grant_valid : 1'h0;
  assign GEN_7 = T_1195 ? io_in_3_grant_ready : GEN_5;
  assign T_1200 = io_out_grant_bits_client_xact_id == 3'h4;
  assign GEN_8 = T_1200 ? io_out_grant_valid : 1'h0;
  assign GEN_9 = T_1200 ? io_in_4_grant_ready : GEN_7;
endmodule
module L2BroadcastHub(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  BroadcastVoluntaryReleaseTracker_1051_clk;
  wire  BroadcastVoluntaryReleaseTracker_1051_reset;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_valid;
  wire [25:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_block;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_beat;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type;
  wire [11:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_union;
  wire [4:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_data;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_valid;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_addr_beat;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_xact_id;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_manager_xact_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_g_type;
  wire [4:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_data;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_valid;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_bits_manager_xact_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_valid;
  wire [25:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_addr_block;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_p_type;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_client_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_release_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_release_valid;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_beat;
  wire [25:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_block;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_xact_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_voluntary;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_r_type;
  wire [4:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_data;
  wire [1:0] BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_incoherent_0;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_valid;
  wire [25:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_block;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_beat;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_a_type;
  wire [11:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_union;
  wire [4:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_data;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_ready;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_valid;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_addr_beat;
  wire [2:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_client_xact_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_manager_xact_id;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_g_type;
  wire [4:0] BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_data;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_matches_iacq;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_matches_irel;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_matches_oprb;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_alloc_iacq;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_alloc_irel;
  wire  BroadcastVoluntaryReleaseTracker_1051_io_alloc_oprb;
  wire  BroadcastAcquireTracker_1052_clk;
  wire  BroadcastAcquireTracker_1052_reset;
  wire  BroadcastAcquireTracker_1052_io_inner_acquire_ready;
  wire  BroadcastAcquireTracker_1052_io_inner_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_1052_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_data;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_id;
  wire  BroadcastAcquireTracker_1052_io_inner_grant_ready;
  wire  BroadcastAcquireTracker_1052_io_inner_grant_valid;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_addr_beat;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_1052_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_data;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_grant_bits_client_id;
  wire  BroadcastAcquireTracker_1052_io_inner_finish_ready;
  wire  BroadcastAcquireTracker_1052_io_inner_finish_valid;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_finish_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_1052_io_inner_probe_ready;
  wire  BroadcastAcquireTracker_1052_io_inner_probe_valid;
  wire [25:0] BroadcastAcquireTracker_1052_io_inner_probe_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_probe_bits_p_type;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_probe_bits_client_id;
  wire  BroadcastAcquireTracker_1052_io_inner_release_ready;
  wire  BroadcastAcquireTracker_1052_io_inner_release_valid;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_release_bits_addr_beat;
  wire [25:0] BroadcastAcquireTracker_1052_io_inner_release_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_release_bits_client_xact_id;
  wire  BroadcastAcquireTracker_1052_io_inner_release_bits_voluntary;
  wire [2:0] BroadcastAcquireTracker_1052_io_inner_release_bits_r_type;
  wire [4:0] BroadcastAcquireTracker_1052_io_inner_release_bits_data;
  wire [1:0] BroadcastAcquireTracker_1052_io_inner_release_bits_client_id;
  wire  BroadcastAcquireTracker_1052_io_incoherent_0;
  wire  BroadcastAcquireTracker_1052_io_outer_acquire_ready;
  wire  BroadcastAcquireTracker_1052_io_outer_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_block;
  wire [2:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_1052_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_1052_io_outer_acquire_bits_data;
  wire  BroadcastAcquireTracker_1052_io_outer_grant_ready;
  wire  BroadcastAcquireTracker_1052_io_outer_grant_valid;
  wire [2:0] BroadcastAcquireTracker_1052_io_outer_grant_bits_addr_beat;
  wire [2:0] BroadcastAcquireTracker_1052_io_outer_grant_bits_client_xact_id;
  wire  BroadcastAcquireTracker_1052_io_outer_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_1052_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_1052_io_outer_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_1052_io_outer_grant_bits_data;
  wire  BroadcastAcquireTracker_1052_io_matches_iacq;
  wire  BroadcastAcquireTracker_1052_io_matches_irel;
  wire  BroadcastAcquireTracker_1052_io_matches_oprb;
  wire  BroadcastAcquireTracker_1052_io_alloc_iacq;
  wire  BroadcastAcquireTracker_1052_io_alloc_irel;
  wire  BroadcastAcquireTracker_1052_io_alloc_oprb;
  wire  BroadcastAcquireTracker_28_1053_clk;
  wire  BroadcastAcquireTracker_28_1053_reset;
  wire  BroadcastAcquireTracker_28_1053_io_inner_acquire_ready;
  wire  BroadcastAcquireTracker_28_1053_io_inner_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_data;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_grant_ready;
  wire  BroadcastAcquireTracker_28_1053_io_inner_grant_valid;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_addr_beat;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_data;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_finish_ready;
  wire  BroadcastAcquireTracker_28_1053_io_inner_finish_valid;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_finish_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_probe_ready;
  wire  BroadcastAcquireTracker_28_1053_io_inner_probe_valid;
  wire [25:0] BroadcastAcquireTracker_28_1053_io_inner_probe_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_probe_bits_p_type;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_probe_bits_client_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_release_ready;
  wire  BroadcastAcquireTracker_28_1053_io_inner_release_valid;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_beat;
  wire [25:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_xact_id;
  wire  BroadcastAcquireTracker_28_1053_io_inner_release_bits_voluntary;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_r_type;
  wire [4:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_data;
  wire [1:0] BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_id;
  wire  BroadcastAcquireTracker_28_1053_io_incoherent_0;
  wire  BroadcastAcquireTracker_28_1053_io_outer_acquire_ready;
  wire  BroadcastAcquireTracker_28_1053_io_outer_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_block;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_data;
  wire  BroadcastAcquireTracker_28_1053_io_outer_grant_ready;
  wire  BroadcastAcquireTracker_28_1053_io_outer_grant_valid;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_outer_grant_bits_addr_beat;
  wire [2:0] BroadcastAcquireTracker_28_1053_io_outer_grant_bits_client_xact_id;
  wire  BroadcastAcquireTracker_28_1053_io_outer_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_28_1053_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_28_1053_io_outer_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_28_1053_io_outer_grant_bits_data;
  wire  BroadcastAcquireTracker_28_1053_io_matches_iacq;
  wire  BroadcastAcquireTracker_28_1053_io_matches_irel;
  wire  BroadcastAcquireTracker_28_1053_io_matches_oprb;
  wire  BroadcastAcquireTracker_28_1053_io_alloc_iacq;
  wire  BroadcastAcquireTracker_28_1053_io_alloc_irel;
  wire  BroadcastAcquireTracker_28_1053_io_alloc_oprb;
  wire  BroadcastAcquireTracker_29_1054_clk;
  wire  BroadcastAcquireTracker_29_1054_reset;
  wire  BroadcastAcquireTracker_29_1054_io_inner_acquire_ready;
  wire  BroadcastAcquireTracker_29_1054_io_inner_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_data;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_grant_ready;
  wire  BroadcastAcquireTracker_29_1054_io_inner_grant_valid;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_addr_beat;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_data;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_finish_ready;
  wire  BroadcastAcquireTracker_29_1054_io_inner_finish_valid;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_finish_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_probe_ready;
  wire  BroadcastAcquireTracker_29_1054_io_inner_probe_valid;
  wire [25:0] BroadcastAcquireTracker_29_1054_io_inner_probe_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_probe_bits_p_type;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_probe_bits_client_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_release_ready;
  wire  BroadcastAcquireTracker_29_1054_io_inner_release_valid;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_beat;
  wire [25:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_xact_id;
  wire  BroadcastAcquireTracker_29_1054_io_inner_release_bits_voluntary;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_r_type;
  wire [4:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_data;
  wire [1:0] BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_id;
  wire  BroadcastAcquireTracker_29_1054_io_incoherent_0;
  wire  BroadcastAcquireTracker_29_1054_io_outer_acquire_ready;
  wire  BroadcastAcquireTracker_29_1054_io_outer_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_block;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_data;
  wire  BroadcastAcquireTracker_29_1054_io_outer_grant_ready;
  wire  BroadcastAcquireTracker_29_1054_io_outer_grant_valid;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_outer_grant_bits_addr_beat;
  wire [2:0] BroadcastAcquireTracker_29_1054_io_outer_grant_bits_client_xact_id;
  wire  BroadcastAcquireTracker_29_1054_io_outer_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_29_1054_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_29_1054_io_outer_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_29_1054_io_outer_grant_bits_data;
  wire  BroadcastAcquireTracker_29_1054_io_matches_iacq;
  wire  BroadcastAcquireTracker_29_1054_io_matches_irel;
  wire  BroadcastAcquireTracker_29_1054_io_matches_oprb;
  wire  BroadcastAcquireTracker_29_1054_io_alloc_iacq;
  wire  BroadcastAcquireTracker_29_1054_io_alloc_irel;
  wire  BroadcastAcquireTracker_29_1054_io_alloc_oprb;
  wire  BroadcastAcquireTracker_30_1055_clk;
  wire  BroadcastAcquireTracker_30_1055_reset;
  wire  BroadcastAcquireTracker_30_1055_io_inner_acquire_ready;
  wire  BroadcastAcquireTracker_30_1055_io_inner_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_data;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_grant_ready;
  wire  BroadcastAcquireTracker_30_1055_io_inner_grant_valid;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_addr_beat;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_data;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_finish_ready;
  wire  BroadcastAcquireTracker_30_1055_io_inner_finish_valid;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_finish_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_probe_ready;
  wire  BroadcastAcquireTracker_30_1055_io_inner_probe_valid;
  wire [25:0] BroadcastAcquireTracker_30_1055_io_inner_probe_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_probe_bits_p_type;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_probe_bits_client_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_release_ready;
  wire  BroadcastAcquireTracker_30_1055_io_inner_release_valid;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_beat;
  wire [25:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_block;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_xact_id;
  wire  BroadcastAcquireTracker_30_1055_io_inner_release_bits_voluntary;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_r_type;
  wire [4:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_data;
  wire [1:0] BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_id;
  wire  BroadcastAcquireTracker_30_1055_io_incoherent_0;
  wire  BroadcastAcquireTracker_30_1055_io_outer_acquire_ready;
  wire  BroadcastAcquireTracker_30_1055_io_outer_acquire_valid;
  wire [25:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_block;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_client_xact_id;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_beat;
  wire  BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_a_type;
  wire [11:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_union;
  wire [4:0] BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_data;
  wire  BroadcastAcquireTracker_30_1055_io_outer_grant_ready;
  wire  BroadcastAcquireTracker_30_1055_io_outer_grant_valid;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_outer_grant_bits_addr_beat;
  wire [2:0] BroadcastAcquireTracker_30_1055_io_outer_grant_bits_client_xact_id;
  wire  BroadcastAcquireTracker_30_1055_io_outer_grant_bits_manager_xact_id;
  wire  BroadcastAcquireTracker_30_1055_io_outer_grant_bits_is_builtin_type;
  wire [3:0] BroadcastAcquireTracker_30_1055_io_outer_grant_bits_g_type;
  wire [4:0] BroadcastAcquireTracker_30_1055_io_outer_grant_bits_data;
  wire  BroadcastAcquireTracker_30_1055_io_matches_iacq;
  wire  BroadcastAcquireTracker_30_1055_io_matches_irel;
  wire  BroadcastAcquireTracker_30_1055_io_matches_oprb;
  wire  BroadcastAcquireTracker_30_1055_io_alloc_iacq;
  wire  BroadcastAcquireTracker_30_1055_io_alloc_irel;
  wire  BroadcastAcquireTracker_30_1055_io_alloc_oprb;
  reg [63:0] sdq_0;
  reg [63:0] GEN_68;
  reg [63:0] sdq_1;
  reg [63:0] GEN_69;
  reg [63:0] sdq_2;
  reg [63:0] GEN_70;
  reg [63:0] sdq_3;
  reg [63:0] GEN_71;
  reg [63:0] sdq_4;
  reg [63:0] GEN_72;
  reg [63:0] sdq_5;
  reg [63:0] GEN_73;
  reg [63:0] sdq_6;
  reg [63:0] GEN_74;
  reg [63:0] sdq_7;
  reg [63:0] GEN_75;
  reg [7:0] sdq_val;
  reg [31:0] GEN_76;
  wire [7:0] T_1063;
  wire  T_1064;
  wire  T_1065;
  wire  T_1066;
  wire  T_1067;
  wire  T_1068;
  wire  T_1069;
  wire  T_1070;
  wire  T_1071;
  wire [2:0] T_1080;
  wire [2:0] T_1081;
  wire [2:0] T_1082;
  wire [2:0] T_1083;
  wire [2:0] T_1084;
  wire [2:0] T_1085;
  wire [2:0] sdq_alloc_id;
  wire [7:0] GEN_59;
  wire  T_1088;
  wire  sdq_rdy;
  wire  T_1090;
  wire  T_1091;
  wire  T_1092;
  wire [2:0] T_1101_0;
  wire [2:0] T_1101_1;
  wire [2:0] T_1101_2;
  wire  T_1103;
  wire  T_1104;
  wire  T_1105;
  wire  T_1108;
  wire  T_1109;
  wire  T_1110;
  wire  T_1111;
  wire  T_1112;
  wire  T_1113;
  wire  T_1114;
  wire [2:0] T_1123_0;
  wire [2:0] T_1123_1;
  wire [2:0] T_1123_2;
  wire  T_1125;
  wire  T_1126;
  wire  T_1127;
  wire  T_1130;
  wire  T_1131;
  wire  T_1132;
  wire  T_1133;
  wire  T_1134;
  wire  T_1135;
  wire  T_1136;
  wire [2:0] T_1145_0;
  wire [2:0] T_1145_1;
  wire [2:0] T_1145_2;
  wire  T_1147;
  wire  T_1148;
  wire  T_1149;
  wire  T_1152;
  wire  T_1153;
  wire  T_1154;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1158;
  wire [2:0] T_1167_0;
  wire [2:0] T_1167_1;
  wire [2:0] T_1167_2;
  wire  T_1169;
  wire  T_1170;
  wire  T_1171;
  wire  T_1174;
  wire  T_1175;
  wire  T_1176;
  wire  T_1177;
  wire  T_1178;
  wire  T_1179;
  wire  T_1180;
  wire [2:0] T_1189_0;
  wire [2:0] T_1189_1;
  wire [2:0] T_1189_2;
  wire  T_1191;
  wire  T_1192;
  wire  T_1193;
  wire  T_1196;
  wire  T_1197;
  wire  T_1198;
  wire  T_1199;
  wire  T_1200;
  wire  T_1201;
  wire  T_1202;
  wire  sdq_enq;
  wire [63:0] GEN_0;
  wire [2:0] GEN_60;
  wire [63:0] GEN_5;
  wire [2:0] GEN_61;
  wire [63:0] GEN_6;
  wire [2:0] GEN_62;
  wire [63:0] GEN_7;
  wire [2:0] GEN_63;
  wire [63:0] GEN_8;
  wire [63:0] GEN_9;
  wire [63:0] GEN_10;
  wire [63:0] GEN_11;
  wire [63:0] GEN_12;
  wire [63:0] GEN_14;
  wire [63:0] GEN_15;
  wire [63:0] GEN_16;
  wire [63:0] GEN_17;
  wire [63:0] GEN_18;
  wire [63:0] GEN_19;
  wire [63:0] GEN_20;
  wire [63:0] GEN_21;
  wire  T_1203;
  wire  T_1204;
  wire  irel_vs_iacq_conflict;
  wire [2:0] T_1251_idx;
  wire [1:0] T_1251_loc;
  wire [4:0] T_1297;
  wire [2:0] T_1344_idx;
  wire [1:0] T_1344_loc;
  wire [4:0] T_1390;
  wire [2:0] T_1437_idx;
  wire [1:0] T_1437_loc;
  wire [4:0] T_1483;
  wire [2:0] T_1530_idx;
  wire [1:0] T_1530_loc;
  wire [4:0] T_1576;
  wire [2:0] T_1623_idx;
  wire [1:0] T_1623_loc;
  wire [4:0] T_1669;
  wire  T_1671;
  wire  T_1672;
  wire  T_1678_0;
  wire  T_1678_1;
  wire  T_1678_2;
  wire  T_1678_3;
  wire  T_1678_4;
  wire [1:0] T_1680;
  wire [1:0] T_1681;
  wire [2:0] T_1682;
  wire [4:0] T_1683;
  wire  T_1684;
  wire  T_1685;
  wire  T_1686;
  wire  T_1687;
  wire  T_1688;
  wire [4:0] T_1696;
  wire [4:0] T_1697;
  wire [4:0] T_1698;
  wire [4:0] T_1699;
  wire [4:0] T_1700;
  wire  T_1706_0;
  wire  T_1706_1;
  wire  T_1706_2;
  wire  T_1706_3;
  wire  T_1706_4;
  wire [1:0] T_1708;
  wire [1:0] T_1709;
  wire [2:0] T_1710;
  wire [4:0] T_1711;
  wire [4:0] GEN_64;
  wire  T_1713;
  wire  T_1715;
  wire  T_1717;
  wire [4:0] T_1718;
  wire  T_1720;
  wire  T_1721;
  wire  T_1722;
  wire  T_1723;
  wire  T_1724;
  wire  T_1725;
  wire  T_1726;
  wire  T_1727;
  wire  T_1728;
  wire  T_1731;
  wire  T_1732;
  wire  T_1733;
  wire  T_1736;
  wire  T_1737;
  wire  T_1738;
  wire  T_1741;
  wire  T_1742;
  wire  T_1743;
  wire  T_1746;
  wire  T_1747;
  wire  T_1748;
  wire  T_1749;
  wire  T_1750;
  wire [2:0] T_1756_0;
  wire [2:0] T_1756_1;
  wire [2:0] T_1756_2;
  wire  T_1758;
  wire  T_1759;
  wire  T_1760;
  wire  T_1763;
  wire  T_1764;
  wire  vwbdq_enq;
  reg [2:0] rel_data_cnt;
  reg [31:0] GEN_77;
  wire [3:0] T_1769;
  wire [2:0] T_1770;
  wire [2:0] GEN_22;
  reg [63:0] vwbdq_0;
  reg [63:0] GEN_78;
  reg [63:0] vwbdq_1;
  reg [63:0] GEN_79;
  reg [63:0] vwbdq_2;
  reg [63:0] GEN_80;
  reg [63:0] vwbdq_3;
  reg [63:0] GEN_81;
  reg [63:0] vwbdq_4;
  reg [63:0] GEN_82;
  reg [63:0] vwbdq_5;
  reg [63:0] GEN_83;
  reg [63:0] vwbdq_6;
  reg [63:0] GEN_84;
  reg [63:0] vwbdq_7;
  reg [63:0] GEN_85;
  wire [63:0] GEN_1;
  wire [63:0] GEN_23;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [63:0] GEN_26;
  wire [63:0] GEN_27;
  wire [63:0] GEN_28;
  wire [63:0] GEN_29;
  wire [63:0] GEN_30;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [2:0] T_1823_idx;
  wire [1:0] T_1823_loc;
  wire [4:0] T_1869;
  wire [2:0] T_1916_idx;
  wire [1:0] T_1916_loc;
  wire [4:0] T_1962;
  wire [2:0] T_2009_idx;
  wire [1:0] T_2009_loc;
  wire [4:0] T_2055;
  wire [2:0] T_2102_idx;
  wire [1:0] T_2102_loc;
  wire [4:0] T_2148;
  wire [2:0] T_2195_idx;
  wire [1:0] T_2195_loc;
  wire [4:0] T_2241;
  wire  T_2247_0;
  wire  T_2247_1;
  wire  T_2247_2;
  wire  T_2247_3;
  wire  T_2247_4;
  wire [1:0] T_2249;
  wire [1:0] T_2250;
  wire [2:0] T_2251;
  wire [4:0] T_2252;
  wire  T_2253;
  wire  T_2254;
  wire  T_2255;
  wire  T_2256;
  wire  T_2257;
  wire [4:0] T_2265;
  wire [4:0] T_2266;
  wire [4:0] T_2267;
  wire [4:0] T_2268;
  wire [4:0] T_2269;
  wire  T_2275_0;
  wire  T_2275_1;
  wire  T_2275_2;
  wire  T_2275_3;
  wire  T_2275_4;
  wire [1:0] T_2277;
  wire [1:0] T_2278;
  wire [2:0] T_2279;
  wire [4:0] T_2280;
  wire  T_2282;
  wire  T_2284;
  wire  T_2288;
  wire [4:0] T_2289;
  wire  T_2291;
  wire  T_2292;
  wire  T_2297;
  wire  T_2298;
  wire  T_2302;
  wire  T_2303;
  wire  T_2307;
  wire  T_2308;
  wire  T_2312;
  wire  T_2313;
  wire  T_2317;
  wire  T_2318;
  wire  LockingRRArbiter_31_2320_clk;
  wire  LockingRRArbiter_31_2320_reset;
  wire  LockingRRArbiter_31_2320_io_in_0_ready;
  wire  LockingRRArbiter_31_2320_io_in_0_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_in_0_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_in_0_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_in_0_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_in_0_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_in_0_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_in_0_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_in_0_bits_client_id;
  wire  LockingRRArbiter_31_2320_io_in_1_ready;
  wire  LockingRRArbiter_31_2320_io_in_1_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_in_1_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_in_1_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_in_1_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_in_1_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_in_1_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_in_1_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_in_1_bits_client_id;
  wire  LockingRRArbiter_31_2320_io_in_2_ready;
  wire  LockingRRArbiter_31_2320_io_in_2_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_in_2_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_in_2_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_in_2_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_in_2_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_in_2_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_in_2_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_in_2_bits_client_id;
  wire  LockingRRArbiter_31_2320_io_in_3_ready;
  wire  LockingRRArbiter_31_2320_io_in_3_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_in_3_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_in_3_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_in_3_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_in_3_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_in_3_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_in_3_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_in_3_bits_client_id;
  wire  LockingRRArbiter_31_2320_io_in_4_ready;
  wire  LockingRRArbiter_31_2320_io_in_4_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_in_4_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_in_4_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_in_4_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_in_4_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_in_4_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_in_4_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_in_4_bits_client_id;
  wire  LockingRRArbiter_31_2320_io_out_ready;
  wire  LockingRRArbiter_31_2320_io_out_valid;
  wire [2:0] LockingRRArbiter_31_2320_io_out_bits_addr_beat;
  wire [1:0] LockingRRArbiter_31_2320_io_out_bits_client_xact_id;
  wire [2:0] LockingRRArbiter_31_2320_io_out_bits_manager_xact_id;
  wire  LockingRRArbiter_31_2320_io_out_bits_is_builtin_type;
  wire [3:0] LockingRRArbiter_31_2320_io_out_bits_g_type;
  wire [63:0] LockingRRArbiter_31_2320_io_out_bits_data;
  wire [1:0] LockingRRArbiter_31_2320_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_31_2320_io_chosen;
  wire  LockingRRArbiter_32_2321_clk;
  wire  LockingRRArbiter_32_2321_reset;
  wire  LockingRRArbiter_32_2321_io_in_0_ready;
  wire  LockingRRArbiter_32_2321_io_in_0_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_in_0_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_in_0_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_in_0_bits_client_id;
  wire  LockingRRArbiter_32_2321_io_in_1_ready;
  wire  LockingRRArbiter_32_2321_io_in_1_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_in_1_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_in_1_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_in_1_bits_client_id;
  wire  LockingRRArbiter_32_2321_io_in_2_ready;
  wire  LockingRRArbiter_32_2321_io_in_2_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_in_2_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_in_2_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_in_2_bits_client_id;
  wire  LockingRRArbiter_32_2321_io_in_3_ready;
  wire  LockingRRArbiter_32_2321_io_in_3_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_in_3_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_in_3_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_in_3_bits_client_id;
  wire  LockingRRArbiter_32_2321_io_in_4_ready;
  wire  LockingRRArbiter_32_2321_io_in_4_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_in_4_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_in_4_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_in_4_bits_client_id;
  wire  LockingRRArbiter_32_2321_io_out_ready;
  wire  LockingRRArbiter_32_2321_io_out_valid;
  wire [25:0] LockingRRArbiter_32_2321_io_out_bits_addr_block;
  wire [1:0] LockingRRArbiter_32_2321_io_out_bits_p_type;
  wire [1:0] LockingRRArbiter_32_2321_io_out_bits_client_id;
  wire [2:0] LockingRRArbiter_32_2321_io_chosen;
  wire  T_2323;
  wire  T_2324;
  wire  T_2326;
  wire  T_2327;
  wire  T_2329;
  wire  T_2330;
  wire  T_2332;
  wire  T_2333;
  wire  T_2335;
  wire  T_2336;
  wire  T_2342_0;
  wire  T_2342_1;
  wire  T_2342_2;
  wire  T_2342_3;
  wire  T_2342_4;
  wire  GEN_2;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  outer_arb_clk;
  wire  outer_arb_reset;
  wire  outer_arb_io_in_0_acquire_ready;
  wire  outer_arb_io_in_0_acquire_valid;
  wire [25:0] outer_arb_io_in_0_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_0_acquire_bits_addr_beat;
  wire  outer_arb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_0_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_0_acquire_bits_union;
  wire [4:0] outer_arb_io_in_0_acquire_bits_data;
  wire  outer_arb_io_in_0_grant_ready;
  wire  outer_arb_io_in_0_grant_valid;
  wire [2:0] outer_arb_io_in_0_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_0_grant_bits_client_xact_id;
  wire  outer_arb_io_in_0_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_0_grant_bits_g_type;
  wire [4:0] outer_arb_io_in_0_grant_bits_data;
  wire  outer_arb_io_in_1_acquire_ready;
  wire  outer_arb_io_in_1_acquire_valid;
  wire [25:0] outer_arb_io_in_1_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_1_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_1_acquire_bits_addr_beat;
  wire  outer_arb_io_in_1_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_1_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_1_acquire_bits_union;
  wire [4:0] outer_arb_io_in_1_acquire_bits_data;
  wire  outer_arb_io_in_1_grant_ready;
  wire  outer_arb_io_in_1_grant_valid;
  wire [2:0] outer_arb_io_in_1_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_1_grant_bits_client_xact_id;
  wire  outer_arb_io_in_1_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_1_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_1_grant_bits_g_type;
  wire [4:0] outer_arb_io_in_1_grant_bits_data;
  wire  outer_arb_io_in_2_acquire_ready;
  wire  outer_arb_io_in_2_acquire_valid;
  wire [25:0] outer_arb_io_in_2_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_2_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_2_acquire_bits_addr_beat;
  wire  outer_arb_io_in_2_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_2_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_2_acquire_bits_union;
  wire [4:0] outer_arb_io_in_2_acquire_bits_data;
  wire  outer_arb_io_in_2_grant_ready;
  wire  outer_arb_io_in_2_grant_valid;
  wire [2:0] outer_arb_io_in_2_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_2_grant_bits_client_xact_id;
  wire  outer_arb_io_in_2_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_2_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_2_grant_bits_g_type;
  wire [4:0] outer_arb_io_in_2_grant_bits_data;
  wire  outer_arb_io_in_3_acquire_ready;
  wire  outer_arb_io_in_3_acquire_valid;
  wire [25:0] outer_arb_io_in_3_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_3_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_3_acquire_bits_addr_beat;
  wire  outer_arb_io_in_3_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_3_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_3_acquire_bits_union;
  wire [4:0] outer_arb_io_in_3_acquire_bits_data;
  wire  outer_arb_io_in_3_grant_ready;
  wire  outer_arb_io_in_3_grant_valid;
  wire [2:0] outer_arb_io_in_3_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_3_grant_bits_client_xact_id;
  wire  outer_arb_io_in_3_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_3_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_3_grant_bits_g_type;
  wire [4:0] outer_arb_io_in_3_grant_bits_data;
  wire  outer_arb_io_in_4_acquire_ready;
  wire  outer_arb_io_in_4_acquire_valid;
  wire [25:0] outer_arb_io_in_4_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_in_4_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_in_4_acquire_bits_addr_beat;
  wire  outer_arb_io_in_4_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_in_4_acquire_bits_a_type;
  wire [11:0] outer_arb_io_in_4_acquire_bits_union;
  wire [4:0] outer_arb_io_in_4_acquire_bits_data;
  wire  outer_arb_io_in_4_grant_ready;
  wire  outer_arb_io_in_4_grant_valid;
  wire [2:0] outer_arb_io_in_4_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_in_4_grant_bits_client_xact_id;
  wire  outer_arb_io_in_4_grant_bits_manager_xact_id;
  wire  outer_arb_io_in_4_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_in_4_grant_bits_g_type;
  wire [4:0] outer_arb_io_in_4_grant_bits_data;
  wire  outer_arb_io_out_acquire_ready;
  wire  outer_arb_io_out_acquire_valid;
  wire [25:0] outer_arb_io_out_acquire_bits_addr_block;
  wire [2:0] outer_arb_io_out_acquire_bits_client_xact_id;
  wire [2:0] outer_arb_io_out_acquire_bits_addr_beat;
  wire  outer_arb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] outer_arb_io_out_acquire_bits_a_type;
  wire [11:0] outer_arb_io_out_acquire_bits_union;
  wire [4:0] outer_arb_io_out_acquire_bits_data;
  wire  outer_arb_io_out_grant_ready;
  wire  outer_arb_io_out_grant_valid;
  wire [2:0] outer_arb_io_out_grant_bits_addr_beat;
  wire [2:0] outer_arb_io_out_grant_bits_client_xact_id;
  wire  outer_arb_io_out_grant_bits_manager_xact_id;
  wire  outer_arb_io_out_grant_bits_is_builtin_type;
  wire [3:0] outer_arb_io_out_grant_bits_g_type;
  wire [4:0] outer_arb_io_out_grant_bits_data;
  wire [2:0] outer_data_ptr_idx;
  wire [1:0] outer_data_ptr_loc;
  wire [1:0] T_2481;
  wire [2:0] T_2482;
  wire  is_in_sdq;
  wire  T_2483;
  wire [2:0] T_2492_0;
  wire [2:0] T_2492_1;
  wire [2:0] T_2492_2;
  wire  T_2494;
  wire  T_2495;
  wire  T_2496;
  wire  T_2499;
  wire  T_2500;
  wire  T_2501;
  wire  T_2502;
  wire  free_sdq;
  wire  T_2504;
  wire [63:0] GEN_3;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] T_2505;
  wire  T_2506;
  wire [63:0] GEN_4;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire [63:0] GEN_55;
  wire [63:0] GEN_56;
  wire [63:0] GEN_57;
  wire [63:0] T_2507;
  wire  T_2508;
  wire [7:0] GEN_88;
  wire [7:0] T_2510;
  wire [7:0] GEN_89;
  wire [8:0] T_2512;
  wire [7:0] T_2513;
  wire [7:0] T_2514;
  wire [7:0] T_2515;
  wire [7:0] T_2516;
  wire [7:0] T_2537;
  wire [7:0] T_2538;
  wire [7:0] T_2539;
  wire [7:0] T_2540;
  wire [7:0] T_2541;
  wire [7:0] T_2542;
  wire [7:0] T_2543;
  wire [7:0] T_2544;
  wire [7:0] GEN_90;
  wire [8:0] T_2546;
  wire [7:0] T_2547;
  wire [7:0] T_2548;
  wire [7:0] T_2549;
  wire [7:0] GEN_58;
  reg  GEN_13;
  reg [31:0] GEN_86;
  reg  GEN_31;
  reg [31:0] GEN_87;
  reg  GEN_65;
  reg [31:0] GEN_91;
  reg  GEN_66;
  reg [31:0] GEN_92;
  reg  GEN_67;
  reg [31:0] GEN_93;
  BroadcastVoluntaryReleaseTracker BroadcastVoluntaryReleaseTracker_1051 (
    .clk(BroadcastVoluntaryReleaseTracker_1051_clk),
    .reset(BroadcastVoluntaryReleaseTracker_1051_reset),
    .io_inner_acquire_ready(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_ready),
    .io_inner_acquire_valid(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_ready),
    .io_inner_grant_valid(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_ready),
    .io_inner_finish_valid(BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_ready),
    .io_inner_probe_valid(BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_ready),
    .io_inner_release_valid(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_id),
    .io_incoherent_0(BroadcastVoluntaryReleaseTracker_1051_io_incoherent_0),
    .io_outer_acquire_ready(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_ready),
    .io_outer_acquire_valid(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_data),
    .io_outer_grant_ready(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_ready),
    .io_outer_grant_valid(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_data),
    .io_matches_iacq(BroadcastVoluntaryReleaseTracker_1051_io_matches_iacq),
    .io_matches_irel(BroadcastVoluntaryReleaseTracker_1051_io_matches_irel),
    .io_matches_oprb(BroadcastVoluntaryReleaseTracker_1051_io_matches_oprb),
    .io_alloc_iacq(BroadcastVoluntaryReleaseTracker_1051_io_alloc_iacq),
    .io_alloc_irel(BroadcastVoluntaryReleaseTracker_1051_io_alloc_irel),
    .io_alloc_oprb(BroadcastVoluntaryReleaseTracker_1051_io_alloc_oprb)
  );
  BroadcastAcquireTracker BroadcastAcquireTracker_1052 (
    .clk(BroadcastAcquireTracker_1052_clk),
    .reset(BroadcastAcquireTracker_1052_reset),
    .io_inner_acquire_ready(BroadcastAcquireTracker_1052_io_inner_acquire_ready),
    .io_inner_acquire_valid(BroadcastAcquireTracker_1052_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BroadcastAcquireTracker_1052_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BroadcastAcquireTracker_1052_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BroadcastAcquireTracker_1052_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BroadcastAcquireTracker_1052_io_inner_grant_ready),
    .io_inner_grant_valid(BroadcastAcquireTracker_1052_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BroadcastAcquireTracker_1052_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BroadcastAcquireTracker_1052_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BroadcastAcquireTracker_1052_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BroadcastAcquireTracker_1052_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BroadcastAcquireTracker_1052_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BroadcastAcquireTracker_1052_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BroadcastAcquireTracker_1052_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BroadcastAcquireTracker_1052_io_inner_finish_ready),
    .io_inner_finish_valid(BroadcastAcquireTracker_1052_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BroadcastAcquireTracker_1052_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BroadcastAcquireTracker_1052_io_inner_probe_ready),
    .io_inner_probe_valid(BroadcastAcquireTracker_1052_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BroadcastAcquireTracker_1052_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BroadcastAcquireTracker_1052_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BroadcastAcquireTracker_1052_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BroadcastAcquireTracker_1052_io_inner_release_ready),
    .io_inner_release_valid(BroadcastAcquireTracker_1052_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BroadcastAcquireTracker_1052_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BroadcastAcquireTracker_1052_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BroadcastAcquireTracker_1052_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BroadcastAcquireTracker_1052_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BroadcastAcquireTracker_1052_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BroadcastAcquireTracker_1052_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BroadcastAcquireTracker_1052_io_inner_release_bits_client_id),
    .io_incoherent_0(BroadcastAcquireTracker_1052_io_incoherent_0),
    .io_outer_acquire_ready(BroadcastAcquireTracker_1052_io_outer_acquire_ready),
    .io_outer_acquire_valid(BroadcastAcquireTracker_1052_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BroadcastAcquireTracker_1052_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BroadcastAcquireTracker_1052_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BroadcastAcquireTracker_1052_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BroadcastAcquireTracker_1052_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BroadcastAcquireTracker_1052_io_outer_acquire_bits_data),
    .io_outer_grant_ready(BroadcastAcquireTracker_1052_io_outer_grant_ready),
    .io_outer_grant_valid(BroadcastAcquireTracker_1052_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BroadcastAcquireTracker_1052_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BroadcastAcquireTracker_1052_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BroadcastAcquireTracker_1052_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BroadcastAcquireTracker_1052_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BroadcastAcquireTracker_1052_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BroadcastAcquireTracker_1052_io_outer_grant_bits_data),
    .io_matches_iacq(BroadcastAcquireTracker_1052_io_matches_iacq),
    .io_matches_irel(BroadcastAcquireTracker_1052_io_matches_irel),
    .io_matches_oprb(BroadcastAcquireTracker_1052_io_matches_oprb),
    .io_alloc_iacq(BroadcastAcquireTracker_1052_io_alloc_iacq),
    .io_alloc_irel(BroadcastAcquireTracker_1052_io_alloc_irel),
    .io_alloc_oprb(BroadcastAcquireTracker_1052_io_alloc_oprb)
  );
  BroadcastAcquireTracker_28 BroadcastAcquireTracker_28_1053 (
    .clk(BroadcastAcquireTracker_28_1053_clk),
    .reset(BroadcastAcquireTracker_28_1053_reset),
    .io_inner_acquire_ready(BroadcastAcquireTracker_28_1053_io_inner_acquire_ready),
    .io_inner_acquire_valid(BroadcastAcquireTracker_28_1053_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BroadcastAcquireTracker_28_1053_io_inner_grant_ready),
    .io_inner_grant_valid(BroadcastAcquireTracker_28_1053_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BroadcastAcquireTracker_28_1053_io_inner_finish_ready),
    .io_inner_finish_valid(BroadcastAcquireTracker_28_1053_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BroadcastAcquireTracker_28_1053_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BroadcastAcquireTracker_28_1053_io_inner_probe_ready),
    .io_inner_probe_valid(BroadcastAcquireTracker_28_1053_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BroadcastAcquireTracker_28_1053_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BroadcastAcquireTracker_28_1053_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BroadcastAcquireTracker_28_1053_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BroadcastAcquireTracker_28_1053_io_inner_release_ready),
    .io_inner_release_valid(BroadcastAcquireTracker_28_1053_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BroadcastAcquireTracker_28_1053_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BroadcastAcquireTracker_28_1053_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BroadcastAcquireTracker_28_1053_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_id),
    .io_incoherent_0(BroadcastAcquireTracker_28_1053_io_incoherent_0),
    .io_outer_acquire_ready(BroadcastAcquireTracker_28_1053_io_outer_acquire_ready),
    .io_outer_acquire_valid(BroadcastAcquireTracker_28_1053_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_data),
    .io_outer_grant_ready(BroadcastAcquireTracker_28_1053_io_outer_grant_ready),
    .io_outer_grant_valid(BroadcastAcquireTracker_28_1053_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BroadcastAcquireTracker_28_1053_io_outer_grant_bits_data),
    .io_matches_iacq(BroadcastAcquireTracker_28_1053_io_matches_iacq),
    .io_matches_irel(BroadcastAcquireTracker_28_1053_io_matches_irel),
    .io_matches_oprb(BroadcastAcquireTracker_28_1053_io_matches_oprb),
    .io_alloc_iacq(BroadcastAcquireTracker_28_1053_io_alloc_iacq),
    .io_alloc_irel(BroadcastAcquireTracker_28_1053_io_alloc_irel),
    .io_alloc_oprb(BroadcastAcquireTracker_28_1053_io_alloc_oprb)
  );
  BroadcastAcquireTracker_29 BroadcastAcquireTracker_29_1054 (
    .clk(BroadcastAcquireTracker_29_1054_clk),
    .reset(BroadcastAcquireTracker_29_1054_reset),
    .io_inner_acquire_ready(BroadcastAcquireTracker_29_1054_io_inner_acquire_ready),
    .io_inner_acquire_valid(BroadcastAcquireTracker_29_1054_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BroadcastAcquireTracker_29_1054_io_inner_grant_ready),
    .io_inner_grant_valid(BroadcastAcquireTracker_29_1054_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BroadcastAcquireTracker_29_1054_io_inner_finish_ready),
    .io_inner_finish_valid(BroadcastAcquireTracker_29_1054_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BroadcastAcquireTracker_29_1054_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BroadcastAcquireTracker_29_1054_io_inner_probe_ready),
    .io_inner_probe_valid(BroadcastAcquireTracker_29_1054_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BroadcastAcquireTracker_29_1054_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BroadcastAcquireTracker_29_1054_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BroadcastAcquireTracker_29_1054_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BroadcastAcquireTracker_29_1054_io_inner_release_ready),
    .io_inner_release_valid(BroadcastAcquireTracker_29_1054_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BroadcastAcquireTracker_29_1054_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BroadcastAcquireTracker_29_1054_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BroadcastAcquireTracker_29_1054_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_id),
    .io_incoherent_0(BroadcastAcquireTracker_29_1054_io_incoherent_0),
    .io_outer_acquire_ready(BroadcastAcquireTracker_29_1054_io_outer_acquire_ready),
    .io_outer_acquire_valid(BroadcastAcquireTracker_29_1054_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_data),
    .io_outer_grant_ready(BroadcastAcquireTracker_29_1054_io_outer_grant_ready),
    .io_outer_grant_valid(BroadcastAcquireTracker_29_1054_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BroadcastAcquireTracker_29_1054_io_outer_grant_bits_data),
    .io_matches_iacq(BroadcastAcquireTracker_29_1054_io_matches_iacq),
    .io_matches_irel(BroadcastAcquireTracker_29_1054_io_matches_irel),
    .io_matches_oprb(BroadcastAcquireTracker_29_1054_io_matches_oprb),
    .io_alloc_iacq(BroadcastAcquireTracker_29_1054_io_alloc_iacq),
    .io_alloc_irel(BroadcastAcquireTracker_29_1054_io_alloc_irel),
    .io_alloc_oprb(BroadcastAcquireTracker_29_1054_io_alloc_oprb)
  );
  BroadcastAcquireTracker_30 BroadcastAcquireTracker_30_1055 (
    .clk(BroadcastAcquireTracker_30_1055_clk),
    .reset(BroadcastAcquireTracker_30_1055_reset),
    .io_inner_acquire_ready(BroadcastAcquireTracker_30_1055_io_inner_acquire_ready),
    .io_inner_acquire_valid(BroadcastAcquireTracker_30_1055_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(BroadcastAcquireTracker_30_1055_io_inner_grant_ready),
    .io_inner_grant_valid(BroadcastAcquireTracker_30_1055_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(BroadcastAcquireTracker_30_1055_io_inner_finish_ready),
    .io_inner_finish_valid(BroadcastAcquireTracker_30_1055_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(BroadcastAcquireTracker_30_1055_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(BroadcastAcquireTracker_30_1055_io_inner_probe_ready),
    .io_inner_probe_valid(BroadcastAcquireTracker_30_1055_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(BroadcastAcquireTracker_30_1055_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(BroadcastAcquireTracker_30_1055_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(BroadcastAcquireTracker_30_1055_io_inner_probe_bits_client_id),
    .io_inner_release_ready(BroadcastAcquireTracker_30_1055_io_inner_release_ready),
    .io_inner_release_valid(BroadcastAcquireTracker_30_1055_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(BroadcastAcquireTracker_30_1055_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(BroadcastAcquireTracker_30_1055_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(BroadcastAcquireTracker_30_1055_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_id),
    .io_incoherent_0(BroadcastAcquireTracker_30_1055_io_incoherent_0),
    .io_outer_acquire_ready(BroadcastAcquireTracker_30_1055_io_outer_acquire_ready),
    .io_outer_acquire_valid(BroadcastAcquireTracker_30_1055_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_data),
    .io_outer_grant_ready(BroadcastAcquireTracker_30_1055_io_outer_grant_ready),
    .io_outer_grant_valid(BroadcastAcquireTracker_30_1055_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(BroadcastAcquireTracker_30_1055_io_outer_grant_bits_data),
    .io_matches_iacq(BroadcastAcquireTracker_30_1055_io_matches_iacq),
    .io_matches_irel(BroadcastAcquireTracker_30_1055_io_matches_irel),
    .io_matches_oprb(BroadcastAcquireTracker_30_1055_io_matches_oprb),
    .io_alloc_iacq(BroadcastAcquireTracker_30_1055_io_alloc_iacq),
    .io_alloc_irel(BroadcastAcquireTracker_30_1055_io_alloc_irel),
    .io_alloc_oprb(BroadcastAcquireTracker_30_1055_io_alloc_oprb)
  );
  LockingRRArbiter_31 LockingRRArbiter_31_2320 (
    .clk(LockingRRArbiter_31_2320_clk),
    .reset(LockingRRArbiter_31_2320_reset),
    .io_in_0_ready(LockingRRArbiter_31_2320_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_31_2320_io_in_0_valid),
    .io_in_0_bits_addr_beat(LockingRRArbiter_31_2320_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(LockingRRArbiter_31_2320_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(LockingRRArbiter_31_2320_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(LockingRRArbiter_31_2320_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(LockingRRArbiter_31_2320_io_in_0_bits_g_type),
    .io_in_0_bits_data(LockingRRArbiter_31_2320_io_in_0_bits_data),
    .io_in_0_bits_client_id(LockingRRArbiter_31_2320_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_31_2320_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_31_2320_io_in_1_valid),
    .io_in_1_bits_addr_beat(LockingRRArbiter_31_2320_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(LockingRRArbiter_31_2320_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(LockingRRArbiter_31_2320_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(LockingRRArbiter_31_2320_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(LockingRRArbiter_31_2320_io_in_1_bits_g_type),
    .io_in_1_bits_data(LockingRRArbiter_31_2320_io_in_1_bits_data),
    .io_in_1_bits_client_id(LockingRRArbiter_31_2320_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_31_2320_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_31_2320_io_in_2_valid),
    .io_in_2_bits_addr_beat(LockingRRArbiter_31_2320_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(LockingRRArbiter_31_2320_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(LockingRRArbiter_31_2320_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(LockingRRArbiter_31_2320_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(LockingRRArbiter_31_2320_io_in_2_bits_g_type),
    .io_in_2_bits_data(LockingRRArbiter_31_2320_io_in_2_bits_data),
    .io_in_2_bits_client_id(LockingRRArbiter_31_2320_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_31_2320_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_31_2320_io_in_3_valid),
    .io_in_3_bits_addr_beat(LockingRRArbiter_31_2320_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(LockingRRArbiter_31_2320_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(LockingRRArbiter_31_2320_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(LockingRRArbiter_31_2320_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(LockingRRArbiter_31_2320_io_in_3_bits_g_type),
    .io_in_3_bits_data(LockingRRArbiter_31_2320_io_in_3_bits_data),
    .io_in_3_bits_client_id(LockingRRArbiter_31_2320_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_31_2320_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_31_2320_io_in_4_valid),
    .io_in_4_bits_addr_beat(LockingRRArbiter_31_2320_io_in_4_bits_addr_beat),
    .io_in_4_bits_client_xact_id(LockingRRArbiter_31_2320_io_in_4_bits_client_xact_id),
    .io_in_4_bits_manager_xact_id(LockingRRArbiter_31_2320_io_in_4_bits_manager_xact_id),
    .io_in_4_bits_is_builtin_type(LockingRRArbiter_31_2320_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_g_type(LockingRRArbiter_31_2320_io_in_4_bits_g_type),
    .io_in_4_bits_data(LockingRRArbiter_31_2320_io_in_4_bits_data),
    .io_in_4_bits_client_id(LockingRRArbiter_31_2320_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_31_2320_io_out_ready),
    .io_out_valid(LockingRRArbiter_31_2320_io_out_valid),
    .io_out_bits_addr_beat(LockingRRArbiter_31_2320_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(LockingRRArbiter_31_2320_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(LockingRRArbiter_31_2320_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(LockingRRArbiter_31_2320_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(LockingRRArbiter_31_2320_io_out_bits_g_type),
    .io_out_bits_data(LockingRRArbiter_31_2320_io_out_bits_data),
    .io_out_bits_client_id(LockingRRArbiter_31_2320_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_31_2320_io_chosen)
  );
  LockingRRArbiter_32 LockingRRArbiter_32_2321 (
    .clk(LockingRRArbiter_32_2321_clk),
    .reset(LockingRRArbiter_32_2321_reset),
    .io_in_0_ready(LockingRRArbiter_32_2321_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_32_2321_io_in_0_valid),
    .io_in_0_bits_addr_block(LockingRRArbiter_32_2321_io_in_0_bits_addr_block),
    .io_in_0_bits_p_type(LockingRRArbiter_32_2321_io_in_0_bits_p_type),
    .io_in_0_bits_client_id(LockingRRArbiter_32_2321_io_in_0_bits_client_id),
    .io_in_1_ready(LockingRRArbiter_32_2321_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_32_2321_io_in_1_valid),
    .io_in_1_bits_addr_block(LockingRRArbiter_32_2321_io_in_1_bits_addr_block),
    .io_in_1_bits_p_type(LockingRRArbiter_32_2321_io_in_1_bits_p_type),
    .io_in_1_bits_client_id(LockingRRArbiter_32_2321_io_in_1_bits_client_id),
    .io_in_2_ready(LockingRRArbiter_32_2321_io_in_2_ready),
    .io_in_2_valid(LockingRRArbiter_32_2321_io_in_2_valid),
    .io_in_2_bits_addr_block(LockingRRArbiter_32_2321_io_in_2_bits_addr_block),
    .io_in_2_bits_p_type(LockingRRArbiter_32_2321_io_in_2_bits_p_type),
    .io_in_2_bits_client_id(LockingRRArbiter_32_2321_io_in_2_bits_client_id),
    .io_in_3_ready(LockingRRArbiter_32_2321_io_in_3_ready),
    .io_in_3_valid(LockingRRArbiter_32_2321_io_in_3_valid),
    .io_in_3_bits_addr_block(LockingRRArbiter_32_2321_io_in_3_bits_addr_block),
    .io_in_3_bits_p_type(LockingRRArbiter_32_2321_io_in_3_bits_p_type),
    .io_in_3_bits_client_id(LockingRRArbiter_32_2321_io_in_3_bits_client_id),
    .io_in_4_ready(LockingRRArbiter_32_2321_io_in_4_ready),
    .io_in_4_valid(LockingRRArbiter_32_2321_io_in_4_valid),
    .io_in_4_bits_addr_block(LockingRRArbiter_32_2321_io_in_4_bits_addr_block),
    .io_in_4_bits_p_type(LockingRRArbiter_32_2321_io_in_4_bits_p_type),
    .io_in_4_bits_client_id(LockingRRArbiter_32_2321_io_in_4_bits_client_id),
    .io_out_ready(LockingRRArbiter_32_2321_io_out_ready),
    .io_out_valid(LockingRRArbiter_32_2321_io_out_valid),
    .io_out_bits_addr_block(LockingRRArbiter_32_2321_io_out_bits_addr_block),
    .io_out_bits_p_type(LockingRRArbiter_32_2321_io_out_bits_p_type),
    .io_out_bits_client_id(LockingRRArbiter_32_2321_io_out_bits_client_id),
    .io_chosen(LockingRRArbiter_32_2321_io_chosen)
  );
  ClientUncachedTileLinkIOArbiter outer_arb (
    .clk(outer_arb_clk),
    .reset(outer_arb_reset),
    .io_in_0_acquire_ready(outer_arb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(outer_arb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(outer_arb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(outer_arb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(outer_arb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(outer_arb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(outer_arb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(outer_arb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(outer_arb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(outer_arb_io_in_0_grant_ready),
    .io_in_0_grant_valid(outer_arb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(outer_arb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(outer_arb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(outer_arb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(outer_arb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(outer_arb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(outer_arb_io_in_0_grant_bits_data),
    .io_in_1_acquire_ready(outer_arb_io_in_1_acquire_ready),
    .io_in_1_acquire_valid(outer_arb_io_in_1_acquire_valid),
    .io_in_1_acquire_bits_addr_block(outer_arb_io_in_1_acquire_bits_addr_block),
    .io_in_1_acquire_bits_client_xact_id(outer_arb_io_in_1_acquire_bits_client_xact_id),
    .io_in_1_acquire_bits_addr_beat(outer_arb_io_in_1_acquire_bits_addr_beat),
    .io_in_1_acquire_bits_is_builtin_type(outer_arb_io_in_1_acquire_bits_is_builtin_type),
    .io_in_1_acquire_bits_a_type(outer_arb_io_in_1_acquire_bits_a_type),
    .io_in_1_acquire_bits_union(outer_arb_io_in_1_acquire_bits_union),
    .io_in_1_acquire_bits_data(outer_arb_io_in_1_acquire_bits_data),
    .io_in_1_grant_ready(outer_arb_io_in_1_grant_ready),
    .io_in_1_grant_valid(outer_arb_io_in_1_grant_valid),
    .io_in_1_grant_bits_addr_beat(outer_arb_io_in_1_grant_bits_addr_beat),
    .io_in_1_grant_bits_client_xact_id(outer_arb_io_in_1_grant_bits_client_xact_id),
    .io_in_1_grant_bits_manager_xact_id(outer_arb_io_in_1_grant_bits_manager_xact_id),
    .io_in_1_grant_bits_is_builtin_type(outer_arb_io_in_1_grant_bits_is_builtin_type),
    .io_in_1_grant_bits_g_type(outer_arb_io_in_1_grant_bits_g_type),
    .io_in_1_grant_bits_data(outer_arb_io_in_1_grant_bits_data),
    .io_in_2_acquire_ready(outer_arb_io_in_2_acquire_ready),
    .io_in_2_acquire_valid(outer_arb_io_in_2_acquire_valid),
    .io_in_2_acquire_bits_addr_block(outer_arb_io_in_2_acquire_bits_addr_block),
    .io_in_2_acquire_bits_client_xact_id(outer_arb_io_in_2_acquire_bits_client_xact_id),
    .io_in_2_acquire_bits_addr_beat(outer_arb_io_in_2_acquire_bits_addr_beat),
    .io_in_2_acquire_bits_is_builtin_type(outer_arb_io_in_2_acquire_bits_is_builtin_type),
    .io_in_2_acquire_bits_a_type(outer_arb_io_in_2_acquire_bits_a_type),
    .io_in_2_acquire_bits_union(outer_arb_io_in_2_acquire_bits_union),
    .io_in_2_acquire_bits_data(outer_arb_io_in_2_acquire_bits_data),
    .io_in_2_grant_ready(outer_arb_io_in_2_grant_ready),
    .io_in_2_grant_valid(outer_arb_io_in_2_grant_valid),
    .io_in_2_grant_bits_addr_beat(outer_arb_io_in_2_grant_bits_addr_beat),
    .io_in_2_grant_bits_client_xact_id(outer_arb_io_in_2_grant_bits_client_xact_id),
    .io_in_2_grant_bits_manager_xact_id(outer_arb_io_in_2_grant_bits_manager_xact_id),
    .io_in_2_grant_bits_is_builtin_type(outer_arb_io_in_2_grant_bits_is_builtin_type),
    .io_in_2_grant_bits_g_type(outer_arb_io_in_2_grant_bits_g_type),
    .io_in_2_grant_bits_data(outer_arb_io_in_2_grant_bits_data),
    .io_in_3_acquire_ready(outer_arb_io_in_3_acquire_ready),
    .io_in_3_acquire_valid(outer_arb_io_in_3_acquire_valid),
    .io_in_3_acquire_bits_addr_block(outer_arb_io_in_3_acquire_bits_addr_block),
    .io_in_3_acquire_bits_client_xact_id(outer_arb_io_in_3_acquire_bits_client_xact_id),
    .io_in_3_acquire_bits_addr_beat(outer_arb_io_in_3_acquire_bits_addr_beat),
    .io_in_3_acquire_bits_is_builtin_type(outer_arb_io_in_3_acquire_bits_is_builtin_type),
    .io_in_3_acquire_bits_a_type(outer_arb_io_in_3_acquire_bits_a_type),
    .io_in_3_acquire_bits_union(outer_arb_io_in_3_acquire_bits_union),
    .io_in_3_acquire_bits_data(outer_arb_io_in_3_acquire_bits_data),
    .io_in_3_grant_ready(outer_arb_io_in_3_grant_ready),
    .io_in_3_grant_valid(outer_arb_io_in_3_grant_valid),
    .io_in_3_grant_bits_addr_beat(outer_arb_io_in_3_grant_bits_addr_beat),
    .io_in_3_grant_bits_client_xact_id(outer_arb_io_in_3_grant_bits_client_xact_id),
    .io_in_3_grant_bits_manager_xact_id(outer_arb_io_in_3_grant_bits_manager_xact_id),
    .io_in_3_grant_bits_is_builtin_type(outer_arb_io_in_3_grant_bits_is_builtin_type),
    .io_in_3_grant_bits_g_type(outer_arb_io_in_3_grant_bits_g_type),
    .io_in_3_grant_bits_data(outer_arb_io_in_3_grant_bits_data),
    .io_in_4_acquire_ready(outer_arb_io_in_4_acquire_ready),
    .io_in_4_acquire_valid(outer_arb_io_in_4_acquire_valid),
    .io_in_4_acquire_bits_addr_block(outer_arb_io_in_4_acquire_bits_addr_block),
    .io_in_4_acquire_bits_client_xact_id(outer_arb_io_in_4_acquire_bits_client_xact_id),
    .io_in_4_acquire_bits_addr_beat(outer_arb_io_in_4_acquire_bits_addr_beat),
    .io_in_4_acquire_bits_is_builtin_type(outer_arb_io_in_4_acquire_bits_is_builtin_type),
    .io_in_4_acquire_bits_a_type(outer_arb_io_in_4_acquire_bits_a_type),
    .io_in_4_acquire_bits_union(outer_arb_io_in_4_acquire_bits_union),
    .io_in_4_acquire_bits_data(outer_arb_io_in_4_acquire_bits_data),
    .io_in_4_grant_ready(outer_arb_io_in_4_grant_ready),
    .io_in_4_grant_valid(outer_arb_io_in_4_grant_valid),
    .io_in_4_grant_bits_addr_beat(outer_arb_io_in_4_grant_bits_addr_beat),
    .io_in_4_grant_bits_client_xact_id(outer_arb_io_in_4_grant_bits_client_xact_id),
    .io_in_4_grant_bits_manager_xact_id(outer_arb_io_in_4_grant_bits_manager_xact_id),
    .io_in_4_grant_bits_is_builtin_type(outer_arb_io_in_4_grant_bits_is_builtin_type),
    .io_in_4_grant_bits_g_type(outer_arb_io_in_4_grant_bits_g_type),
    .io_in_4_grant_bits_data(outer_arb_io_in_4_grant_bits_data),
    .io_out_acquire_ready(outer_arb_io_out_acquire_ready),
    .io_out_acquire_valid(outer_arb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(outer_arb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(outer_arb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(outer_arb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(outer_arb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(outer_arb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(outer_arb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(outer_arb_io_out_acquire_bits_data),
    .io_out_grant_ready(outer_arb_io_out_grant_ready),
    .io_out_grant_valid(outer_arb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(outer_arb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(outer_arb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(outer_arb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(outer_arb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(outer_arb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(outer_arb_io_out_grant_bits_data)
  );
  assign io_inner_acquire_ready = T_1723;
  assign io_inner_grant_valid = LockingRRArbiter_31_2320_io_out_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = LockingRRArbiter_31_2320_io_out_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = LockingRRArbiter_31_2320_io_out_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = LockingRRArbiter_31_2320_io_out_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = LockingRRArbiter_31_2320_io_out_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = LockingRRArbiter_31_2320_io_out_bits_client_id;
  assign io_inner_finish_ready = GEN_2;
  assign io_inner_probe_valid = LockingRRArbiter_32_2321_io_out_valid;
  assign io_inner_probe_bits_addr_block = LockingRRArbiter_32_2321_io_out_bits_addr_block;
  assign io_inner_probe_bits_p_type = LockingRRArbiter_32_2321_io_out_bits_p_type;
  assign io_inner_probe_bits_client_id = LockingRRArbiter_32_2321_io_out_bits_client_id;
  assign io_inner_release_ready = T_2292;
  assign io_outer_acquire_valid = outer_arb_io_out_acquire_valid;
  assign io_outer_acquire_bits_addr_block = outer_arb_io_out_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_arb_io_out_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = outer_arb_io_out_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = outer_arb_io_out_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = outer_arb_io_out_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = outer_arb_io_out_acquire_bits_union;
  assign io_outer_acquire_bits_data = T_2507;
  assign io_outer_grant_ready = outer_arb_io_out_grant_ready;
  assign BroadcastVoluntaryReleaseTracker_1051_clk = clk;
  assign BroadcastVoluntaryReleaseTracker_1051_reset = reset;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_valid = T_1725;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_data = T_1297;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_ready = LockingRRArbiter_31_2320_io_in_0_ready;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_valid = T_2324;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_ready = LockingRRArbiter_32_2321_io_in_0_ready;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_valid = io_inner_release_valid;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_data = T_1869;
  assign BroadcastVoluntaryReleaseTracker_1051_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_incoherent_0 = io_incoherent_0;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_ready = outer_arb_io_in_0_acquire_ready;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_valid = outer_arb_io_in_0_grant_valid;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_addr_beat = outer_arb_io_in_0_grant_bits_addr_beat;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_client_xact_id = outer_arb_io_in_0_grant_bits_client_xact_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_0_grant_bits_manager_xact_id;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_0_grant_bits_is_builtin_type;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_g_type = outer_arb_io_in_0_grant_bits_g_type;
  assign BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_bits_data = outer_arb_io_in_0_grant_bits_data;
  assign BroadcastVoluntaryReleaseTracker_1051_io_alloc_iacq = T_1728;
  assign BroadcastVoluntaryReleaseTracker_1051_io_alloc_irel = T_2298;
  assign BroadcastVoluntaryReleaseTracker_1051_io_alloc_oprb = GEN_13;
  assign BroadcastAcquireTracker_1052_clk = clk;
  assign BroadcastAcquireTracker_1052_reset = reset;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_valid = T_1725;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_data = T_1390;
  assign BroadcastAcquireTracker_1052_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BroadcastAcquireTracker_1052_io_inner_grant_ready = LockingRRArbiter_31_2320_io_in_1_ready;
  assign BroadcastAcquireTracker_1052_io_inner_finish_valid = T_2327;
  assign BroadcastAcquireTracker_1052_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BroadcastAcquireTracker_1052_io_inner_probe_ready = LockingRRArbiter_32_2321_io_in_1_ready;
  assign BroadcastAcquireTracker_1052_io_inner_release_valid = io_inner_release_valid;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_data = T_1962;
  assign BroadcastAcquireTracker_1052_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BroadcastAcquireTracker_1052_io_incoherent_0 = io_incoherent_0;
  assign BroadcastAcquireTracker_1052_io_outer_acquire_ready = outer_arb_io_in_1_acquire_ready;
  assign BroadcastAcquireTracker_1052_io_outer_grant_valid = outer_arb_io_in_1_grant_valid;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_addr_beat = outer_arb_io_in_1_grant_bits_addr_beat;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_client_xact_id = outer_arb_io_in_1_grant_bits_client_xact_id;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_1_grant_bits_manager_xact_id;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_1_grant_bits_is_builtin_type;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_g_type = outer_arb_io_in_1_grant_bits_g_type;
  assign BroadcastAcquireTracker_1052_io_outer_grant_bits_data = outer_arb_io_in_1_grant_bits_data;
  assign BroadcastAcquireTracker_1052_io_alloc_iacq = T_1733;
  assign BroadcastAcquireTracker_1052_io_alloc_irel = T_2303;
  assign BroadcastAcquireTracker_1052_io_alloc_oprb = GEN_31;
  assign BroadcastAcquireTracker_28_1053_clk = clk;
  assign BroadcastAcquireTracker_28_1053_reset = reset;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_valid = T_1725;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_data = T_1483;
  assign BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BroadcastAcquireTracker_28_1053_io_inner_grant_ready = LockingRRArbiter_31_2320_io_in_2_ready;
  assign BroadcastAcquireTracker_28_1053_io_inner_finish_valid = T_2330;
  assign BroadcastAcquireTracker_28_1053_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BroadcastAcquireTracker_28_1053_io_inner_probe_ready = LockingRRArbiter_32_2321_io_in_2_ready;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_valid = io_inner_release_valid;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_data = T_2055;
  assign BroadcastAcquireTracker_28_1053_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BroadcastAcquireTracker_28_1053_io_incoherent_0 = io_incoherent_0;
  assign BroadcastAcquireTracker_28_1053_io_outer_acquire_ready = outer_arb_io_in_2_acquire_ready;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_valid = outer_arb_io_in_2_grant_valid;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_addr_beat = outer_arb_io_in_2_grant_bits_addr_beat;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_client_xact_id = outer_arb_io_in_2_grant_bits_client_xact_id;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_2_grant_bits_manager_xact_id;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_2_grant_bits_is_builtin_type;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_g_type = outer_arb_io_in_2_grant_bits_g_type;
  assign BroadcastAcquireTracker_28_1053_io_outer_grant_bits_data = outer_arb_io_in_2_grant_bits_data;
  assign BroadcastAcquireTracker_28_1053_io_alloc_iacq = T_1738;
  assign BroadcastAcquireTracker_28_1053_io_alloc_irel = T_2308;
  assign BroadcastAcquireTracker_28_1053_io_alloc_oprb = GEN_65;
  assign BroadcastAcquireTracker_29_1054_clk = clk;
  assign BroadcastAcquireTracker_29_1054_reset = reset;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_valid = T_1725;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_data = T_1576;
  assign BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BroadcastAcquireTracker_29_1054_io_inner_grant_ready = LockingRRArbiter_31_2320_io_in_3_ready;
  assign BroadcastAcquireTracker_29_1054_io_inner_finish_valid = T_2333;
  assign BroadcastAcquireTracker_29_1054_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BroadcastAcquireTracker_29_1054_io_inner_probe_ready = LockingRRArbiter_32_2321_io_in_3_ready;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_valid = io_inner_release_valid;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_data = T_2148;
  assign BroadcastAcquireTracker_29_1054_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BroadcastAcquireTracker_29_1054_io_incoherent_0 = io_incoherent_0;
  assign BroadcastAcquireTracker_29_1054_io_outer_acquire_ready = outer_arb_io_in_3_acquire_ready;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_valid = outer_arb_io_in_3_grant_valid;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_addr_beat = outer_arb_io_in_3_grant_bits_addr_beat;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_client_xact_id = outer_arb_io_in_3_grant_bits_client_xact_id;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_3_grant_bits_manager_xact_id;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_3_grant_bits_is_builtin_type;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_g_type = outer_arb_io_in_3_grant_bits_g_type;
  assign BroadcastAcquireTracker_29_1054_io_outer_grant_bits_data = outer_arb_io_in_3_grant_bits_data;
  assign BroadcastAcquireTracker_29_1054_io_alloc_iacq = T_1743;
  assign BroadcastAcquireTracker_29_1054_io_alloc_irel = T_2313;
  assign BroadcastAcquireTracker_29_1054_io_alloc_oprb = GEN_66;
  assign BroadcastAcquireTracker_30_1055_clk = clk;
  assign BroadcastAcquireTracker_30_1055_reset = reset;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_valid = T_1725;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_union = io_inner_acquire_bits_union;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_data = T_1669;
  assign BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_client_id = io_inner_acquire_bits_client_id;
  assign BroadcastAcquireTracker_30_1055_io_inner_grant_ready = LockingRRArbiter_31_2320_io_in_4_ready;
  assign BroadcastAcquireTracker_30_1055_io_inner_finish_valid = T_2336;
  assign BroadcastAcquireTracker_30_1055_io_inner_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign BroadcastAcquireTracker_30_1055_io_inner_probe_ready = LockingRRArbiter_32_2321_io_in_4_ready;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_valid = io_inner_release_valid;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_r_type = io_inner_release_bits_r_type;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_data = T_2241;
  assign BroadcastAcquireTracker_30_1055_io_inner_release_bits_client_id = io_inner_release_bits_client_id;
  assign BroadcastAcquireTracker_30_1055_io_incoherent_0 = io_incoherent_0;
  assign BroadcastAcquireTracker_30_1055_io_outer_acquire_ready = outer_arb_io_in_4_acquire_ready;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_valid = outer_arb_io_in_4_grant_valid;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_addr_beat = outer_arb_io_in_4_grant_bits_addr_beat;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_client_xact_id = outer_arb_io_in_4_grant_bits_client_xact_id;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_manager_xact_id = outer_arb_io_in_4_grant_bits_manager_xact_id;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_is_builtin_type = outer_arb_io_in_4_grant_bits_is_builtin_type;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_g_type = outer_arb_io_in_4_grant_bits_g_type;
  assign BroadcastAcquireTracker_30_1055_io_outer_grant_bits_data = outer_arb_io_in_4_grant_bits_data;
  assign BroadcastAcquireTracker_30_1055_io_alloc_iacq = T_1748;
  assign BroadcastAcquireTracker_30_1055_io_alloc_irel = T_2318;
  assign BroadcastAcquireTracker_30_1055_io_alloc_oprb = GEN_67;
  assign T_1063 = ~ sdq_val;
  assign T_1064 = T_1063[0];
  assign T_1065 = T_1063[1];
  assign T_1066 = T_1063[2];
  assign T_1067 = T_1063[3];
  assign T_1068 = T_1063[4];
  assign T_1069 = T_1063[5];
  assign T_1070 = T_1063[6];
  assign T_1071 = T_1063[7];
  assign T_1080 = T_1070 ? 3'h6 : 3'h7;
  assign T_1081 = T_1069 ? 3'h5 : T_1080;
  assign T_1082 = T_1068 ? 3'h4 : T_1081;
  assign T_1083 = T_1067 ? {{1'd0}, 2'h3} : T_1082;
  assign T_1084 = T_1066 ? {{1'd0}, 2'h2} : T_1083;
  assign T_1085 = T_1065 ? {{2'd0}, 1'h1} : T_1084;
  assign sdq_alloc_id = T_1064 ? {{2'd0}, 1'h0} : T_1085;
  assign GEN_59 = {{7'd0}, 1'h0};
  assign T_1088 = T_1063 == GEN_59;
  assign sdq_rdy = T_1088 == 1'h0;
  assign T_1090 = BroadcastVoluntaryReleaseTracker_1051_io_alloc_iacq | BroadcastVoluntaryReleaseTracker_1051_io_matches_iacq;
  assign T_1091 = BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_ready & BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_valid;
  assign T_1092 = T_1090 & T_1091;
  assign T_1101_0 = 3'h2;
  assign T_1101_1 = 3'h3;
  assign T_1101_2 = 3'h4;
  assign T_1103 = T_1101_0 == BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type;
  assign T_1104 = T_1101_1 == BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type;
  assign T_1105 = T_1101_2 == BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_a_type;
  assign T_1108 = T_1103 | T_1104;
  assign T_1109 = T_1108 | T_1105;
  assign T_1110 = BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_bits_is_builtin_type & T_1109;
  assign T_1111 = T_1092 & T_1110;
  assign T_1112 = BroadcastAcquireTracker_1052_io_alloc_iacq | BroadcastAcquireTracker_1052_io_matches_iacq;
  assign T_1113 = BroadcastAcquireTracker_1052_io_inner_acquire_ready & BroadcastAcquireTracker_1052_io_inner_acquire_valid;
  assign T_1114 = T_1112 & T_1113;
  assign T_1123_0 = 3'h2;
  assign T_1123_1 = 3'h3;
  assign T_1123_2 = 3'h4;
  assign T_1125 = T_1123_0 == BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type;
  assign T_1126 = T_1123_1 == BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type;
  assign T_1127 = T_1123_2 == BroadcastAcquireTracker_1052_io_inner_acquire_bits_a_type;
  assign T_1130 = T_1125 | T_1126;
  assign T_1131 = T_1130 | T_1127;
  assign T_1132 = BroadcastAcquireTracker_1052_io_inner_acquire_bits_is_builtin_type & T_1131;
  assign T_1133 = T_1114 & T_1132;
  assign T_1134 = BroadcastAcquireTracker_28_1053_io_alloc_iacq | BroadcastAcquireTracker_28_1053_io_matches_iacq;
  assign T_1135 = BroadcastAcquireTracker_28_1053_io_inner_acquire_ready & BroadcastAcquireTracker_28_1053_io_inner_acquire_valid;
  assign T_1136 = T_1134 & T_1135;
  assign T_1145_0 = 3'h2;
  assign T_1145_1 = 3'h3;
  assign T_1145_2 = 3'h4;
  assign T_1147 = T_1145_0 == BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type;
  assign T_1148 = T_1145_1 == BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type;
  assign T_1149 = T_1145_2 == BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_a_type;
  assign T_1152 = T_1147 | T_1148;
  assign T_1153 = T_1152 | T_1149;
  assign T_1154 = BroadcastAcquireTracker_28_1053_io_inner_acquire_bits_is_builtin_type & T_1153;
  assign T_1155 = T_1136 & T_1154;
  assign T_1156 = BroadcastAcquireTracker_29_1054_io_alloc_iacq | BroadcastAcquireTracker_29_1054_io_matches_iacq;
  assign T_1157 = BroadcastAcquireTracker_29_1054_io_inner_acquire_ready & BroadcastAcquireTracker_29_1054_io_inner_acquire_valid;
  assign T_1158 = T_1156 & T_1157;
  assign T_1167_0 = 3'h2;
  assign T_1167_1 = 3'h3;
  assign T_1167_2 = 3'h4;
  assign T_1169 = T_1167_0 == BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type;
  assign T_1170 = T_1167_1 == BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type;
  assign T_1171 = T_1167_2 == BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_a_type;
  assign T_1174 = T_1169 | T_1170;
  assign T_1175 = T_1174 | T_1171;
  assign T_1176 = BroadcastAcquireTracker_29_1054_io_inner_acquire_bits_is_builtin_type & T_1175;
  assign T_1177 = T_1158 & T_1176;
  assign T_1178 = BroadcastAcquireTracker_30_1055_io_alloc_iacq | BroadcastAcquireTracker_30_1055_io_matches_iacq;
  assign T_1179 = BroadcastAcquireTracker_30_1055_io_inner_acquire_ready & BroadcastAcquireTracker_30_1055_io_inner_acquire_valid;
  assign T_1180 = T_1178 & T_1179;
  assign T_1189_0 = 3'h2;
  assign T_1189_1 = 3'h3;
  assign T_1189_2 = 3'h4;
  assign T_1191 = T_1189_0 == BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type;
  assign T_1192 = T_1189_1 == BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type;
  assign T_1193 = T_1189_2 == BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_a_type;
  assign T_1196 = T_1191 | T_1192;
  assign T_1197 = T_1196 | T_1193;
  assign T_1198 = BroadcastAcquireTracker_30_1055_io_inner_acquire_bits_is_builtin_type & T_1197;
  assign T_1199 = T_1180 & T_1198;
  assign T_1200 = T_1111 | T_1133;
  assign T_1201 = T_1200 | T_1155;
  assign T_1202 = T_1201 | T_1177;
  assign sdq_enq = T_1202 | T_1199;
  assign GEN_0 = io_inner_acquire_bits_data;
  assign GEN_60 = {{2'd0}, 1'h0};
  assign GEN_5 = GEN_60 == sdq_alloc_id ? GEN_0 : sdq_0;
  assign GEN_61 = {{2'd0}, 1'h1};
  assign GEN_6 = GEN_61 == sdq_alloc_id ? GEN_0 : sdq_1;
  assign GEN_62 = {{1'd0}, 2'h2};
  assign GEN_7 = GEN_62 == sdq_alloc_id ? GEN_0 : sdq_2;
  assign GEN_63 = {{1'd0}, 2'h3};
  assign GEN_8 = GEN_63 == sdq_alloc_id ? GEN_0 : sdq_3;
  assign GEN_9 = 3'h4 == sdq_alloc_id ? GEN_0 : sdq_4;
  assign GEN_10 = 3'h5 == sdq_alloc_id ? GEN_0 : sdq_5;
  assign GEN_11 = 3'h6 == sdq_alloc_id ? GEN_0 : sdq_6;
  assign GEN_12 = 3'h7 == sdq_alloc_id ? GEN_0 : sdq_7;
  assign GEN_14 = sdq_enq ? GEN_5 : sdq_0;
  assign GEN_15 = sdq_enq ? GEN_6 : sdq_1;
  assign GEN_16 = sdq_enq ? GEN_7 : sdq_2;
  assign GEN_17 = sdq_enq ? GEN_8 : sdq_3;
  assign GEN_18 = sdq_enq ? GEN_9 : sdq_4;
  assign GEN_19 = sdq_enq ? GEN_10 : sdq_5;
  assign GEN_20 = sdq_enq ? GEN_11 : sdq_6;
  assign GEN_21 = sdq_enq ? GEN_12 : sdq_7;
  assign T_1203 = io_inner_acquire_valid & io_inner_release_valid;
  assign T_1204 = io_inner_release_bits_addr_block == io_inner_acquire_bits_addr_block;
  assign irel_vs_iacq_conflict = T_1203 & T_1204;
  assign T_1251_idx = sdq_alloc_id;
  assign T_1251_loc = 2'h0;
  assign T_1297 = {T_1251_idx,T_1251_loc};
  assign T_1344_idx = sdq_alloc_id;
  assign T_1344_loc = 2'h0;
  assign T_1390 = {T_1344_idx,T_1344_loc};
  assign T_1437_idx = sdq_alloc_id;
  assign T_1437_loc = 2'h0;
  assign T_1483 = {T_1437_idx,T_1437_loc};
  assign T_1530_idx = sdq_alloc_id;
  assign T_1530_loc = 2'h0;
  assign T_1576 = {T_1530_idx,T_1530_loc};
  assign T_1623_idx = sdq_alloc_id;
  assign T_1623_loc = 2'h0;
  assign T_1669 = {T_1623_idx,T_1623_loc};
  assign T_1671 = irel_vs_iacq_conflict == 1'h0;
  assign T_1672 = sdq_rdy & T_1671;
  assign T_1678_0 = BroadcastVoluntaryReleaseTracker_1051_io_inner_acquire_ready;
  assign T_1678_1 = BroadcastAcquireTracker_1052_io_inner_acquire_ready;
  assign T_1678_2 = BroadcastAcquireTracker_28_1053_io_inner_acquire_ready;
  assign T_1678_3 = BroadcastAcquireTracker_29_1054_io_inner_acquire_ready;
  assign T_1678_4 = BroadcastAcquireTracker_30_1055_io_inner_acquire_ready;
  assign T_1680 = {T_1678_1,T_1678_0};
  assign T_1681 = {T_1678_4,T_1678_3};
  assign T_1682 = {T_1681,T_1678_2};
  assign T_1683 = {T_1682,T_1680};
  assign T_1684 = T_1683[0];
  assign T_1685 = T_1683[1];
  assign T_1686 = T_1683[2];
  assign T_1687 = T_1683[3];
  assign T_1688 = T_1683[4];
  assign T_1696 = T_1688 ? 5'h10 : 5'h0;
  assign T_1697 = T_1687 ? 5'h8 : T_1696;
  assign T_1698 = T_1686 ? 5'h4 : T_1697;
  assign T_1699 = T_1685 ? 5'h2 : T_1698;
  assign T_1700 = T_1684 ? 5'h1 : T_1699;
  assign T_1706_0 = BroadcastVoluntaryReleaseTracker_1051_io_matches_iacq;
  assign T_1706_1 = BroadcastAcquireTracker_1052_io_matches_iacq;
  assign T_1706_2 = BroadcastAcquireTracker_28_1053_io_matches_iacq;
  assign T_1706_3 = BroadcastAcquireTracker_29_1054_io_matches_iacq;
  assign T_1706_4 = BroadcastAcquireTracker_30_1055_io_matches_iacq;
  assign T_1708 = {T_1706_1,T_1706_0};
  assign T_1709 = {T_1706_4,T_1706_3};
  assign T_1710 = {T_1709,T_1706_2};
  assign T_1711 = {T_1710,T_1708};
  assign GEN_64 = {{4'd0}, 1'h0};
  assign T_1713 = T_1711 != GEN_64;
  assign T_1715 = T_1713 == 1'h0;
  assign T_1717 = T_1683 != GEN_64;
  assign T_1718 = T_1711 & T_1683;
  assign T_1720 = T_1718 != GEN_64;
  assign T_1721 = T_1715 ? T_1717 : T_1720;
  assign T_1722 = T_1721 & T_1672;
  assign T_1723 = T_1722 & sdq_rdy;
  assign T_1724 = io_inner_acquire_valid & sdq_rdy;
  assign T_1725 = T_1724 & T_1672;
  assign T_1726 = T_1700[0];
  assign T_1727 = T_1726 & T_1715;
  assign T_1728 = T_1727 & T_1672;
  assign T_1731 = T_1700[1];
  assign T_1732 = T_1731 & T_1715;
  assign T_1733 = T_1732 & T_1672;
  assign T_1736 = T_1700[2];
  assign T_1737 = T_1736 & T_1715;
  assign T_1738 = T_1737 & T_1672;
  assign T_1741 = T_1700[3];
  assign T_1742 = T_1741 & T_1715;
  assign T_1743 = T_1742 & T_1672;
  assign T_1746 = T_1700[4];
  assign T_1747 = T_1746 & T_1715;
  assign T_1748 = T_1747 & T_1672;
  assign T_1749 = io_inner_release_ready & io_inner_release_valid;
  assign T_1750 = T_1749 & io_inner_release_bits_voluntary;
  assign T_1756_0 = 3'h0;
  assign T_1756_1 = 3'h1;
  assign T_1756_2 = 3'h2;
  assign T_1758 = T_1756_0 == io_inner_release_bits_r_type;
  assign T_1759 = T_1756_1 == io_inner_release_bits_r_type;
  assign T_1760 = T_1756_2 == io_inner_release_bits_r_type;
  assign T_1763 = T_1758 | T_1759;
  assign T_1764 = T_1763 | T_1760;
  assign vwbdq_enq = T_1750 & T_1764;
  assign T_1769 = rel_data_cnt + GEN_61;
  assign T_1770 = T_1769[2:0];
  assign GEN_22 = vwbdq_enq ? T_1770 : rel_data_cnt;
  assign GEN_1 = io_inner_release_bits_data;
  assign GEN_23 = GEN_60 == rel_data_cnt ? GEN_1 : vwbdq_0;
  assign GEN_24 = GEN_61 == rel_data_cnt ? GEN_1 : vwbdq_1;
  assign GEN_25 = GEN_62 == rel_data_cnt ? GEN_1 : vwbdq_2;
  assign GEN_26 = GEN_63 == rel_data_cnt ? GEN_1 : vwbdq_3;
  assign GEN_27 = 3'h4 == rel_data_cnt ? GEN_1 : vwbdq_4;
  assign GEN_28 = 3'h5 == rel_data_cnt ? GEN_1 : vwbdq_5;
  assign GEN_29 = 3'h6 == rel_data_cnt ? GEN_1 : vwbdq_6;
  assign GEN_30 = 3'h7 == rel_data_cnt ? GEN_1 : vwbdq_7;
  assign GEN_32 = vwbdq_enq ? GEN_23 : vwbdq_0;
  assign GEN_33 = vwbdq_enq ? GEN_24 : vwbdq_1;
  assign GEN_34 = vwbdq_enq ? GEN_25 : vwbdq_2;
  assign GEN_35 = vwbdq_enq ? GEN_26 : vwbdq_3;
  assign GEN_36 = vwbdq_enq ? GEN_27 : vwbdq_4;
  assign GEN_37 = vwbdq_enq ? GEN_28 : vwbdq_5;
  assign GEN_38 = vwbdq_enq ? GEN_29 : vwbdq_6;
  assign GEN_39 = vwbdq_enq ? GEN_30 : vwbdq_7;
  assign T_1823_idx = rel_data_cnt;
  assign T_1823_loc = 2'h1;
  assign T_1869 = {T_1823_idx,T_1823_loc};
  assign T_1916_idx = rel_data_cnt;
  assign T_1916_loc = 2'h2;
  assign T_1962 = {T_1916_idx,T_1916_loc};
  assign T_2009_idx = rel_data_cnt;
  assign T_2009_loc = 2'h2;
  assign T_2055 = {T_2009_idx,T_2009_loc};
  assign T_2102_idx = rel_data_cnt;
  assign T_2102_loc = 2'h2;
  assign T_2148 = {T_2102_idx,T_2102_loc};
  assign T_2195_idx = rel_data_cnt;
  assign T_2195_loc = 2'h2;
  assign T_2241 = {T_2195_idx,T_2195_loc};
  assign T_2247_0 = BroadcastVoluntaryReleaseTracker_1051_io_inner_release_ready;
  assign T_2247_1 = BroadcastAcquireTracker_1052_io_inner_release_ready;
  assign T_2247_2 = BroadcastAcquireTracker_28_1053_io_inner_release_ready;
  assign T_2247_3 = BroadcastAcquireTracker_29_1054_io_inner_release_ready;
  assign T_2247_4 = BroadcastAcquireTracker_30_1055_io_inner_release_ready;
  assign T_2249 = {T_2247_1,T_2247_0};
  assign T_2250 = {T_2247_4,T_2247_3};
  assign T_2251 = {T_2250,T_2247_2};
  assign T_2252 = {T_2251,T_2249};
  assign T_2253 = T_2252[0];
  assign T_2254 = T_2252[1];
  assign T_2255 = T_2252[2];
  assign T_2256 = T_2252[3];
  assign T_2257 = T_2252[4];
  assign T_2265 = T_2257 ? 5'h10 : 5'h0;
  assign T_2266 = T_2256 ? 5'h8 : T_2265;
  assign T_2267 = T_2255 ? 5'h4 : T_2266;
  assign T_2268 = T_2254 ? 5'h2 : T_2267;
  assign T_2269 = T_2253 ? 5'h1 : T_2268;
  assign T_2275_0 = BroadcastVoluntaryReleaseTracker_1051_io_matches_irel;
  assign T_2275_1 = BroadcastAcquireTracker_1052_io_matches_irel;
  assign T_2275_2 = BroadcastAcquireTracker_28_1053_io_matches_irel;
  assign T_2275_3 = BroadcastAcquireTracker_29_1054_io_matches_irel;
  assign T_2275_4 = BroadcastAcquireTracker_30_1055_io_matches_irel;
  assign T_2277 = {T_2275_1,T_2275_0};
  assign T_2278 = {T_2275_4,T_2275_3};
  assign T_2279 = {T_2278,T_2275_2};
  assign T_2280 = {T_2279,T_2277};
  assign T_2282 = T_2280 != GEN_64;
  assign T_2284 = T_2282 == 1'h0;
  assign T_2288 = T_2252 != GEN_64;
  assign T_2289 = T_2280 & T_2252;
  assign T_2291 = T_2289 != GEN_64;
  assign T_2292 = T_2284 ? T_2288 : T_2291;
  assign T_2297 = T_2269[0];
  assign T_2298 = T_2297 & T_2284;
  assign T_2302 = T_2269[1];
  assign T_2303 = T_2302 & T_2284;
  assign T_2307 = T_2269[2];
  assign T_2308 = T_2307 & T_2284;
  assign T_2312 = T_2269[3];
  assign T_2313 = T_2312 & T_2284;
  assign T_2317 = T_2269[4];
  assign T_2318 = T_2317 & T_2284;
  assign LockingRRArbiter_31_2320_clk = clk;
  assign LockingRRArbiter_31_2320_reset = reset;
  assign LockingRRArbiter_31_2320_io_in_0_valid = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_valid;
  assign LockingRRArbiter_31_2320_io_in_0_bits_addr_beat = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_31_2320_io_in_0_bits_client_xact_id = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_31_2320_io_in_0_bits_manager_xact_id = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_31_2320_io_in_0_bits_is_builtin_type = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_31_2320_io_in_0_bits_g_type = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_31_2320_io_in_0_bits_data = {{59'd0}, BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_data};
  assign LockingRRArbiter_31_2320_io_in_0_bits_client_id = BroadcastVoluntaryReleaseTracker_1051_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_31_2320_io_in_1_valid = BroadcastAcquireTracker_1052_io_inner_grant_valid;
  assign LockingRRArbiter_31_2320_io_in_1_bits_addr_beat = BroadcastAcquireTracker_1052_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_31_2320_io_in_1_bits_client_xact_id = BroadcastAcquireTracker_1052_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_31_2320_io_in_1_bits_manager_xact_id = BroadcastAcquireTracker_1052_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_31_2320_io_in_1_bits_is_builtin_type = BroadcastAcquireTracker_1052_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_31_2320_io_in_1_bits_g_type = BroadcastAcquireTracker_1052_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_31_2320_io_in_1_bits_data = {{59'd0}, BroadcastAcquireTracker_1052_io_inner_grant_bits_data};
  assign LockingRRArbiter_31_2320_io_in_1_bits_client_id = BroadcastAcquireTracker_1052_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_31_2320_io_in_2_valid = BroadcastAcquireTracker_28_1053_io_inner_grant_valid;
  assign LockingRRArbiter_31_2320_io_in_2_bits_addr_beat = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_31_2320_io_in_2_bits_client_xact_id = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_31_2320_io_in_2_bits_manager_xact_id = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_31_2320_io_in_2_bits_is_builtin_type = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_31_2320_io_in_2_bits_g_type = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_31_2320_io_in_2_bits_data = {{59'd0}, BroadcastAcquireTracker_28_1053_io_inner_grant_bits_data};
  assign LockingRRArbiter_31_2320_io_in_2_bits_client_id = BroadcastAcquireTracker_28_1053_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_31_2320_io_in_3_valid = BroadcastAcquireTracker_29_1054_io_inner_grant_valid;
  assign LockingRRArbiter_31_2320_io_in_3_bits_addr_beat = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_31_2320_io_in_3_bits_client_xact_id = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_31_2320_io_in_3_bits_manager_xact_id = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_31_2320_io_in_3_bits_is_builtin_type = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_31_2320_io_in_3_bits_g_type = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_31_2320_io_in_3_bits_data = {{59'd0}, BroadcastAcquireTracker_29_1054_io_inner_grant_bits_data};
  assign LockingRRArbiter_31_2320_io_in_3_bits_client_id = BroadcastAcquireTracker_29_1054_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_31_2320_io_in_4_valid = BroadcastAcquireTracker_30_1055_io_inner_grant_valid;
  assign LockingRRArbiter_31_2320_io_in_4_bits_addr_beat = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_addr_beat;
  assign LockingRRArbiter_31_2320_io_in_4_bits_client_xact_id = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_xact_id;
  assign LockingRRArbiter_31_2320_io_in_4_bits_manager_xact_id = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_manager_xact_id;
  assign LockingRRArbiter_31_2320_io_in_4_bits_is_builtin_type = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_is_builtin_type;
  assign LockingRRArbiter_31_2320_io_in_4_bits_g_type = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_g_type;
  assign LockingRRArbiter_31_2320_io_in_4_bits_data = {{59'd0}, BroadcastAcquireTracker_30_1055_io_inner_grant_bits_data};
  assign LockingRRArbiter_31_2320_io_in_4_bits_client_id = BroadcastAcquireTracker_30_1055_io_inner_grant_bits_client_id;
  assign LockingRRArbiter_31_2320_io_out_ready = io_inner_grant_ready;
  assign LockingRRArbiter_32_2321_clk = clk;
  assign LockingRRArbiter_32_2321_reset = reset;
  assign LockingRRArbiter_32_2321_io_in_0_valid = BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_valid;
  assign LockingRRArbiter_32_2321_io_in_0_bits_addr_block = BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_32_2321_io_in_0_bits_p_type = BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_32_2321_io_in_0_bits_client_id = BroadcastVoluntaryReleaseTracker_1051_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_32_2321_io_in_1_valid = BroadcastAcquireTracker_1052_io_inner_probe_valid;
  assign LockingRRArbiter_32_2321_io_in_1_bits_addr_block = BroadcastAcquireTracker_1052_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_32_2321_io_in_1_bits_p_type = BroadcastAcquireTracker_1052_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_32_2321_io_in_1_bits_client_id = BroadcastAcquireTracker_1052_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_32_2321_io_in_2_valid = BroadcastAcquireTracker_28_1053_io_inner_probe_valid;
  assign LockingRRArbiter_32_2321_io_in_2_bits_addr_block = BroadcastAcquireTracker_28_1053_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_32_2321_io_in_2_bits_p_type = BroadcastAcquireTracker_28_1053_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_32_2321_io_in_2_bits_client_id = BroadcastAcquireTracker_28_1053_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_32_2321_io_in_3_valid = BroadcastAcquireTracker_29_1054_io_inner_probe_valid;
  assign LockingRRArbiter_32_2321_io_in_3_bits_addr_block = BroadcastAcquireTracker_29_1054_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_32_2321_io_in_3_bits_p_type = BroadcastAcquireTracker_29_1054_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_32_2321_io_in_3_bits_client_id = BroadcastAcquireTracker_29_1054_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_32_2321_io_in_4_valid = BroadcastAcquireTracker_30_1055_io_inner_probe_valid;
  assign LockingRRArbiter_32_2321_io_in_4_bits_addr_block = BroadcastAcquireTracker_30_1055_io_inner_probe_bits_addr_block;
  assign LockingRRArbiter_32_2321_io_in_4_bits_p_type = BroadcastAcquireTracker_30_1055_io_inner_probe_bits_p_type;
  assign LockingRRArbiter_32_2321_io_in_4_bits_client_id = BroadcastAcquireTracker_30_1055_io_inner_probe_bits_client_id;
  assign LockingRRArbiter_32_2321_io_out_ready = io_inner_probe_ready;
  assign T_2323 = io_inner_finish_bits_manager_xact_id == GEN_60;
  assign T_2324 = io_inner_finish_valid & T_2323;
  assign T_2326 = io_inner_finish_bits_manager_xact_id == GEN_61;
  assign T_2327 = io_inner_finish_valid & T_2326;
  assign T_2329 = io_inner_finish_bits_manager_xact_id == GEN_62;
  assign T_2330 = io_inner_finish_valid & T_2329;
  assign T_2332 = io_inner_finish_bits_manager_xact_id == GEN_63;
  assign T_2333 = io_inner_finish_valid & T_2332;
  assign T_2335 = io_inner_finish_bits_manager_xact_id == 3'h4;
  assign T_2336 = io_inner_finish_valid & T_2335;
  assign T_2342_0 = BroadcastVoluntaryReleaseTracker_1051_io_inner_finish_ready;
  assign T_2342_1 = BroadcastAcquireTracker_1052_io_inner_finish_ready;
  assign T_2342_2 = BroadcastAcquireTracker_28_1053_io_inner_finish_ready;
  assign T_2342_3 = BroadcastAcquireTracker_29_1054_io_inner_finish_ready;
  assign T_2342_4 = BroadcastAcquireTracker_30_1055_io_inner_finish_ready;
  assign GEN_2 = GEN_43;
  assign GEN_40 = GEN_61 == io_inner_finish_bits_manager_xact_id ? T_2342_1 : T_2342_0;
  assign GEN_41 = GEN_62 == io_inner_finish_bits_manager_xact_id ? T_2342_2 : GEN_40;
  assign GEN_42 = GEN_63 == io_inner_finish_bits_manager_xact_id ? T_2342_3 : GEN_41;
  assign GEN_43 = 3'h4 == io_inner_finish_bits_manager_xact_id ? T_2342_4 : GEN_42;
  assign outer_arb_clk = clk;
  assign outer_arb_reset = reset;
  assign outer_arb_io_in_0_acquire_valid = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_valid;
  assign outer_arb_io_in_0_acquire_bits_addr_block = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_0_acquire_bits_client_xact_id = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_0_acquire_bits_addr_beat = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_0_acquire_bits_is_builtin_type = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_0_acquire_bits_a_type = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_0_acquire_bits_union = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_union;
  assign outer_arb_io_in_0_acquire_bits_data = BroadcastVoluntaryReleaseTracker_1051_io_outer_acquire_bits_data;
  assign outer_arb_io_in_0_grant_ready = BroadcastVoluntaryReleaseTracker_1051_io_outer_grant_ready;
  assign outer_arb_io_in_1_acquire_valid = BroadcastAcquireTracker_1052_io_outer_acquire_valid;
  assign outer_arb_io_in_1_acquire_bits_addr_block = BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_1_acquire_bits_client_xact_id = BroadcastAcquireTracker_1052_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_1_acquire_bits_addr_beat = BroadcastAcquireTracker_1052_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_1_acquire_bits_is_builtin_type = BroadcastAcquireTracker_1052_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_1_acquire_bits_a_type = BroadcastAcquireTracker_1052_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_1_acquire_bits_union = BroadcastAcquireTracker_1052_io_outer_acquire_bits_union;
  assign outer_arb_io_in_1_acquire_bits_data = BroadcastAcquireTracker_1052_io_outer_acquire_bits_data;
  assign outer_arb_io_in_1_grant_ready = BroadcastAcquireTracker_1052_io_outer_grant_ready;
  assign outer_arb_io_in_2_acquire_valid = BroadcastAcquireTracker_28_1053_io_outer_acquire_valid;
  assign outer_arb_io_in_2_acquire_bits_addr_block = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_2_acquire_bits_client_xact_id = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_2_acquire_bits_addr_beat = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_2_acquire_bits_is_builtin_type = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_2_acquire_bits_a_type = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_2_acquire_bits_union = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_union;
  assign outer_arb_io_in_2_acquire_bits_data = BroadcastAcquireTracker_28_1053_io_outer_acquire_bits_data;
  assign outer_arb_io_in_2_grant_ready = BroadcastAcquireTracker_28_1053_io_outer_grant_ready;
  assign outer_arb_io_in_3_acquire_valid = BroadcastAcquireTracker_29_1054_io_outer_acquire_valid;
  assign outer_arb_io_in_3_acquire_bits_addr_block = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_3_acquire_bits_client_xact_id = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_3_acquire_bits_addr_beat = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_3_acquire_bits_is_builtin_type = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_3_acquire_bits_a_type = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_3_acquire_bits_union = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_union;
  assign outer_arb_io_in_3_acquire_bits_data = BroadcastAcquireTracker_29_1054_io_outer_acquire_bits_data;
  assign outer_arb_io_in_3_grant_ready = BroadcastAcquireTracker_29_1054_io_outer_grant_ready;
  assign outer_arb_io_in_4_acquire_valid = BroadcastAcquireTracker_30_1055_io_outer_acquire_valid;
  assign outer_arb_io_in_4_acquire_bits_addr_block = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_block;
  assign outer_arb_io_in_4_acquire_bits_client_xact_id = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_client_xact_id;
  assign outer_arb_io_in_4_acquire_bits_addr_beat = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_addr_beat;
  assign outer_arb_io_in_4_acquire_bits_is_builtin_type = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_is_builtin_type;
  assign outer_arb_io_in_4_acquire_bits_a_type = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_a_type;
  assign outer_arb_io_in_4_acquire_bits_union = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_union;
  assign outer_arb_io_in_4_acquire_bits_data = BroadcastAcquireTracker_30_1055_io_outer_acquire_bits_data;
  assign outer_arb_io_in_4_grant_ready = BroadcastAcquireTracker_30_1055_io_outer_grant_ready;
  assign outer_arb_io_out_acquire_ready = io_outer_acquire_ready;
  assign outer_arb_io_out_grant_valid = io_outer_grant_valid;
  assign outer_arb_io_out_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign outer_arb_io_out_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign outer_arb_io_out_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign outer_arb_io_out_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign outer_arb_io_out_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign outer_arb_io_out_grant_bits_data = io_outer_grant_bits_data[4:0];
  assign outer_data_ptr_idx = T_2482;
  assign outer_data_ptr_loc = T_2481;
  assign T_2481 = outer_arb_io_out_acquire_bits_data[1:0];
  assign T_2482 = outer_arb_io_out_acquire_bits_data[4:2];
  assign is_in_sdq = outer_data_ptr_loc == 2'h0;
  assign T_2483 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_2492_0 = 3'h2;
  assign T_2492_1 = 3'h3;
  assign T_2492_2 = 3'h4;
  assign T_2494 = T_2492_0 == io_outer_acquire_bits_a_type;
  assign T_2495 = T_2492_1 == io_outer_acquire_bits_a_type;
  assign T_2496 = T_2492_2 == io_outer_acquire_bits_a_type;
  assign T_2499 = T_2494 | T_2495;
  assign T_2500 = T_2499 | T_2496;
  assign T_2501 = io_outer_acquire_bits_is_builtin_type & T_2500;
  assign T_2502 = T_2483 & T_2501;
  assign free_sdq = T_2502 & is_in_sdq;
  assign T_2504 = 2'h1 == outer_data_ptr_loc;
  assign GEN_3 = GEN_50;
  assign GEN_44 = GEN_61 == outer_data_ptr_idx ? vwbdq_1 : vwbdq_0;
  assign GEN_45 = GEN_62 == outer_data_ptr_idx ? vwbdq_2 : GEN_44;
  assign GEN_46 = GEN_63 == outer_data_ptr_idx ? vwbdq_3 : GEN_45;
  assign GEN_47 = 3'h4 == outer_data_ptr_idx ? vwbdq_4 : GEN_46;
  assign GEN_48 = 3'h5 == outer_data_ptr_idx ? vwbdq_5 : GEN_47;
  assign GEN_49 = 3'h6 == outer_data_ptr_idx ? vwbdq_6 : GEN_48;
  assign GEN_50 = 3'h7 == outer_data_ptr_idx ? vwbdq_7 : GEN_49;
  assign T_2505 = T_2504 ? GEN_3 : io_inner_release_bits_data;
  assign T_2506 = 2'h0 == outer_data_ptr_loc;
  assign GEN_4 = GEN_57;
  assign GEN_51 = GEN_61 == outer_data_ptr_idx ? sdq_1 : sdq_0;
  assign GEN_52 = GEN_62 == outer_data_ptr_idx ? sdq_2 : GEN_51;
  assign GEN_53 = GEN_63 == outer_data_ptr_idx ? sdq_3 : GEN_52;
  assign GEN_54 = 3'h4 == outer_data_ptr_idx ? sdq_4 : GEN_53;
  assign GEN_55 = 3'h5 == outer_data_ptr_idx ? sdq_5 : GEN_54;
  assign GEN_56 = 3'h6 == outer_data_ptr_idx ? sdq_6 : GEN_55;
  assign GEN_57 = 3'h7 == outer_data_ptr_idx ? sdq_7 : GEN_56;
  assign T_2507 = T_2506 ? GEN_4 : T_2505;
  assign T_2508 = io_outer_acquire_valid | sdq_enq;
  assign GEN_88 = {{7'd0}, 1'h1};
  assign T_2510 = GEN_88 << outer_data_ptr_idx;
  assign GEN_89 = {{7'd0}, free_sdq};
  assign T_2512 = 8'h0 - GEN_89;
  assign T_2513 = T_2512[7:0];
  assign T_2514 = T_2510 & T_2513;
  assign T_2515 = ~ T_2514;
  assign T_2516 = sdq_val & T_2515;
  assign T_2537 = T_1071 ? 8'h80 : 8'h0;
  assign T_2538 = T_1070 ? 8'h40 : T_2537;
  assign T_2539 = T_1069 ? 8'h20 : T_2538;
  assign T_2540 = T_1068 ? 8'h10 : T_2539;
  assign T_2541 = T_1067 ? 8'h8 : T_2540;
  assign T_2542 = T_1066 ? 8'h4 : T_2541;
  assign T_2543 = T_1065 ? 8'h2 : T_2542;
  assign T_2544 = T_1064 ? 8'h1 : T_2543;
  assign GEN_90 = {{7'd0}, sdq_enq};
  assign T_2546 = 8'h0 - GEN_90;
  assign T_2547 = T_2546[7:0];
  assign T_2548 = T_2544 & T_2547;
  assign T_2549 = T_2516 | T_2548;
  assign GEN_58 = T_2508 ? T_2549 : sdq_val;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_68 = {2{$random}};
  sdq_0 = GEN_68[63:0];
  GEN_69 = {2{$random}};
  sdq_1 = GEN_69[63:0];
  GEN_70 = {2{$random}};
  sdq_2 = GEN_70[63:0];
  GEN_71 = {2{$random}};
  sdq_3 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  sdq_4 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  sdq_5 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  sdq_6 = GEN_74[63:0];
  GEN_75 = {2{$random}};
  sdq_7 = GEN_75[63:0];
  GEN_76 = {1{$random}};
  sdq_val = GEN_76[7:0];
  GEN_77 = {1{$random}};
  rel_data_cnt = GEN_77[2:0];
  GEN_78 = {2{$random}};
  vwbdq_0 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  vwbdq_1 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  vwbdq_2 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  vwbdq_3 = GEN_81[63:0];
  GEN_82 = {2{$random}};
  vwbdq_4 = GEN_82[63:0];
  GEN_83 = {2{$random}};
  vwbdq_5 = GEN_83[63:0];
  GEN_84 = {2{$random}};
  vwbdq_6 = GEN_84[63:0];
  GEN_85 = {2{$random}};
  vwbdq_7 = GEN_85[63:0];
  GEN_86 = {1{$random}};
  GEN_13 = GEN_86[0:0];
  GEN_87 = {1{$random}};
  GEN_31 = GEN_87[0:0];
  GEN_91 = {1{$random}};
  GEN_65 = GEN_91[0:0];
  GEN_92 = {1{$random}};
  GEN_66 = GEN_92[0:0];
  GEN_93 = {1{$random}};
  GEN_67 = GEN_93[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      sdq_0 <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      sdq_1 <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      sdq_2 <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      sdq_3 <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      sdq_4 <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      sdq_5 <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      sdq_6 <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      sdq_7 <= GEN_21;
    end
    if(reset) begin
      sdq_val <= 8'h0;
    end else begin
      sdq_val <= GEN_58;
    end
    if(reset) begin
      rel_data_cnt <= 3'h0;
    end else begin
      rel_data_cnt <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      vwbdq_0 <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      vwbdq_1 <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      vwbdq_2 <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      vwbdq_3 <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      vwbdq_4 <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      vwbdq_5 <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      vwbdq_6 <= GEN_38;
    end
    if(1'h0) begin
    end else begin
      vwbdq_7 <= GEN_39;
    end
  end
endmodule
module MMIOTileLinkManager(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [1:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input  [1:0] io_inner_acquire_bits_client_id,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [1:0] io_inner_grant_bits_client_xact_id,
  output [2:0] io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output [1:0] io_inner_grant_bits_client_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input  [2:0] io_inner_finish_bits_manager_xact_id,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output [1:0] io_inner_probe_bits_client_id,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [1:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input  [1:0] io_inner_release_bits_client_id,
  input   io_incoherent_0,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [1:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [1:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data
);
  wire  T_952;
  wire [2:0] T_961_0;
  wire  T_963;
  wire  T_966;
  wire  multibeat_fire;
  wire [2:0] GEN_43;
  wire  T_968;
  wire  multibeat_start;
  wire  T_970;
  wire  multibeat_end;
  reg [5:0] xact_pending;
  reg [31:0] GEN_54;
  wire [5:0] T_972;
  wire  T_973;
  wire  T_974;
  wire  T_975;
  wire  T_976;
  wire  T_977;
  wire [2:0] T_985;
  wire [2:0] T_986;
  wire [2:0] T_987;
  wire [2:0] T_988;
  wire [2:0] xact_id_sel;
  reg [2:0] xact_id_reg;
  reg [31:0] GEN_58;
  wire [2:0] GEN_4;
  reg  xact_multibeat;
  reg [31:0] GEN_59;
  wire [2:0] outer_xact_id;
  wire [5:0] GEN_44;
  wire  T_992;
  wire  xact_free;
  reg [1:0] xact_buffer_0_client_id;
  reg [31:0] GEN_60;
  reg [1:0] xact_buffer_0_client_xact_id;
  reg [31:0] GEN_61;
  reg [1:0] xact_buffer_1_client_id;
  reg [31:0] GEN_64;
  reg [1:0] xact_buffer_1_client_xact_id;
  reg [31:0] GEN_65;
  reg [1:0] xact_buffer_2_client_id;
  reg [31:0] GEN_66;
  reg [1:0] xact_buffer_2_client_xact_id;
  reg [31:0] GEN_67;
  reg [1:0] xact_buffer_3_client_id;
  reg [31:0] GEN_68;
  reg [1:0] xact_buffer_3_client_xact_id;
  reg [31:0] GEN_69;
  reg [1:0] xact_buffer_4_client_id;
  reg [31:0] GEN_70;
  reg [1:0] xact_buffer_4_client_xact_id;
  reg [31:0] GEN_71;
  reg [1:0] xact_buffer_5_client_id;
  reg [31:0] GEN_72;
  reg [1:0] xact_buffer_5_client_xact_id;
  reg [31:0] GEN_73;
  wire  T_1451;
  wire  T_1452;
  wire [2:0] T_1462_0;
  wire  T_1464;
  wire  T_1467;
  wire  T_1469;
  wire  T_1472;
  wire  T_1473;
  wire [3:0] GEN_45;
  wire [3:0] T_1475;
  wire [3:0] T_1477;
  wire [5:0] GEN_46;
  wire [5:0] T_1478;
  wire  T_1479;
  wire [7:0] GEN_47;
  wire [7:0] T_1481;
  wire [7:0] T_1483;
  wire [7:0] T_1484;
  wire [7:0] GEN_48;
  wire [7:0] T_1485;
  wire  T_1486;
  wire [2:0] T_1494_0;
  wire [3:0] GEN_49;
  wire  T_1496;
  wire [1:0] T_1504_0;
  wire [1:0] T_1504_1;
  wire [3:0] GEN_50;
  wire  T_1506;
  wire [3:0] GEN_51;
  wire  T_1507;
  wire  T_1510;
  wire  T_1511;
  wire  T_1514;
  wire  T_1516;
  wire  T_1517;
  wire  T_1518;
  wire [3:0] GEN_52;
  wire  T_1523;
  wire  T_1524;
  wire  T_1526;
  wire  T_1529;
  wire  T_1530;
  wire [7:0] T_1532;
  wire [7:0] T_1534;
  wire [7:0] T_1535;
  wire [7:0] T_1536;
  wire [2:0] T_1546_0;
  wire  T_1548;
  wire  T_1551;
  wire  T_1553;
  wire  T_1556;
  wire  T_1557;
  wire [1:0] GEN_0;
  wire [1:0] GEN_5;
  wire [2:0] GEN_55;
  wire [1:0] GEN_6;
  wire [2:0] GEN_56;
  wire [1:0] GEN_7;
  wire [2:0] GEN_57;
  wire [1:0] GEN_8;
  wire [1:0] GEN_9;
  wire [1:0] GEN_10;
  wire [1:0] GEN_1;
  wire [1:0] GEN_11;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [1:0] GEN_14;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_18;
  wire [1:0] GEN_19;
  wire [1:0] GEN_20;
  wire [1:0] GEN_21;
  wire [1:0] GEN_22;
  wire [1:0] GEN_23;
  wire [1:0] GEN_25;
  wire [1:0] GEN_26;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [1:0] GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire [1:0] GEN_2;
  wire [1:0] GEN_62;
  wire [1:0] GEN_33;
  wire [1:0] GEN_34;
  wire [1:0] GEN_35;
  wire [2:0] GEN_63;
  wire [1:0] GEN_36;
  wire [1:0] GEN_37;
  wire [1:0] GEN_3;
  wire [1:0] GEN_38;
  wire [1:0] GEN_39;
  wire [1:0] GEN_40;
  wire [1:0] GEN_41;
  wire [1:0] GEN_42;
  reg [25:0] GEN_17;
  reg [31:0] GEN_74;
  reg [1:0] GEN_24;
  reg [31:0] GEN_75;
  reg [1:0] GEN_53;
  reg [31:0] GEN_76;
  assign io_inner_acquire_ready = T_1451;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = GEN_3;
  assign io_inner_grant_bits_manager_xact_id = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_client_id = GEN_2;
  assign io_inner_finish_ready = 1'h1;
  assign io_inner_probe_valid = 1'h0;
  assign io_inner_probe_bits_addr_block = GEN_17;
  assign io_inner_probe_bits_p_type = GEN_24;
  assign io_inner_probe_bits_client_id = GEN_53;
  assign io_inner_release_ready = 1'h0;
  assign io_outer_acquire_valid = T_1452;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = outer_xact_id[1:0];
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign T_952 = io_outer_acquire_ready & io_outer_acquire_valid;
  assign T_961_0 = 3'h3;
  assign T_963 = T_961_0 == io_outer_acquire_bits_a_type;
  assign T_966 = io_outer_acquire_bits_is_builtin_type & T_963;
  assign multibeat_fire = T_952 & T_966;
  assign GEN_43 = {{2'd0}, 1'h0};
  assign T_968 = io_outer_acquire_bits_addr_beat == GEN_43;
  assign multibeat_start = multibeat_fire & T_968;
  assign T_970 = io_outer_acquire_bits_addr_beat == 3'h7;
  assign multibeat_end = multibeat_fire & T_970;
  assign T_972 = ~ xact_pending;
  assign T_973 = T_972[0];
  assign T_974 = T_972[1];
  assign T_975 = T_972[2];
  assign T_976 = T_972[3];
  assign T_977 = T_972[4];
  assign T_985 = T_977 ? 3'h4 : 3'h5;
  assign T_986 = T_976 ? {{1'd0}, 2'h3} : T_985;
  assign T_987 = T_975 ? {{1'd0}, 2'h2} : T_986;
  assign T_988 = T_974 ? {{2'd0}, 1'h1} : T_987;
  assign xact_id_sel = T_973 ? {{2'd0}, 1'h0} : T_988;
  assign GEN_4 = multibeat_start ? xact_id_sel : xact_id_reg;
  assign outer_xact_id = xact_multibeat ? xact_id_reg : xact_id_sel;
  assign GEN_44 = {{5'd0}, 1'h0};
  assign T_992 = T_972 == GEN_44;
  assign xact_free = T_992 == 1'h0;
  assign T_1451 = io_outer_acquire_ready & xact_free;
  assign T_1452 = io_inner_acquire_valid & xact_free;
  assign T_1462_0 = 3'h3;
  assign T_1464 = T_1462_0 == io_outer_acquire_bits_a_type;
  assign T_1467 = io_outer_acquire_bits_is_builtin_type & T_1464;
  assign T_1469 = T_1467 == 1'h0;
  assign T_1472 = T_1469 | T_970;
  assign T_1473 = T_952 & T_1472;
  assign GEN_45 = {{3'd0}, 1'h1};
  assign T_1475 = GEN_45 << io_outer_acquire_bits_client_xact_id;
  assign T_1477 = T_1473 ? T_1475 : {{3'd0}, 1'h0};
  assign GEN_46 = {{2'd0}, T_1477};
  assign T_1478 = xact_pending | GEN_46;
  assign T_1479 = io_inner_finish_ready & io_inner_finish_valid;
  assign GEN_47 = {{7'd0}, 1'h1};
  assign T_1481 = GEN_47 << io_inner_finish_bits_manager_xact_id;
  assign T_1483 = T_1479 ? T_1481 : {{7'd0}, 1'h0};
  assign T_1484 = ~ T_1483;
  assign GEN_48 = {{2'd0}, T_1478};
  assign T_1485 = GEN_48 & T_1484;
  assign T_1486 = io_inner_grant_ready & io_inner_grant_valid;
  assign T_1494_0 = 3'h5;
  assign GEN_49 = {{1'd0}, T_1494_0};
  assign T_1496 = GEN_49 == io_inner_grant_bits_g_type;
  assign T_1504_0 = 2'h0;
  assign T_1504_1 = 2'h1;
  assign GEN_50 = {{2'd0}, T_1504_0};
  assign T_1506 = GEN_50 == io_inner_grant_bits_g_type;
  assign GEN_51 = {{2'd0}, T_1504_1};
  assign T_1507 = GEN_51 == io_inner_grant_bits_g_type;
  assign T_1510 = T_1506 | T_1507;
  assign T_1511 = io_inner_grant_bits_is_builtin_type ? T_1496 : T_1510;
  assign T_1514 = T_1511 == 1'h0;
  assign T_1516 = io_inner_grant_bits_addr_beat == 3'h7;
  assign T_1517 = T_1514 | T_1516;
  assign T_1518 = T_1486 & T_1517;
  assign GEN_52 = {{1'd0}, 3'h0};
  assign T_1523 = io_inner_grant_bits_g_type == GEN_52;
  assign T_1524 = io_inner_grant_bits_is_builtin_type & T_1523;
  assign T_1526 = T_1524 == 1'h0;
  assign T_1529 = T_1526 == 1'h0;
  assign T_1530 = T_1518 & T_1529;
  assign T_1532 = GEN_47 << io_inner_grant_bits_manager_xact_id;
  assign T_1534 = T_1530 ? T_1532 : {{7'd0}, 1'h0};
  assign T_1535 = ~ T_1534;
  assign T_1536 = T_1485 & T_1535;
  assign T_1546_0 = 3'h3;
  assign T_1548 = T_1546_0 == io_outer_acquire_bits_a_type;
  assign T_1551 = io_outer_acquire_bits_is_builtin_type & T_1548;
  assign T_1553 = T_1551 == 1'h0;
  assign T_1556 = T_1553 | T_970;
  assign T_1557 = T_952 & T_1556;
  assign GEN_0 = io_inner_acquire_bits_client_id;
  assign GEN_5 = GEN_43 == outer_xact_id ? GEN_0 : xact_buffer_0_client_id;
  assign GEN_55 = {{2'd0}, 1'h1};
  assign GEN_6 = GEN_55 == outer_xact_id ? GEN_0 : xact_buffer_1_client_id;
  assign GEN_56 = {{1'd0}, 2'h2};
  assign GEN_7 = GEN_56 == outer_xact_id ? GEN_0 : xact_buffer_2_client_id;
  assign GEN_57 = {{1'd0}, 2'h3};
  assign GEN_8 = GEN_57 == outer_xact_id ? GEN_0 : xact_buffer_3_client_id;
  assign GEN_9 = 3'h4 == outer_xact_id ? GEN_0 : xact_buffer_4_client_id;
  assign GEN_10 = 3'h5 == outer_xact_id ? GEN_0 : xact_buffer_5_client_id;
  assign GEN_1 = io_inner_acquire_bits_client_xact_id;
  assign GEN_11 = GEN_43 == outer_xact_id ? GEN_1 : xact_buffer_0_client_xact_id;
  assign GEN_12 = GEN_55 == outer_xact_id ? GEN_1 : xact_buffer_1_client_xact_id;
  assign GEN_13 = GEN_56 == outer_xact_id ? GEN_1 : xact_buffer_2_client_xact_id;
  assign GEN_14 = GEN_57 == outer_xact_id ? GEN_1 : xact_buffer_3_client_xact_id;
  assign GEN_15 = 3'h4 == outer_xact_id ? GEN_1 : xact_buffer_4_client_xact_id;
  assign GEN_16 = 3'h5 == outer_xact_id ? GEN_1 : xact_buffer_5_client_xact_id;
  assign GEN_18 = T_1557 ? GEN_5 : xact_buffer_0_client_id;
  assign GEN_19 = T_1557 ? GEN_6 : xact_buffer_1_client_id;
  assign GEN_20 = T_1557 ? GEN_7 : xact_buffer_2_client_id;
  assign GEN_21 = T_1557 ? GEN_8 : xact_buffer_3_client_id;
  assign GEN_22 = T_1557 ? GEN_9 : xact_buffer_4_client_id;
  assign GEN_23 = T_1557 ? GEN_10 : xact_buffer_5_client_id;
  assign GEN_25 = T_1557 ? GEN_11 : xact_buffer_0_client_xact_id;
  assign GEN_26 = T_1557 ? GEN_12 : xact_buffer_1_client_xact_id;
  assign GEN_27 = T_1557 ? GEN_13 : xact_buffer_2_client_xact_id;
  assign GEN_28 = T_1557 ? GEN_14 : xact_buffer_3_client_xact_id;
  assign GEN_29 = T_1557 ? GEN_15 : xact_buffer_4_client_xact_id;
  assign GEN_30 = T_1557 ? GEN_16 : xact_buffer_5_client_xact_id;
  assign GEN_31 = multibeat_start ? 1'h1 : xact_multibeat;
  assign GEN_32 = multibeat_end ? 1'h0 : GEN_31;
  assign GEN_2 = GEN_37;
  assign GEN_62 = {{1'd0}, 1'h1};
  assign GEN_33 = GEN_62 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_id : xact_buffer_0_client_id;
  assign GEN_34 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_id : GEN_33;
  assign GEN_35 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_id : GEN_34;
  assign GEN_63 = {{1'd0}, io_outer_grant_bits_client_xact_id};
  assign GEN_36 = 3'h4 == GEN_63 ? xact_buffer_4_client_id : GEN_35;
  assign GEN_37 = 3'h5 == GEN_63 ? xact_buffer_5_client_id : GEN_36;
  assign GEN_3 = GEN_42;
  assign GEN_38 = GEN_62 == io_outer_grant_bits_client_xact_id ? xact_buffer_1_client_xact_id : xact_buffer_0_client_xact_id;
  assign GEN_39 = 2'h2 == io_outer_grant_bits_client_xact_id ? xact_buffer_2_client_xact_id : GEN_38;
  assign GEN_40 = 2'h3 == io_outer_grant_bits_client_xact_id ? xact_buffer_3_client_xact_id : GEN_39;
  assign GEN_41 = 3'h4 == GEN_63 ? xact_buffer_4_client_xact_id : GEN_40;
  assign GEN_42 = 3'h5 == GEN_63 ? xact_buffer_5_client_xact_id : GEN_41;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_54 = {1{$random}};
  xact_pending = GEN_54[5:0];
  GEN_58 = {1{$random}};
  xact_id_reg = GEN_58[2:0];
  GEN_59 = {1{$random}};
  xact_multibeat = GEN_59[0:0];
  GEN_60 = {1{$random}};
  xact_buffer_0_client_id = GEN_60[1:0];
  GEN_61 = {1{$random}};
  xact_buffer_0_client_xact_id = GEN_61[1:0];
  GEN_64 = {1{$random}};
  xact_buffer_1_client_id = GEN_64[1:0];
  GEN_65 = {1{$random}};
  xact_buffer_1_client_xact_id = GEN_65[1:0];
  GEN_66 = {1{$random}};
  xact_buffer_2_client_id = GEN_66[1:0];
  GEN_67 = {1{$random}};
  xact_buffer_2_client_xact_id = GEN_67[1:0];
  GEN_68 = {1{$random}};
  xact_buffer_3_client_id = GEN_68[1:0];
  GEN_69 = {1{$random}};
  xact_buffer_3_client_xact_id = GEN_69[1:0];
  GEN_70 = {1{$random}};
  xact_buffer_4_client_id = GEN_70[1:0];
  GEN_71 = {1{$random}};
  xact_buffer_4_client_xact_id = GEN_71[1:0];
  GEN_72 = {1{$random}};
  xact_buffer_5_client_id = GEN_72[1:0];
  GEN_73 = {1{$random}};
  xact_buffer_5_client_xact_id = GEN_73[1:0];
  GEN_74 = {1{$random}};
  GEN_17 = GEN_74[25:0];
  GEN_75 = {1{$random}};
  GEN_24 = GEN_75[1:0];
  GEN_76 = {1{$random}};
  GEN_53 = GEN_76[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      xact_pending <= 6'h0;
    end else begin
      xact_pending <= T_1536[5:0];
    end
    if(1'h0) begin
    end else begin
      xact_id_reg <= GEN_4;
    end
    if(reset) begin
      xact_multibeat <= 1'h0;
    end else begin
      xact_multibeat <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_0_client_id <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_0_client_xact_id <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_1_client_id <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_1_client_xact_id <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_2_client_id <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_2_client_xact_id <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_3_client_id <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_3_client_xact_id <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_4_client_id <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_4_client_xact_id <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_5_client_id <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      xact_buffer_5_client_xact_id <= GEN_30;
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_34(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module TileLinkMemoryInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [2:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [2:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [2:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [2:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data
);
  wire  ClientUncachedTileLinkIOArbiter_34_3008_clk;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_reset;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_ready;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_block;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_data;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_ready;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_valid;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_addr_beat;
  wire [2:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_data;
  wire [25:0] T_3010;
  ClientUncachedTileLinkIOArbiter_34 ClientUncachedTileLinkIOArbiter_34_3008 (
    .clk(ClientUncachedTileLinkIOArbiter_34_3008_clk),
    .reset(ClientUncachedTileLinkIOArbiter_34_3008_reset),
    .io_in_0_acquire_ready(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_ready),
    .io_in_0_grant_valid(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_data),
    .io_out_acquire_ready(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_ready),
    .io_out_acquire_valid(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_ready),
    .io_out_grant_valid(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = T_3010;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_34_3008_clk = clk;
  assign ClientUncachedTileLinkIOArbiter_34_3008_reset = reset;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_in_0_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIOArbiter_34_3008_io_out_grant_bits_data = io_out_0_grant_bits_data;
  assign T_3010 = ClientUncachedTileLinkIOArbiter_34_3008_io_out_acquire_bits_addr_block >> 1'h0;
endmodule
module LockingRRArbiter_35(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [2:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [2:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [2:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_8;
  wire [25:0] GEN_1;
  wire [25:0] GEN_9;
  wire [2:0] GEN_2;
  wire [2:0] GEN_10;
  wire [2:0] GEN_3;
  wire [2:0] GEN_11;
  wire  GEN_4;
  wire  GEN_12;
  wire [2:0] GEN_5;
  wire [2:0] GEN_13;
  wire [11:0] GEN_6;
  wire [11:0] GEN_14;
  wire [63:0] GEN_7;
  wire [63:0] GEN_15;
  reg [2:0] T_766;
  reg [31:0] GEN_24;
  reg  T_768;
  reg [31:0] GEN_25;
  wire [2:0] GEN_22;
  wire  T_770;
  wire [2:0] T_779_0;
  wire  T_781;
  wire  T_784;
  wire  T_785;
  wire  T_786;
  wire [2:0] GEN_23;
  wire [3:0] T_790;
  wire [2:0] T_791;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire  GEN_18;
  reg  lastGrant;
  reg [31:0] GEN_26;
  wire  GEN_19;
  wire  T_796;
  wire  T_798;
  wire  T_801;
  wire  T_805;
  wire  T_807;
  wire  T_811;
  wire  T_813;
  wire  T_814;
  wire  T_815;
  wire  T_818;
  wire  T_819;
  wire  GEN_20;
  wire  GEN_21;
  assign io_in_0_ready = T_815;
  assign io_in_1_ready = T_819;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_18;
  assign choice = GEN_21;
  assign GEN_0 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_2 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_4 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_6 = GEN_14;
  assign GEN_14 = io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_7 = GEN_15;
  assign GEN_15 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_22 = {{2'd0}, 1'h0};
  assign T_770 = T_766 != GEN_22;
  assign T_779_0 = 3'h3;
  assign T_781 = T_779_0 == io_out_bits_a_type;
  assign T_784 = io_out_bits_is_builtin_type & T_781;
  assign T_785 = io_out_ready & io_out_valid;
  assign T_786 = T_785 & T_784;
  assign GEN_23 = {{2'd0}, 1'h1};
  assign T_790 = T_766 + GEN_23;
  assign T_791 = T_790[2:0];
  assign GEN_16 = T_786 ? io_chosen : T_768;
  assign GEN_17 = T_786 ? T_791 : T_766;
  assign GEN_18 = T_770 ? T_768 : choice;
  assign GEN_19 = T_785 ? io_chosen : lastGrant;
  assign T_796 = 1'h1 > lastGrant;
  assign T_798 = io_in_1_valid & T_796;
  assign T_801 = T_798 | io_in_0_valid;
  assign T_805 = T_798 == 1'h0;
  assign T_807 = T_801 == 1'h0;
  assign T_811 = T_796 | T_807;
  assign T_813 = T_768 == 1'h0;
  assign T_814 = T_770 ? T_813 : T_805;
  assign T_815 = T_814 & io_out_ready;
  assign T_818 = T_770 ? T_768 : T_811;
  assign T_819 = T_818 & io_out_ready;
  assign GEN_20 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_21 = T_798 ? 1'h1 : GEN_20;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_24 = {1{$random}};
  T_766 = GEN_24[2:0];
  GEN_25 = {1{$random}};
  T_768 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  lastGrant = GEN_26[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_766 <= 3'h0;
    end else begin
      T_766 <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      T_768 <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_19;
    end
  end
endmodule
module ReorderQueue(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits_data,
  input  [2:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [2:0] io_deq_tag,
  output  io_deq_data,
  output  io_deq_matches
);
  reg  roq_data [0:5];
  reg [31:0] GEN_15;
  wire  roq_data_T_104_data;
  wire [2:0] roq_data_T_104_addr;
  wire  roq_data_T_104_en;
  wire  roq_data_T_111_data;
  wire [2:0] roq_data_T_111_addr;
  wire  roq_data_T_111_mask;
  wire  roq_data_T_111_en;
  reg [2:0] roq_tags_0;
  reg [31:0] GEN_16;
  reg [2:0] roq_tags_1;
  reg [31:0] GEN_17;
  reg [2:0] roq_tags_2;
  reg [31:0] GEN_18;
  reg [2:0] roq_tags_3;
  reg [31:0] GEN_19;
  reg [2:0] roq_tags_4;
  reg [31:0] GEN_20;
  reg [2:0] roq_tags_5;
  reg [31:0] GEN_27;
  wire  T_50_0;
  wire  T_50_1;
  wire  T_50_2;
  wire  T_50_3;
  wire  T_50_4;
  wire  T_50_5;
  reg  roq_free_0;
  reg [31:0] GEN_40;
  reg  roq_free_1;
  reg [31:0] GEN_51;
  reg  roq_free_2;
  reg [31:0] GEN_52;
  reg  roq_free_3;
  reg [31:0] GEN_53;
  reg  roq_free_4;
  reg [31:0] GEN_54;
  reg  roq_free_5;
  reg [31:0] GEN_55;
  wire [2:0] T_61;
  wire [2:0] T_62;
  wire [2:0] T_63;
  wire [2:0] T_64;
  wire [2:0] roq_enq_addr;
  wire  T_65;
  wire  T_67;
  wire  T_68;
  wire  T_69;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire  T_75;
  wire  T_76;
  wire  T_77;
  wire  T_79;
  wire  T_80;
  wire  T_81;
  wire  T_83;
  wire  T_84;
  wire  T_85;
  wire  T_87;
  wire  T_88;
  wire [2:0] T_95;
  wire [2:0] T_96;
  wire [2:0] T_97;
  wire [2:0] T_98;
  wire [2:0] roq_deq_addr;
  wire  T_99;
  wire  T_100;
  wire  T_101;
  wire  T_102;
  wire  T_103;
  wire  T_105;
  wire  T_106;
  wire  T_107;
  wire  T_108;
  wire  T_109;
  wire  T_110;
  wire [2:0] GEN_0;
  wire [2:0] GEN_47;
  wire [2:0] GEN_3;
  wire [2:0] GEN_48;
  wire [2:0] GEN_4;
  wire [2:0] GEN_49;
  wire [2:0] GEN_5;
  wire [2:0] GEN_50;
  wire [2:0] GEN_6;
  wire [2:0] GEN_7;
  wire [2:0] GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [2:0] GEN_21;
  wire [2:0] GEN_22;
  wire [2:0] GEN_23;
  wire [2:0] GEN_24;
  wire [2:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_2;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  assign io_enq_ready = T_103;
  assign io_deq_data = roq_data_T_104_data;
  assign io_deq_matches = T_109;
  assign roq_data_T_104_addr = roq_deq_addr;
  assign roq_data_T_104_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_T_104_data = roq_data[roq_data_T_104_addr];
  `else
  assign roq_data_T_104_data = roq_data_T_104_addr >= 3'h6 ? $random : roq_data[roq_data_T_104_addr];
  `endif
  assign roq_data_T_111_data = io_enq_bits_data;
  assign roq_data_T_111_addr = roq_enq_addr;
  assign roq_data_T_111_mask = T_110;
  assign roq_data_T_111_en = T_110;
  assign T_50_0 = 1'h1;
  assign T_50_1 = 1'h1;
  assign T_50_2 = 1'h1;
  assign T_50_3 = 1'h1;
  assign T_50_4 = 1'h1;
  assign T_50_5 = 1'h1;
  assign T_61 = roq_free_4 ? 3'h4 : 3'h5;
  assign T_62 = roq_free_3 ? {{1'd0}, 2'h3} : T_61;
  assign T_63 = roq_free_2 ? {{1'd0}, 2'h2} : T_62;
  assign T_64 = roq_free_1 ? {{2'd0}, 1'h1} : T_63;
  assign roq_enq_addr = roq_free_0 ? {{2'd0}, 1'h0} : T_64;
  assign T_65 = roq_tags_0 == io_deq_tag;
  assign T_67 = roq_free_0 == 1'h0;
  assign T_68 = T_65 & T_67;
  assign T_69 = roq_tags_1 == io_deq_tag;
  assign T_71 = roq_free_1 == 1'h0;
  assign T_72 = T_69 & T_71;
  assign T_73 = roq_tags_2 == io_deq_tag;
  assign T_75 = roq_free_2 == 1'h0;
  assign T_76 = T_73 & T_75;
  assign T_77 = roq_tags_3 == io_deq_tag;
  assign T_79 = roq_free_3 == 1'h0;
  assign T_80 = T_77 & T_79;
  assign T_81 = roq_tags_4 == io_deq_tag;
  assign T_83 = roq_free_4 == 1'h0;
  assign T_84 = T_81 & T_83;
  assign T_85 = roq_tags_5 == io_deq_tag;
  assign T_87 = roq_free_5 == 1'h0;
  assign T_88 = T_85 & T_87;
  assign T_95 = T_84 ? 3'h4 : 3'h5;
  assign T_96 = T_80 ? {{1'd0}, 2'h3} : T_95;
  assign T_97 = T_76 ? {{1'd0}, 2'h2} : T_96;
  assign T_98 = T_72 ? {{2'd0}, 1'h1} : T_97;
  assign roq_deq_addr = T_68 ? {{2'd0}, 1'h0} : T_98;
  assign T_99 = roq_free_0 | roq_free_1;
  assign T_100 = T_99 | roq_free_2;
  assign T_101 = T_100 | roq_free_3;
  assign T_102 = T_101 | roq_free_4;
  assign T_103 = T_102 | roq_free_5;
  assign T_105 = T_68 | T_72;
  assign T_106 = T_105 | T_76;
  assign T_107 = T_106 | T_80;
  assign T_108 = T_107 | T_84;
  assign T_109 = T_108 | T_88;
  assign T_110 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_47 = {{2'd0}, 1'h0};
  assign GEN_3 = GEN_47 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_48 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_48 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_49 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_49 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_50 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_50 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_7 = 3'h4 == roq_enq_addr ? GEN_0 : roq_tags_4;
  assign GEN_8 = 3'h5 == roq_enq_addr ? GEN_0 : roq_tags_5;
  assign GEN_1 = 1'h0;
  assign GEN_9 = GEN_47 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_10 = GEN_48 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_11 = GEN_49 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_12 = GEN_50 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_13 = 3'h4 == roq_enq_addr ? GEN_1 : roq_free_4;
  assign GEN_14 = 3'h5 == roq_enq_addr ? GEN_1 : roq_free_5;
  assign GEN_21 = T_110 ? GEN_3 : roq_tags_0;
  assign GEN_22 = T_110 ? GEN_4 : roq_tags_1;
  assign GEN_23 = T_110 ? GEN_5 : roq_tags_2;
  assign GEN_24 = T_110 ? GEN_6 : roq_tags_3;
  assign GEN_25 = T_110 ? GEN_7 : roq_tags_4;
  assign GEN_26 = T_110 ? GEN_8 : roq_tags_5;
  assign GEN_28 = T_110 ? GEN_9 : roq_free_0;
  assign GEN_29 = T_110 ? GEN_10 : roq_free_1;
  assign GEN_30 = T_110 ? GEN_11 : roq_free_2;
  assign GEN_31 = T_110 ? GEN_12 : roq_free_3;
  assign GEN_32 = T_110 ? GEN_13 : roq_free_4;
  assign GEN_33 = T_110 ? GEN_14 : roq_free_5;
  assign GEN_2 = 1'h1;
  assign GEN_34 = GEN_47 == roq_deq_addr ? GEN_2 : GEN_28;
  assign GEN_35 = GEN_48 == roq_deq_addr ? GEN_2 : GEN_29;
  assign GEN_36 = GEN_49 == roq_deq_addr ? GEN_2 : GEN_30;
  assign GEN_37 = GEN_50 == roq_deq_addr ? GEN_2 : GEN_31;
  assign GEN_38 = 3'h4 == roq_deq_addr ? GEN_2 : GEN_32;
  assign GEN_39 = 3'h5 == roq_deq_addr ? GEN_2 : GEN_33;
  assign GEN_41 = io_deq_valid ? GEN_34 : GEN_28;
  assign GEN_42 = io_deq_valid ? GEN_35 : GEN_29;
  assign GEN_43 = io_deq_valid ? GEN_36 : GEN_30;
  assign GEN_44 = io_deq_valid ? GEN_37 : GEN_31;
  assign GEN_45 = io_deq_valid ? GEN_38 : GEN_32;
  assign GEN_46 = io_deq_valid ? GEN_39 : GEN_33;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data[initvar] = GEN_15[0:0];
  GEN_16 = {1{$random}};
  roq_tags_0 = GEN_16[2:0];
  GEN_17 = {1{$random}};
  roq_tags_1 = GEN_17[2:0];
  GEN_18 = {1{$random}};
  roq_tags_2 = GEN_18[2:0];
  GEN_19 = {1{$random}};
  roq_tags_3 = GEN_19[2:0];
  GEN_20 = {1{$random}};
  roq_tags_4 = GEN_20[2:0];
  GEN_27 = {1{$random}};
  roq_tags_5 = GEN_27[2:0];
  GEN_40 = {1{$random}};
  roq_free_0 = GEN_40[0:0];
  GEN_51 = {1{$random}};
  roq_free_1 = GEN_51[0:0];
  GEN_52 = {1{$random}};
  roq_free_2 = GEN_52[0:0];
  GEN_53 = {1{$random}};
  roq_free_3 = GEN_53[0:0];
  GEN_54 = {1{$random}};
  roq_free_4 = GEN_54[0:0];
  GEN_55 = {1{$random}};
  roq_free_5 = GEN_55[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_T_111_en & roq_data_T_111_mask) begin
      roq_data[roq_data_T_111_addr] <= roq_data_T_111_data;
    end
    if(1'h0) begin
    end else begin
      roq_tags_0 <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      roq_tags_1 <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      roq_tags_2 <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      roq_tags_3 <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      roq_tags_4 <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      roq_tags_5 <= GEN_26;
    end
    if(reset) begin
      roq_free_0 <= T_50_0;
    end else begin
      roq_free_0 <= GEN_41;
    end
    if(reset) begin
      roq_free_1 <= T_50_1;
    end else begin
      roq_free_1 <= GEN_42;
    end
    if(reset) begin
      roq_free_2 <= T_50_2;
    end else begin
      roq_free_2 <= GEN_43;
    end
    if(reset) begin
      roq_free_3 <= T_50_3;
    end else begin
      roq_free_3 <= GEN_44;
    end
    if(reset) begin
      roq_free_4 <= T_50_4;
    end else begin
      roq_free_4 <= GEN_45;
    end
    if(reset) begin
      roq_free_5 <= T_50_5;
    end else begin
      roq_free_5 <= GEN_46;
    end
  end
endmodule
module ClientTileLinkIOUnwrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [2:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_probe_ready,
  output  io_in_probe_valid,
  output [25:0] io_in_probe_bits_addr_block,
  output [1:0] io_in_probe_bits_p_type,
  output  io_in_release_ready,
  input   io_in_release_valid,
  input  [2:0] io_in_release_bits_addr_beat,
  input  [25:0] io_in_release_bits_addr_block,
  input  [2:0] io_in_release_bits_client_xact_id,
  input   io_in_release_bits_voluntary,
  input  [2:0] io_in_release_bits_r_type,
  input  [63:0] io_in_release_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [2:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  output  io_in_grant_bits_manager_id,
  output  io_in_finish_ready,
  input   io_in_finish_valid,
  input   io_in_finish_bits_manager_xact_id,
  input   io_in_finish_bits_manager_id,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  wire  acqArb_clk;
  wire  acqArb_reset;
  wire  acqArb_io_in_0_ready;
  wire  acqArb_io_in_0_valid;
  wire [25:0] acqArb_io_in_0_bits_addr_block;
  wire [2:0] acqArb_io_in_0_bits_client_xact_id;
  wire [2:0] acqArb_io_in_0_bits_addr_beat;
  wire  acqArb_io_in_0_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_0_bits_a_type;
  wire [11:0] acqArb_io_in_0_bits_union;
  wire [63:0] acqArb_io_in_0_bits_data;
  wire  acqArb_io_in_1_ready;
  wire  acqArb_io_in_1_valid;
  wire [25:0] acqArb_io_in_1_bits_addr_block;
  wire [2:0] acqArb_io_in_1_bits_client_xact_id;
  wire [2:0] acqArb_io_in_1_bits_addr_beat;
  wire  acqArb_io_in_1_bits_is_builtin_type;
  wire [2:0] acqArb_io_in_1_bits_a_type;
  wire [11:0] acqArb_io_in_1_bits_union;
  wire [63:0] acqArb_io_in_1_bits_data;
  wire  acqArb_io_out_ready;
  wire  acqArb_io_out_valid;
  wire [25:0] acqArb_io_out_bits_addr_block;
  wire [2:0] acqArb_io_out_bits_client_xact_id;
  wire [2:0] acqArb_io_out_bits_addr_beat;
  wire  acqArb_io_out_bits_is_builtin_type;
  wire [2:0] acqArb_io_out_bits_a_type;
  wire [11:0] acqArb_io_out_bits_union;
  wire [63:0] acqArb_io_out_bits_data;
  wire  acqArb_io_chosen;
  wire  acqRoq_clk;
  wire  acqRoq_reset;
  wire  acqRoq_io_enq_ready;
  wire  acqRoq_io_enq_valid;
  wire  acqRoq_io_enq_bits_data;
  wire [2:0] acqRoq_io_enq_bits_tag;
  wire  acqRoq_io_deq_valid;
  wire [2:0] acqRoq_io_deq_tag;
  wire  acqRoq_io_deq_data;
  wire  acqRoq_io_deq_matches;
  wire  relRoq_clk;
  wire  relRoq_reset;
  wire  relRoq_io_enq_ready;
  wire  relRoq_io_enq_valid;
  wire  relRoq_io_enq_bits_data;
  wire [2:0] relRoq_io_enq_bits_tag;
  wire  relRoq_io_deq_valid;
  wire [2:0] relRoq_io_deq_tag;
  wire  relRoq_io_deq_data;
  wire  relRoq_io_deq_matches;
  wire [2:0] T_1366_0;
  wire  T_1368;
  wire  T_1371;
  wire [2:0] GEN_0;
  wire  T_1373;
  wire  acq_roq_enq;
  wire [2:0] T_1381_0;
  wire [2:0] T_1381_1;
  wire [2:0] T_1381_2;
  wire  T_1383;
  wire  T_1384;
  wire  T_1385;
  wire  T_1388;
  wire  T_1389;
  wire  T_1392;
  wire  rel_roq_enq;
  wire  T_1395;
  wire  acq_roq_ready;
  wire  T_1397;
  wire  rel_roq_ready;
  wire  T_1398;
  wire  T_1399;
  wire  T_1400;
  wire [2:0] T_1403;
  wire [11:0] T_1407;
  wire [25:0] T_1436_addr_block;
  wire [2:0] T_1436_client_xact_id;
  wire [2:0] T_1436_addr_beat;
  wire  T_1436_is_builtin_type;
  wire [2:0] T_1436_a_type;
  wire [11:0] T_1436_union;
  wire [63:0] T_1436_data;
  wire  T_1464;
  wire  T_1465;
  wire  T_1466;
  wire  T_1467;
  wire [7:0] GEN_2;
  wire [7:0] T_1489;
  wire [8:0] T_1536;
  wire [11:0] T_1554;
  wire [25:0] T_1589_addr_block;
  wire [2:0] T_1589_client_xact_id;
  wire [2:0] T_1589_addr_beat;
  wire  T_1589_is_builtin_type;
  wire [2:0] T_1589_a_type;
  wire [11:0] T_1589_union;
  wire [63:0] T_1589_data;
  wire  T_1617;
  wire  T_1618;
  wire [2:0] T_1626_0;
  wire [3:0] GEN_3;
  wire  T_1628;
  wire  T_1636_0;
  wire [3:0] GEN_4;
  wire  T_1638;
  wire  T_1641;
  wire  T_1644;
  wire  T_1646;
  wire  T_1647;
  wire [2:0] T_1656_0;
  wire [3:0] GEN_5;
  wire  T_1658;
  wire  T_1666_0;
  wire [3:0] GEN_6;
  wire  T_1668;
  wire  T_1671;
  wire  T_1676;
  wire  T_1677;
  wire [3:0] T_1678;
  wire [2:0] acq_grant_addr_beat;
  wire [2:0] acq_grant_client_xact_id;
  wire  acq_grant_manager_xact_id;
  wire  acq_grant_is_builtin_type;
  wire [3:0] acq_grant_g_type;
  wire [63:0] acq_grant_data;
  wire [3:0] T_1734;
  wire [2:0] rel_grant_addr_beat;
  wire [2:0] rel_grant_client_xact_id;
  wire  rel_grant_manager_xact_id;
  wire  rel_grant_is_builtin_type;
  wire [3:0] rel_grant_g_type;
  wire [63:0] rel_grant_data;
  wire [2:0] T_1788_addr_beat;
  wire [2:0] T_1788_client_xact_id;
  wire  T_1788_manager_xact_id;
  wire  T_1788_is_builtin_type;
  wire [3:0] T_1788_g_type;
  wire [63:0] T_1788_data;
  reg [25:0] GEN_1;
  reg [31:0] GEN_10;
  reg [1:0] GEN_7;
  reg [31:0] GEN_11;
  reg  GEN_8;
  reg [31:0] GEN_12;
  reg  GEN_9;
  reg [31:0] GEN_13;
  LockingRRArbiter_35 acqArb (
    .clk(acqArb_clk),
    .reset(acqArb_reset),
    .io_in_0_ready(acqArb_io_in_0_ready),
    .io_in_0_valid(acqArb_io_in_0_valid),
    .io_in_0_bits_addr_block(acqArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(acqArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(acqArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(acqArb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(acqArb_io_in_0_bits_a_type),
    .io_in_0_bits_union(acqArb_io_in_0_bits_union),
    .io_in_0_bits_data(acqArb_io_in_0_bits_data),
    .io_in_1_ready(acqArb_io_in_1_ready),
    .io_in_1_valid(acqArb_io_in_1_valid),
    .io_in_1_bits_addr_block(acqArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(acqArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(acqArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(acqArb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(acqArb_io_in_1_bits_a_type),
    .io_in_1_bits_union(acqArb_io_in_1_bits_union),
    .io_in_1_bits_data(acqArb_io_in_1_bits_data),
    .io_out_ready(acqArb_io_out_ready),
    .io_out_valid(acqArb_io_out_valid),
    .io_out_bits_addr_block(acqArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(acqArb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(acqArb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(acqArb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(acqArb_io_out_bits_a_type),
    .io_out_bits_union(acqArb_io_out_bits_union),
    .io_out_bits_data(acqArb_io_out_bits_data),
    .io_chosen(acqArb_io_chosen)
  );
  ReorderQueue acqRoq (
    .clk(acqRoq_clk),
    .reset(acqRoq_reset),
    .io_enq_ready(acqRoq_io_enq_ready),
    .io_enq_valid(acqRoq_io_enq_valid),
    .io_enq_bits_data(acqRoq_io_enq_bits_data),
    .io_enq_bits_tag(acqRoq_io_enq_bits_tag),
    .io_deq_valid(acqRoq_io_deq_valid),
    .io_deq_tag(acqRoq_io_deq_tag),
    .io_deq_data(acqRoq_io_deq_data),
    .io_deq_matches(acqRoq_io_deq_matches)
  );
  ReorderQueue relRoq (
    .clk(relRoq_clk),
    .reset(relRoq_reset),
    .io_enq_ready(relRoq_io_enq_ready),
    .io_enq_valid(relRoq_io_enq_valid),
    .io_enq_bits_data(relRoq_io_enq_bits_data),
    .io_enq_bits_tag(relRoq_io_enq_bits_tag),
    .io_deq_valid(relRoq_io_deq_valid),
    .io_deq_tag(relRoq_io_deq_tag),
    .io_deq_data(relRoq_io_deq_data),
    .io_deq_matches(relRoq_io_deq_matches)
  );
  assign io_in_acquire_ready = T_1464;
  assign io_in_probe_valid = 1'h0;
  assign io_in_probe_bits_addr_block = GEN_1;
  assign io_in_probe_bits_p_type = GEN_7;
  assign io_in_release_ready = T_1617;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = T_1788_addr_beat;
  assign io_in_grant_bits_client_xact_id = T_1788_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = T_1788_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = T_1788_is_builtin_type;
  assign io_in_grant_bits_g_type = T_1788_g_type;
  assign io_in_grant_bits_data = T_1788_data;
  assign io_in_grant_bits_manager_id = GEN_8;
  assign io_in_finish_ready = GEN_9;
  assign io_out_acquire_valid = acqArb_io_out_valid;
  assign io_out_acquire_bits_addr_block = acqArb_io_out_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = acqArb_io_out_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = acqArb_io_out_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = acqArb_io_out_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = acqArb_io_out_bits_a_type;
  assign io_out_acquire_bits_union = acqArb_io_out_bits_union;
  assign io_out_acquire_bits_data = acqArb_io_out_bits_data;
  assign io_out_grant_ready = io_in_grant_ready;
  assign acqArb_clk = clk;
  assign acqArb_reset = reset;
  assign acqArb_io_in_0_valid = T_1400;
  assign acqArb_io_in_0_bits_addr_block = T_1436_addr_block;
  assign acqArb_io_in_0_bits_client_xact_id = T_1436_client_xact_id;
  assign acqArb_io_in_0_bits_addr_beat = T_1436_addr_beat;
  assign acqArb_io_in_0_bits_is_builtin_type = T_1436_is_builtin_type;
  assign acqArb_io_in_0_bits_a_type = T_1436_a_type;
  assign acqArb_io_in_0_bits_union = T_1436_union;
  assign acqArb_io_in_0_bits_data = T_1436_data;
  assign acqArb_io_in_1_valid = T_1467;
  assign acqArb_io_in_1_bits_addr_block = T_1589_addr_block;
  assign acqArb_io_in_1_bits_client_xact_id = T_1589_client_xact_id;
  assign acqArb_io_in_1_bits_addr_beat = T_1589_addr_beat;
  assign acqArb_io_in_1_bits_is_builtin_type = T_1589_is_builtin_type;
  assign acqArb_io_in_1_bits_a_type = T_1589_a_type;
  assign acqArb_io_in_1_bits_union = T_1589_union;
  assign acqArb_io_in_1_bits_data = T_1589_data;
  assign acqArb_io_out_ready = io_out_acquire_ready;
  assign acqRoq_clk = clk;
  assign acqRoq_reset = reset;
  assign acqRoq_io_enq_valid = T_1399;
  assign acqRoq_io_enq_bits_data = io_in_acquire_bits_is_builtin_type;
  assign acqRoq_io_enq_bits_tag = io_in_acquire_bits_client_xact_id;
  assign acqRoq_io_deq_valid = T_1647;
  assign acqRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign relRoq_clk = clk;
  assign relRoq_reset = reset;
  assign relRoq_io_enq_valid = T_1466;
  assign relRoq_io_enq_bits_data = io_in_release_bits_voluntary;
  assign relRoq_io_enq_bits_tag = io_in_release_bits_client_xact_id;
  assign relRoq_io_deq_valid = T_1677;
  assign relRoq_io_deq_tag = io_out_grant_bits_client_xact_id;
  assign T_1366_0 = 3'h3;
  assign T_1368 = T_1366_0 == io_in_acquire_bits_a_type;
  assign T_1371 = io_in_acquire_bits_is_builtin_type & T_1368;
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_1373 = io_in_acquire_bits_addr_beat == GEN_0;
  assign acq_roq_enq = T_1371 ? T_1373 : 1'h1;
  assign T_1381_0 = 3'h0;
  assign T_1381_1 = 3'h1;
  assign T_1381_2 = 3'h2;
  assign T_1383 = T_1381_0 == io_in_release_bits_r_type;
  assign T_1384 = T_1381_1 == io_in_release_bits_r_type;
  assign T_1385 = T_1381_2 == io_in_release_bits_r_type;
  assign T_1388 = T_1383 | T_1384;
  assign T_1389 = T_1388 | T_1385;
  assign T_1392 = io_in_release_bits_addr_beat == GEN_0;
  assign rel_roq_enq = T_1389 ? T_1392 : 1'h1;
  assign T_1395 = acq_roq_enq == 1'h0;
  assign acq_roq_ready = T_1395 | acqRoq_io_enq_ready;
  assign T_1397 = rel_roq_enq == 1'h0;
  assign rel_roq_ready = T_1397 | relRoq_io_enq_ready;
  assign T_1398 = io_in_acquire_valid & acqArb_io_in_0_ready;
  assign T_1399 = T_1398 & acq_roq_enq;
  assign T_1400 = io_in_acquire_valid & acq_roq_ready;
  assign T_1403 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_a_type : 3'h1;
  assign T_1407 = io_in_acquire_bits_is_builtin_type ? io_in_acquire_bits_union : {{3'd0}, 9'h1c1};
  assign T_1436_addr_block = io_in_acquire_bits_addr_block;
  assign T_1436_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign T_1436_addr_beat = io_in_acquire_bits_addr_beat;
  assign T_1436_is_builtin_type = 1'h1;
  assign T_1436_a_type = T_1403;
  assign T_1436_union = T_1407;
  assign T_1436_data = io_in_acquire_bits_data;
  assign T_1464 = acq_roq_ready & acqArb_io_in_0_ready;
  assign T_1465 = io_in_release_valid & acqArb_io_in_1_ready;
  assign T_1466 = T_1465 & rel_roq_enq;
  assign T_1467 = io_in_release_valid & rel_roq_ready;
  assign GEN_2 = $signed(8'hff);
  assign T_1489 = $unsigned(GEN_2);
  assign T_1536 = {T_1489,1'h1};
  assign T_1554 = 1'h1 ? {{3'd0}, T_1536} : 12'h0;
  assign T_1589_addr_block = io_in_release_bits_addr_block;
  assign T_1589_client_xact_id = io_in_release_bits_client_xact_id;
  assign T_1589_addr_beat = io_in_release_bits_addr_beat;
  assign T_1589_is_builtin_type = 1'h1;
  assign T_1589_a_type = 3'h3;
  assign T_1589_union = T_1554;
  assign T_1589_data = io_in_release_bits_data;
  assign T_1617 = rel_roq_ready & acqArb_io_in_1_ready;
  assign T_1618 = io_out_grant_ready & io_out_grant_valid;
  assign T_1626_0 = 3'h5;
  assign GEN_3 = {{1'd0}, T_1626_0};
  assign T_1628 = GEN_3 == io_out_grant_bits_g_type;
  assign T_1636_0 = 1'h0;
  assign GEN_4 = {{3'd0}, T_1636_0};
  assign T_1638 = GEN_4 == io_out_grant_bits_g_type;
  assign T_1641 = io_out_grant_bits_is_builtin_type ? T_1628 : T_1638;
  assign T_1644 = io_out_grant_bits_addr_beat == 3'h7;
  assign T_1646 = T_1641 ? T_1644 : 1'h1;
  assign T_1647 = T_1618 & T_1646;
  assign T_1656_0 = 3'h5;
  assign GEN_5 = {{1'd0}, T_1656_0};
  assign T_1658 = GEN_5 == io_out_grant_bits_g_type;
  assign T_1666_0 = 1'h0;
  assign GEN_6 = {{3'd0}, T_1666_0};
  assign T_1668 = GEN_6 == io_out_grant_bits_g_type;
  assign T_1671 = io_out_grant_bits_is_builtin_type ? T_1658 : T_1668;
  assign T_1676 = T_1671 ? T_1644 : 1'h1;
  assign T_1677 = T_1618 & T_1676;
  assign T_1678 = acqRoq_io_deq_data ? io_out_grant_bits_g_type : {{3'd0}, 1'h0};
  assign acq_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign acq_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign acq_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign acq_grant_is_builtin_type = acqRoq_io_deq_data;
  assign acq_grant_g_type = T_1678;
  assign acq_grant_data = io_out_grant_bits_data;
  assign T_1734 = relRoq_io_deq_data ? {{1'd0}, 3'h0} : io_out_grant_bits_g_type;
  assign rel_grant_addr_beat = io_out_grant_bits_addr_beat;
  assign rel_grant_client_xact_id = io_out_grant_bits_client_xact_id;
  assign rel_grant_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign rel_grant_is_builtin_type = 1'h1;
  assign rel_grant_g_type = T_1734;
  assign rel_grant_data = io_out_grant_bits_data;
  assign T_1788_addr_beat = acqRoq_io_deq_matches ? acq_grant_addr_beat : rel_grant_addr_beat;
  assign T_1788_client_xact_id = acqRoq_io_deq_matches ? acq_grant_client_xact_id : rel_grant_client_xact_id;
  assign T_1788_manager_xact_id = acqRoq_io_deq_matches ? acq_grant_manager_xact_id : rel_grant_manager_xact_id;
  assign T_1788_is_builtin_type = acqRoq_io_deq_matches ? acq_grant_is_builtin_type : rel_grant_is_builtin_type;
  assign T_1788_g_type = acqRoq_io_deq_matches ? acq_grant_g_type : rel_grant_g_type;
  assign T_1788_data = acqRoq_io_deq_matches ? acq_grant_data : rel_grant_data;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_10 = {1{$random}};
  GEN_1 = GEN_10[25:0];
  GEN_11 = {1{$random}};
  GEN_7 = GEN_11[1:0];
  GEN_12 = {1{$random}};
  GEN_8 = GEN_12[0:0];
  GEN_13 = {1{$random}};
  GEN_9 = GEN_13[0:0];
  end
`endif
endmodule
module ClientTileLinkIOWrapper(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [2:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [2:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [2:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_probe_ready,
  input   io_out_probe_valid,
  input  [25:0] io_out_probe_bits_addr_block,
  input  [1:0] io_out_probe_bits_p_type,
  input   io_out_release_ready,
  output  io_out_release_valid,
  output [2:0] io_out_release_bits_addr_beat,
  output [25:0] io_out_release_bits_addr_block,
  output [2:0] io_out_release_bits_client_xact_id,
  output  io_out_release_bits_voluntary,
  output [2:0] io_out_release_bits_r_type,
  output [63:0] io_out_release_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [2:0] io_out_grant_bits_client_xact_id,
  input   io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data,
  input   io_out_grant_bits_manager_id,
  input   io_out_finish_ready,
  output  io_out_finish_valid,
  output  io_out_finish_bits_manager_xact_id,
  output  io_out_finish_bits_manager_id
);
  reg [2:0] GEN_0;
  reg [31:0] GEN_9;
  reg [25:0] GEN_1;
  reg [31:0] GEN_10;
  reg [2:0] GEN_2;
  reg [31:0] GEN_11;
  reg  GEN_3;
  reg [31:0] GEN_12;
  reg [2:0] GEN_4;
  reg [31:0] GEN_13;
  reg [63:0] GEN_5;
  reg [63:0] GEN_14;
  reg  GEN_6;
  reg [31:0] GEN_15;
  reg  GEN_7;
  reg [31:0] GEN_16;
  reg  GEN_8;
  reg [31:0] GEN_17;
  assign io_in_acquire_ready = io_out_acquire_ready;
  assign io_in_grant_valid = io_out_grant_valid;
  assign io_in_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_probe_ready = 1'h1;
  assign io_out_release_valid = 1'h0;
  assign io_out_release_bits_addr_beat = GEN_0;
  assign io_out_release_bits_addr_block = GEN_1;
  assign io_out_release_bits_client_xact_id = GEN_2;
  assign io_out_release_bits_voluntary = GEN_3;
  assign io_out_release_bits_r_type = GEN_4;
  assign io_out_release_bits_data = GEN_5;
  assign io_out_grant_ready = io_in_grant_ready;
  assign io_out_finish_valid = GEN_6;
  assign io_out_finish_bits_manager_xact_id = GEN_7;
  assign io_out_finish_bits_manager_id = GEN_8;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  GEN_0 = GEN_9[2:0];
  GEN_10 = {1{$random}};
  GEN_1 = GEN_10[25:0];
  GEN_11 = {1{$random}};
  GEN_2 = GEN_11[2:0];
  GEN_12 = {1{$random}};
  GEN_3 = GEN_12[0:0];
  GEN_13 = {1{$random}};
  GEN_4 = GEN_13[2:0];
  GEN_14 = {2{$random}};
  GEN_5 = GEN_14[63:0];
  GEN_15 = {1{$random}};
  GEN_6 = GEN_15[0:0];
  GEN_16 = {1{$random}};
  GEN_7 = GEN_16[0:0];
  GEN_17 = {1{$random}};
  GEN_8 = GEN_17[0:0];
  end
`endif
endmodule
module ClientTileLinkEnqueuer(
  input   clk,
  input   reset,
  output  io_inner_acquire_ready,
  input   io_inner_acquire_valid,
  input  [25:0] io_inner_acquire_bits_addr_block,
  input  [2:0] io_inner_acquire_bits_client_xact_id,
  input  [2:0] io_inner_acquire_bits_addr_beat,
  input   io_inner_acquire_bits_is_builtin_type,
  input  [2:0] io_inner_acquire_bits_a_type,
  input  [11:0] io_inner_acquire_bits_union,
  input  [63:0] io_inner_acquire_bits_data,
  input   io_inner_probe_ready,
  output  io_inner_probe_valid,
  output [25:0] io_inner_probe_bits_addr_block,
  output [1:0] io_inner_probe_bits_p_type,
  output  io_inner_release_ready,
  input   io_inner_release_valid,
  input  [2:0] io_inner_release_bits_addr_beat,
  input  [25:0] io_inner_release_bits_addr_block,
  input  [2:0] io_inner_release_bits_client_xact_id,
  input   io_inner_release_bits_voluntary,
  input  [2:0] io_inner_release_bits_r_type,
  input  [63:0] io_inner_release_bits_data,
  input   io_inner_grant_ready,
  output  io_inner_grant_valid,
  output [2:0] io_inner_grant_bits_addr_beat,
  output [2:0] io_inner_grant_bits_client_xact_id,
  output  io_inner_grant_bits_manager_xact_id,
  output  io_inner_grant_bits_is_builtin_type,
  output [3:0] io_inner_grant_bits_g_type,
  output [63:0] io_inner_grant_bits_data,
  output  io_inner_grant_bits_manager_id,
  output  io_inner_finish_ready,
  input   io_inner_finish_valid,
  input   io_inner_finish_bits_manager_xact_id,
  input   io_inner_finish_bits_manager_id,
  input   io_outer_acquire_ready,
  output  io_outer_acquire_valid,
  output [25:0] io_outer_acquire_bits_addr_block,
  output [2:0] io_outer_acquire_bits_client_xact_id,
  output [2:0] io_outer_acquire_bits_addr_beat,
  output  io_outer_acquire_bits_is_builtin_type,
  output [2:0] io_outer_acquire_bits_a_type,
  output [11:0] io_outer_acquire_bits_union,
  output [63:0] io_outer_acquire_bits_data,
  output  io_outer_probe_ready,
  input   io_outer_probe_valid,
  input  [25:0] io_outer_probe_bits_addr_block,
  input  [1:0] io_outer_probe_bits_p_type,
  input   io_outer_release_ready,
  output  io_outer_release_valid,
  output [2:0] io_outer_release_bits_addr_beat,
  output [25:0] io_outer_release_bits_addr_block,
  output [2:0] io_outer_release_bits_client_xact_id,
  output  io_outer_release_bits_voluntary,
  output [2:0] io_outer_release_bits_r_type,
  output [63:0] io_outer_release_bits_data,
  output  io_outer_grant_ready,
  input   io_outer_grant_valid,
  input  [2:0] io_outer_grant_bits_addr_beat,
  input  [2:0] io_outer_grant_bits_client_xact_id,
  input   io_outer_grant_bits_manager_xact_id,
  input   io_outer_grant_bits_is_builtin_type,
  input  [3:0] io_outer_grant_bits_g_type,
  input  [63:0] io_outer_grant_bits_data,
  input   io_outer_grant_bits_manager_id,
  input   io_outer_finish_ready,
  output  io_outer_finish_valid,
  output  io_outer_finish_bits_manager_xact_id,
  output  io_outer_finish_bits_manager_id
);
  assign io_inner_acquire_ready = io_outer_acquire_ready;
  assign io_inner_probe_valid = io_outer_probe_valid;
  assign io_inner_probe_bits_addr_block = io_outer_probe_bits_addr_block;
  assign io_inner_probe_bits_p_type = io_outer_probe_bits_p_type;
  assign io_inner_release_ready = io_outer_release_ready;
  assign io_inner_grant_valid = io_outer_grant_valid;
  assign io_inner_grant_bits_addr_beat = io_outer_grant_bits_addr_beat;
  assign io_inner_grant_bits_client_xact_id = io_outer_grant_bits_client_xact_id;
  assign io_inner_grant_bits_manager_xact_id = io_outer_grant_bits_manager_xact_id;
  assign io_inner_grant_bits_is_builtin_type = io_outer_grant_bits_is_builtin_type;
  assign io_inner_grant_bits_g_type = io_outer_grant_bits_g_type;
  assign io_inner_grant_bits_data = io_outer_grant_bits_data;
  assign io_inner_grant_bits_manager_id = io_outer_grant_bits_manager_id;
  assign io_inner_finish_ready = io_outer_finish_ready;
  assign io_outer_acquire_valid = io_inner_acquire_valid;
  assign io_outer_acquire_bits_addr_block = io_inner_acquire_bits_addr_block;
  assign io_outer_acquire_bits_client_xact_id = io_inner_acquire_bits_client_xact_id;
  assign io_outer_acquire_bits_addr_beat = io_inner_acquire_bits_addr_beat;
  assign io_outer_acquire_bits_is_builtin_type = io_inner_acquire_bits_is_builtin_type;
  assign io_outer_acquire_bits_a_type = io_inner_acquire_bits_a_type;
  assign io_outer_acquire_bits_union = io_inner_acquire_bits_union;
  assign io_outer_acquire_bits_data = io_inner_acquire_bits_data;
  assign io_outer_probe_ready = io_inner_probe_ready;
  assign io_outer_release_valid = io_inner_release_valid;
  assign io_outer_release_bits_addr_beat = io_inner_release_bits_addr_beat;
  assign io_outer_release_bits_addr_block = io_inner_release_bits_addr_block;
  assign io_outer_release_bits_client_xact_id = io_inner_release_bits_client_xact_id;
  assign io_outer_release_bits_voluntary = io_inner_release_bits_voluntary;
  assign io_outer_release_bits_r_type = io_inner_release_bits_r_type;
  assign io_outer_release_bits_data = io_inner_release_bits_data;
  assign io_outer_grant_ready = io_inner_grant_ready;
  assign io_outer_finish_valid = io_inner_finish_valid;
  assign io_outer_finish_bits_manager_xact_id = io_inner_finish_bits_manager_xact_id;
  assign io_outer_finish_bits_manager_id = io_inner_finish_bits_manager_id;
endmodule
module ReorderQueue_37(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [4:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [4:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] roq_data_addr_beat [0:5];
  reg [31:0] GEN_15;
  wire [2:0] roq_data_addr_beat_T_324_data;
  wire [2:0] roq_data_addr_beat_T_324_addr;
  wire  roq_data_addr_beat_T_324_en;
  wire [2:0] roq_data_addr_beat_T_353_data;
  wire [2:0] roq_data_addr_beat_T_353_addr;
  wire  roq_data_addr_beat_T_353_mask;
  wire  roq_data_addr_beat_T_353_en;
  reg  roq_data_subblock [0:5];
  reg [31:0] GEN_16;
  wire  roq_data_subblock_T_324_data;
  wire [2:0] roq_data_subblock_T_324_addr;
  wire  roq_data_subblock_T_324_en;
  wire  roq_data_subblock_T_353_data;
  wire [2:0] roq_data_subblock_T_353_addr;
  wire  roq_data_subblock_T_353_mask;
  wire  roq_data_subblock_T_353_en;
  reg [4:0] roq_tags_0;
  reg [31:0] GEN_17;
  reg [4:0] roq_tags_1;
  reg [31:0] GEN_18;
  reg [4:0] roq_tags_2;
  reg [31:0] GEN_19;
  reg [4:0] roq_tags_3;
  reg [31:0] GEN_20;
  reg [4:0] roq_tags_4;
  reg [31:0] GEN_21;
  reg [4:0] roq_tags_5;
  reg [31:0] GEN_22;
  wire  T_270_0;
  wire  T_270_1;
  wire  T_270_2;
  wire  T_270_3;
  wire  T_270_4;
  wire  T_270_5;
  reg  roq_free_0;
  reg [31:0] GEN_29;
  reg  roq_free_1;
  reg [31:0] GEN_42;
  reg  roq_free_2;
  reg [31:0] GEN_53;
  reg  roq_free_3;
  reg [31:0] GEN_54;
  reg  roq_free_4;
  reg [31:0] GEN_55;
  reg  roq_free_5;
  reg [31:0] GEN_56;
  wire [2:0] T_281;
  wire [2:0] T_282;
  wire [2:0] T_283;
  wire [2:0] T_284;
  wire [2:0] roq_enq_addr;
  wire  T_285;
  wire  T_287;
  wire  T_288;
  wire  T_289;
  wire  T_291;
  wire  T_292;
  wire  T_293;
  wire  T_295;
  wire  T_296;
  wire  T_297;
  wire  T_299;
  wire  T_300;
  wire  T_301;
  wire  T_303;
  wire  T_304;
  wire  T_305;
  wire  T_307;
  wire  T_308;
  wire [2:0] T_315;
  wire [2:0] T_316;
  wire [2:0] T_317;
  wire [2:0] T_318;
  wire [2:0] roq_deq_addr;
  wire  T_319;
  wire  T_320;
  wire  T_321;
  wire  T_322;
  wire  T_323;
  wire  T_347;
  wire  T_348;
  wire  T_349;
  wire  T_350;
  wire  T_351;
  wire  T_352;
  wire [4:0] GEN_0;
  wire [2:0] GEN_49;
  wire [4:0] GEN_3;
  wire [2:0] GEN_50;
  wire [4:0] GEN_4;
  wire [2:0] GEN_51;
  wire [4:0] GEN_5;
  wire [2:0] GEN_52;
  wire [4:0] GEN_6;
  wire [4:0] GEN_7;
  wire [4:0] GEN_8;
  wire  GEN_1;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [4:0] GEN_23;
  wire [4:0] GEN_24;
  wire [4:0] GEN_25;
  wire [4:0] GEN_26;
  wire [4:0] GEN_27;
  wire [4:0] GEN_28;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_2;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  assign io_enq_ready = T_323;
  assign io_deq_data_addr_beat = roq_data_addr_beat_T_324_data;
  assign io_deq_data_subblock = roq_data_subblock_T_324_data;
  assign io_deq_matches = T_351;
  assign roq_data_addr_beat_T_324_addr = roq_deq_addr;
  assign roq_data_addr_beat_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_addr_beat_T_324_data = roq_data_addr_beat[roq_data_addr_beat_T_324_addr];
  `else
  assign roq_data_addr_beat_T_324_data = roq_data_addr_beat_T_324_addr >= 3'h6 ? $random : roq_data_addr_beat[roq_data_addr_beat_T_324_addr];
  `endif
  assign roq_data_addr_beat_T_353_data = io_enq_bits_data_addr_beat;
  assign roq_data_addr_beat_T_353_addr = roq_enq_addr;
  assign roq_data_addr_beat_T_353_mask = T_352;
  assign roq_data_addr_beat_T_353_en = T_352;
  assign roq_data_subblock_T_324_addr = roq_deq_addr;
  assign roq_data_subblock_T_324_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_subblock_T_324_data = roq_data_subblock[roq_data_subblock_T_324_addr];
  `else
  assign roq_data_subblock_T_324_data = roq_data_subblock_T_324_addr >= 3'h6 ? $random : roq_data_subblock[roq_data_subblock_T_324_addr];
  `endif
  assign roq_data_subblock_T_353_data = io_enq_bits_data_subblock;
  assign roq_data_subblock_T_353_addr = roq_enq_addr;
  assign roq_data_subblock_T_353_mask = T_352;
  assign roq_data_subblock_T_353_en = T_352;
  assign T_270_0 = 1'h1;
  assign T_270_1 = 1'h1;
  assign T_270_2 = 1'h1;
  assign T_270_3 = 1'h1;
  assign T_270_4 = 1'h1;
  assign T_270_5 = 1'h1;
  assign T_281 = roq_free_4 ? 3'h4 : 3'h5;
  assign T_282 = roq_free_3 ? {{1'd0}, 2'h3} : T_281;
  assign T_283 = roq_free_2 ? {{1'd0}, 2'h2} : T_282;
  assign T_284 = roq_free_1 ? {{2'd0}, 1'h1} : T_283;
  assign roq_enq_addr = roq_free_0 ? {{2'd0}, 1'h0} : T_284;
  assign T_285 = roq_tags_0 == io_deq_tag;
  assign T_287 = roq_free_0 == 1'h0;
  assign T_288 = T_285 & T_287;
  assign T_289 = roq_tags_1 == io_deq_tag;
  assign T_291 = roq_free_1 == 1'h0;
  assign T_292 = T_289 & T_291;
  assign T_293 = roq_tags_2 == io_deq_tag;
  assign T_295 = roq_free_2 == 1'h0;
  assign T_296 = T_293 & T_295;
  assign T_297 = roq_tags_3 == io_deq_tag;
  assign T_299 = roq_free_3 == 1'h0;
  assign T_300 = T_297 & T_299;
  assign T_301 = roq_tags_4 == io_deq_tag;
  assign T_303 = roq_free_4 == 1'h0;
  assign T_304 = T_301 & T_303;
  assign T_305 = roq_tags_5 == io_deq_tag;
  assign T_307 = roq_free_5 == 1'h0;
  assign T_308 = T_305 & T_307;
  assign T_315 = T_304 ? 3'h4 : 3'h5;
  assign T_316 = T_300 ? {{1'd0}, 2'h3} : T_315;
  assign T_317 = T_296 ? {{1'd0}, 2'h2} : T_316;
  assign T_318 = T_292 ? {{2'd0}, 1'h1} : T_317;
  assign roq_deq_addr = T_288 ? {{2'd0}, 1'h0} : T_318;
  assign T_319 = roq_free_0 | roq_free_1;
  assign T_320 = T_319 | roq_free_2;
  assign T_321 = T_320 | roq_free_3;
  assign T_322 = T_321 | roq_free_4;
  assign T_323 = T_322 | roq_free_5;
  assign T_347 = T_288 | T_292;
  assign T_348 = T_347 | T_296;
  assign T_349 = T_348 | T_300;
  assign T_350 = T_349 | T_304;
  assign T_351 = T_350 | T_308;
  assign T_352 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_49 = {{2'd0}, 1'h0};
  assign GEN_3 = GEN_49 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_50 = {{2'd0}, 1'h1};
  assign GEN_4 = GEN_50 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_51 = {{1'd0}, 2'h2};
  assign GEN_5 = GEN_51 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_52 = {{1'd0}, 2'h3};
  assign GEN_6 = GEN_52 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_7 = 3'h4 == roq_enq_addr ? GEN_0 : roq_tags_4;
  assign GEN_8 = 3'h5 == roq_enq_addr ? GEN_0 : roq_tags_5;
  assign GEN_1 = 1'h0;
  assign GEN_9 = GEN_49 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_10 = GEN_50 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_11 = GEN_51 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_12 = GEN_52 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_13 = 3'h4 == roq_enq_addr ? GEN_1 : roq_free_4;
  assign GEN_14 = 3'h5 == roq_enq_addr ? GEN_1 : roq_free_5;
  assign GEN_23 = T_352 ? GEN_3 : roq_tags_0;
  assign GEN_24 = T_352 ? GEN_4 : roq_tags_1;
  assign GEN_25 = T_352 ? GEN_5 : roq_tags_2;
  assign GEN_26 = T_352 ? GEN_6 : roq_tags_3;
  assign GEN_27 = T_352 ? GEN_7 : roq_tags_4;
  assign GEN_28 = T_352 ? GEN_8 : roq_tags_5;
  assign GEN_30 = T_352 ? GEN_9 : roq_free_0;
  assign GEN_31 = T_352 ? GEN_10 : roq_free_1;
  assign GEN_32 = T_352 ? GEN_11 : roq_free_2;
  assign GEN_33 = T_352 ? GEN_12 : roq_free_3;
  assign GEN_34 = T_352 ? GEN_13 : roq_free_4;
  assign GEN_35 = T_352 ? GEN_14 : roq_free_5;
  assign GEN_2 = 1'h1;
  assign GEN_36 = GEN_49 == roq_deq_addr ? GEN_2 : GEN_30;
  assign GEN_37 = GEN_50 == roq_deq_addr ? GEN_2 : GEN_31;
  assign GEN_38 = GEN_51 == roq_deq_addr ? GEN_2 : GEN_32;
  assign GEN_39 = GEN_52 == roq_deq_addr ? GEN_2 : GEN_33;
  assign GEN_40 = 3'h4 == roq_deq_addr ? GEN_2 : GEN_34;
  assign GEN_41 = 3'h5 == roq_deq_addr ? GEN_2 : GEN_35;
  assign GEN_43 = io_deq_valid ? GEN_36 : GEN_30;
  assign GEN_44 = io_deq_valid ? GEN_37 : GEN_31;
  assign GEN_45 = io_deq_valid ? GEN_38 : GEN_32;
  assign GEN_46 = io_deq_valid ? GEN_39 : GEN_33;
  assign GEN_47 = io_deq_valid ? GEN_40 : GEN_34;
  assign GEN_48 = io_deq_valid ? GEN_41 : GEN_35;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data_addr_beat[initvar] = GEN_15[2:0];
  GEN_16 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    roq_data_subblock[initvar] = GEN_16[0:0];
  GEN_17 = {1{$random}};
  roq_tags_0 = GEN_17[4:0];
  GEN_18 = {1{$random}};
  roq_tags_1 = GEN_18[4:0];
  GEN_19 = {1{$random}};
  roq_tags_2 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  roq_tags_3 = GEN_20[4:0];
  GEN_21 = {1{$random}};
  roq_tags_4 = GEN_21[4:0];
  GEN_22 = {1{$random}};
  roq_tags_5 = GEN_22[4:0];
  GEN_29 = {1{$random}};
  roq_free_0 = GEN_29[0:0];
  GEN_42 = {1{$random}};
  roq_free_1 = GEN_42[0:0];
  GEN_53 = {1{$random}};
  roq_free_2 = GEN_53[0:0];
  GEN_54 = {1{$random}};
  roq_free_3 = GEN_54[0:0];
  GEN_55 = {1{$random}};
  roq_free_4 = GEN_55[0:0];
  GEN_56 = {1{$random}};
  roq_free_5 = GEN_56[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_addr_beat_T_353_en & roq_data_addr_beat_T_353_mask) begin
      roq_data_addr_beat[roq_data_addr_beat_T_353_addr] <= roq_data_addr_beat_T_353_data;
    end
    if(roq_data_subblock_T_353_en & roq_data_subblock_T_353_mask) begin
      roq_data_subblock[roq_data_subblock_T_353_addr] <= roq_data_subblock_T_353_data;
    end
    if(1'h0) begin
    end else begin
      roq_tags_0 <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      roq_tags_1 <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      roq_tags_2 <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      roq_tags_3 <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      roq_tags_4 <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      roq_tags_5 <= GEN_28;
    end
    if(reset) begin
      roq_free_0 <= T_270_0;
    end else begin
      roq_free_0 <= GEN_43;
    end
    if(reset) begin
      roq_free_1 <= T_270_1;
    end else begin
      roq_free_1 <= GEN_44;
    end
    if(reset) begin
      roq_free_2 <= T_270_2;
    end else begin
      roq_free_2 <= GEN_45;
    end
    if(reset) begin
      roq_free_3 <= T_270_3;
    end else begin
      roq_free_3 <= GEN_46;
    end
    if(reset) begin
      roq_free_4 <= T_270_4;
    end else begin
      roq_free_4 <= GEN_47;
    end
    if(reset) begin
      roq_free_5 <= T_270_5;
    end else begin
      roq_free_5 <= GEN_48;
    end
  end
endmodule
module NastiIOTileLinkIOIdMapper(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [2:0] io_req_tl_id,
  output [4:0] io_req_nasti_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_nasti_id,
  output [2:0] io_resp_tl_id
);
  assign io_req_ready = 1'h1;
  assign io_req_nasti_id = {{2'd0}, io_req_tl_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_tl_id = io_resp_nasti_id[2:0];
endmodule
module Arbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [2:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [2:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [2:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [2:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire [63:0] GEN_6;
  wire  GEN_7;
  wire  T_652;
  wire  T_654;
  wire  T_656;
  wire  T_657;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_654;
  assign io_out_valid = T_657;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_manager_xact_id : io_in_1_bits_manager_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_is_builtin_type : io_in_1_bits_is_builtin_type;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_g_type : io_in_1_bits_g_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_client_id : io_in_1_bits_client_id;
  assign T_652 = io_in_0_valid == 1'h0;
  assign T_654 = T_652 & io_out_ready;
  assign T_656 = T_652 == 1'h0;
  assign T_657 = T_656 | io_in_1_valid;
endmodule
module NastiIOTileLinkIOConverter(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [2:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [2:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_688_0;
  wire [2:0] T_688_1;
  wire [2:0] T_688_2;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_695;
  wire  T_696;
  wire  has_data;
  wire [2:0] T_705_0;
  wire [2:0] T_705_1;
  wire [2:0] T_705_2;
  wire  T_707;
  wire  T_708;
  wire  T_709;
  wire  T_712;
  wire  T_713;
  wire  is_subblock;
  wire [2:0] T_722_0;
  wire  T_724;
  wire  is_multibeat;
  wire  T_727;
  wire  T_728;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_15;
  wire  T_731;
  wire [2:0] GEN_6;
  wire [3:0] T_733;
  wire [2:0] T_734;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_736;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [4:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [4:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [2:0] get_id_mapper_io_req_tl_id;
  wire [4:0] get_id_mapper_io_req_nasti_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_nasti_id;
  wire [2:0] get_id_mapper_io_resp_tl_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [2:0] put_id_mapper_io_req_tl_id;
  wire [4:0] put_id_mapper_io_req_nasti_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_nasti_id;
  wire [2:0] put_id_mapper_io_resp_tl_id;
  wire [2:0] GEN_7;
  wire  T_761;
  wire  put_id_mask;
  wire  T_763;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_16;
  wire  aw_ready;
  wire  T_765;
  wire  T_767;
  wire  T_768;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_17;
  wire  T_771;
  wire [3:0] T_773;
  wire [2:0] T_774;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_775;
  wire  T_776;
  wire  T_778;
  wire  T_779;
  wire  T_780;
  wire  T_781;
  wire  T_783;
  wire  T_784;
  wire  T_785;
  wire  T_786;
  wire  T_787;
  wire  T_789;
  wire [2:0] T_790;
  wire [28:0] T_791;
  wire [31:0] T_792;
  wire [2:0] T_793;
  wire  T_803;
  wire [2:0] T_804;
  wire  T_805;
  wire [2:0] T_806;
  wire  T_807;
  wire [2:0] T_808;
  wire  T_809;
  wire [2:0] T_810;
  wire  T_811;
  wire [2:0] T_812;
  wire  T_813;
  wire [2:0] T_814;
  wire  T_815;
  wire [2:0] T_816;
  wire  T_817;
  wire [2:0] T_818;
  wire [2:0] T_820;
  wire [2:0] T_823;
  wire [31:0] T_843_addr;
  wire [7:0] T_843_len;
  wire [2:0] T_843_size;
  wire [1:0] T_843_burst;
  wire  T_843_lock;
  wire [3:0] T_843_cache;
  wire [2:0] T_843_prot;
  wire [3:0] T_843_qos;
  wire [3:0] T_843_region;
  wire [4:0] T_843_id;
  wire  T_843_user;
  wire  T_862;
  wire  T_863;
  wire  T_864;
  wire  T_865;
  wire [2:0] T_872;
  wire [31:0] T_885_addr;
  wire [7:0] T_885_len;
  wire [2:0] T_885_size;
  wire [1:0] T_885_burst;
  wire  T_885_lock;
  wire [3:0] T_885_cache;
  wire [2:0] T_885_prot;
  wire [3:0] T_885_qos;
  wire [3:0] T_885_region;
  wire [4:0] T_885_id;
  wire  T_885_user;
  wire  T_904;
  wire  T_906;
  wire  T_907;
  wire [7:0] GEN_9;
  wire [8:0] T_911;
  wire [7:0] T_912;
  wire [7:0] T_918_0;
  wire  T_921;
  wire  T_922;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire [7:0] T_927;
  wire [7:0] T_929;
  wire [7:0] T_930;
  wire  T_932;
  wire  T_933;
  wire [63:0] T_940_data;
  wire  T_940_last;
  wire [4:0] T_940_id;
  wire [7:0] T_940_strb;
  wire  T_940_user;
  wire  T_951;
  wire  T_952;
  wire  T_953;
  wire  T_954;
  wire  T_955;
  wire  T_959;
  wire  T_960;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  T_963;
  wire [2:0] T_971_0;
  wire [3:0] GEN_10;
  wire  T_973;
  wire  T_981_0;
  wire [3:0] GEN_11;
  wire  T_983;
  wire  T_986;
  wire  T_988;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_18;
  wire [3:0] T_993;
  wire [2:0] T_994;
  wire [2:0] GEN_5;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [2:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [2:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_1026;
  wire [2:0] T_1028;
  wire [2:0] T_1056_addr_beat;
  wire [2:0] T_1056_client_xact_id;
  wire  T_1056_manager_xact_id;
  wire  T_1056_is_builtin_type;
  wire [3:0] T_1056_g_type;
  wire [63:0] T_1056_data;
  wire  T_1084;
  wire  T_1085;
  wire  T_1086;
  wire  T_1088;
  wire  T_1091;
  wire  T_1092;
  wire  T_1094;
  wire [2:0] T_1127_addr_beat;
  wire [2:0] T_1127_client_xact_id;
  wire  T_1127_manager_xact_id;
  wire  T_1127_is_builtin_type;
  wire [3:0] T_1127_g_type;
  wire [63:0] T_1127_data;
  wire  T_1155;
  wire  T_1156;
  wire  T_1157;
  wire  T_1159;
  wire  T_1161;
  wire [1:0] GEN_13;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire  T_1167;
  wire  T_1169;
  wire  T_1171;
  wire  T_1172;
  wire  T_1173;
  wire  T_1175;
  reg [4:0] GEN_8;
  reg [31:0] GEN_19;
  reg  GEN_12;
  reg [31:0] GEN_20;
  reg  GEN_14;
  reg [31:0] GEN_21;
  ReorderQueue_37 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  NastiIOTileLinkIOIdMapper get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_tl_id(get_id_mapper_io_req_tl_id),
    .io_req_nasti_id(get_id_mapper_io_req_nasti_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_nasti_id(get_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(get_id_mapper_io_resp_tl_id)
  );
  NastiIOTileLinkIOIdMapper put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_tl_id(put_id_mapper_io_req_tl_id),
    .io_req_nasti_id(put_id_mapper_io_req_nasti_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_nasti_id(put_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(put_id_mapper_io_resp_tl_id)
  );
  Arbiter gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_955;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_865;
  assign io_nasti_aw_bits_addr = T_885_addr;
  assign io_nasti_aw_bits_len = T_885_len;
  assign io_nasti_aw_bits_size = T_885_size;
  assign io_nasti_aw_bits_burst = T_885_burst;
  assign io_nasti_aw_bits_lock = T_885_lock;
  assign io_nasti_aw_bits_cache = T_885_cache;
  assign io_nasti_aw_bits_prot = T_885_prot;
  assign io_nasti_aw_bits_qos = T_885_qos;
  assign io_nasti_aw_bits_region = T_885_region;
  assign io_nasti_aw_bits_id = T_885_id;
  assign io_nasti_aw_bits_user = T_885_user;
  assign io_nasti_w_valid = T_904;
  assign io_nasti_w_bits_data = T_940_data;
  assign io_nasti_w_bits_last = T_940_last;
  assign io_nasti_w_bits_id = T_940_id;
  assign io_nasti_w_bits_strb = T_940_strb;
  assign io_nasti_w_bits_user = T_940_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_789;
  assign io_nasti_ar_bits_addr = T_843_addr;
  assign io_nasti_ar_bits_len = T_843_len;
  assign io_nasti_ar_bits_size = T_843_size;
  assign io_nasti_ar_bits_burst = T_843_burst;
  assign io_nasti_ar_bits_lock = T_843_lock;
  assign io_nasti_ar_bits_cache = T_843_cache;
  assign io_nasti_ar_bits_prot = T_843_prot;
  assign io_nasti_ar_bits_qos = T_843_qos;
  assign io_nasti_ar_bits_region = T_843_region;
  assign io_nasti_ar_bits_id = T_843_id;
  assign io_nasti_ar_bits_user = T_843_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_688_0 = 3'h2;
  assign T_688_1 = 3'h3;
  assign T_688_2 = 3'h4;
  assign T_690 = T_688_0 == io_tl_acquire_bits_a_type;
  assign T_691 = T_688_1 == io_tl_acquire_bits_a_type;
  assign T_692 = T_688_2 == io_tl_acquire_bits_a_type;
  assign T_695 = T_690 | T_691;
  assign T_696 = T_695 | T_692;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_696;
  assign T_705_0 = 3'h2;
  assign T_705_1 = 3'h0;
  assign T_705_2 = 3'h4;
  assign T_707 = T_705_0 == io_tl_acquire_bits_a_type;
  assign T_708 = T_705_1 == io_tl_acquire_bits_a_type;
  assign T_709 = T_705_2 == io_tl_acquire_bits_a_type;
  assign T_712 = T_707 | T_708;
  assign T_713 = T_712 | T_709;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_713;
  assign T_722_0 = 3'h3;
  assign T_724 = T_722_0 == io_tl_acquire_bits_a_type;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_724;
  assign T_727 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_728 = T_727 & is_multibeat;
  assign T_731 = tl_cnt_out == 3'h7;
  assign GEN_6 = {{2'd0}, 1'h1};
  assign T_733 = tl_cnt_out + GEN_6;
  assign T_734 = T_733[2:0];
  assign GEN_0 = T_728 ? T_734 : tl_cnt_out;
  assign tl_wrap_out = T_728 & T_731;
  assign T_736 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_736;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_776;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id;
  assign roq_io_deq_valid = T_779;
  assign roq_io_deq_tag = io_nasti_r_bits_id;
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_781;
  assign get_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_783;
  assign get_id_mapper_io_resp_nasti_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_786;
  assign put_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_787;
  assign put_id_mapper_io_resp_nasti_id = io_nasti_b_bits_id;
  assign GEN_7 = {{2'd0}, 1'h0};
  assign T_761 = io_tl_acquire_bits_addr_beat == GEN_7;
  assign put_id_mask = is_subblock | T_761;
  assign T_763 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_763;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_765 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_767 = roq_io_deq_data_subblock == 1'h0;
  assign T_768 = T_765 & T_767;
  assign T_771 = nasti_cnt_out == 3'h7;
  assign T_773 = nasti_cnt_out + GEN_6;
  assign T_774 = T_773[2:0];
  assign GEN_1 = T_768 ? T_774 : nasti_cnt_out;
  assign nasti_wrap_out = T_768 & T_771;
  assign T_775 = get_valid & io_nasti_ar_ready;
  assign T_776 = T_775 & get_id_mapper_io_req_ready;
  assign T_778 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_779 = T_765 & T_778;
  assign T_780 = get_valid & roq_io_enq_ready;
  assign T_781 = T_780 & io_nasti_ar_ready;
  assign T_783 = T_765 & io_nasti_r_bits_last;
  assign T_784 = put_valid & aw_ready;
  assign T_785 = T_784 & io_nasti_w_ready;
  assign T_786 = T_785 & put_id_mask;
  assign T_787 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_789 = T_780 & get_id_mapper_io_req_ready;
  assign T_790 = io_tl_acquire_bits_union[11:9];
  assign T_791 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_792 = {T_791,T_790};
  assign T_793 = io_tl_acquire_bits_union[8:6];
  assign T_803 = 3'h7 == T_793;
  assign T_804 = T_803 ? {{1'd0}, 2'h3} : 3'h7;
  assign T_805 = 3'h3 == T_793;
  assign T_806 = T_805 ? {{1'd0}, 2'h3} : T_804;
  assign T_807 = 3'h6 == T_793;
  assign T_808 = T_807 ? {{1'd0}, 2'h2} : T_806;
  assign T_809 = 3'h2 == T_793;
  assign T_810 = T_809 ? {{1'd0}, 2'h2} : T_808;
  assign T_811 = 3'h5 == T_793;
  assign T_812 = T_811 ? {{2'd0}, 1'h1} : T_810;
  assign T_813 = 3'h1 == T_793;
  assign T_814 = T_813 ? {{2'd0}, 1'h1} : T_812;
  assign T_815 = 3'h4 == T_793;
  assign T_816 = T_815 ? {{2'd0}, 1'h0} : T_814;
  assign T_817 = 3'h0 == T_793;
  assign T_818 = T_817 ? {{2'd0}, 1'h0} : T_816;
  assign T_820 = is_subblock ? T_818 : {{1'd0}, 2'h3};
  assign T_823 = is_subblock ? {{2'd0}, 1'h0} : 3'h7;
  assign T_843_addr = T_792;
  assign T_843_len = {{5'd0}, T_823};
  assign T_843_size = T_820;
  assign T_843_burst = 2'h1;
  assign T_843_lock = 1'h0;
  assign T_843_cache = {{3'd0}, 1'h0};
  assign T_843_prot = {{2'd0}, 1'h0};
  assign T_843_qos = {{3'd0}, 1'h0};
  assign T_843_region = {{3'd0}, 1'h0};
  assign T_843_id = get_id_mapper_io_req_nasti_id;
  assign T_843_user = 1'h0;
  assign T_862 = w_inflight == 1'h0;
  assign T_863 = put_valid & io_nasti_w_ready;
  assign T_864 = T_863 & put_id_ready;
  assign T_865 = T_864 & T_862;
  assign T_872 = is_multibeat ? 3'h7 : {{2'd0}, 1'h0};
  assign T_885_addr = T_792;
  assign T_885_len = {{5'd0}, T_872};
  assign T_885_size = {{1'd0}, 2'h3};
  assign T_885_burst = 2'h1;
  assign T_885_lock = 1'h0;
  assign T_885_cache = 4'h0;
  assign T_885_prot = 3'h0;
  assign T_885_qos = 4'h0;
  assign T_885_region = 4'h0;
  assign T_885_id = put_id_mapper_io_req_nasti_id;
  assign T_885_user = 1'h0;
  assign T_904 = T_784 & put_id_ready;
  assign T_906 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_907 = io_tl_acquire_bits_is_builtin_type & T_906;
  assign GEN_9 = {{7'd0}, 1'h1};
  assign T_911 = 8'h0 - GEN_9;
  assign T_912 = T_911[7:0];
  assign T_918_0 = T_912;
  assign T_921 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_922 = io_tl_acquire_bits_is_builtin_type & T_921;
  assign T_924 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_925 = io_tl_acquire_bits_is_builtin_type & T_924;
  assign T_926 = T_922 | T_925;
  assign T_927 = io_tl_acquire_bits_union[8:1];
  assign T_929 = T_926 ? T_927 : {{7'd0}, 1'h0};
  assign T_930 = T_907 ? T_918_0 : T_929;
  assign T_932 = T_727 & is_subblock;
  assign T_933 = tl_wrap_out | T_932;
  assign T_940_data = io_tl_acquire_bits_data;
  assign T_940_last = T_933;
  assign T_940_id = GEN_8;
  assign T_940_strb = T_930;
  assign T_940_user = 1'h0;
  assign T_951 = aw_ready & io_nasti_w_ready;
  assign T_952 = T_951 & put_id_ready;
  assign T_953 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_954 = T_953 & get_id_mapper_io_req_ready;
  assign T_955 = has_data ? T_952 : T_954;
  assign T_959 = T_862 & T_727;
  assign T_960 = T_959 & is_multibeat;
  assign GEN_2 = T_960 ? 1'h1 : w_inflight;
  assign GEN_3 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_4 = w_inflight ? GEN_3 : GEN_2;
  assign T_963 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_971_0 = 3'h5;
  assign GEN_10 = {{1'd0}, T_971_0};
  assign T_973 = GEN_10 == io_tl_grant_bits_g_type;
  assign T_981_0 = 1'h0;
  assign GEN_11 = {{3'd0}, T_981_0};
  assign T_983 = GEN_11 == io_tl_grant_bits_g_type;
  assign T_986 = io_tl_grant_bits_is_builtin_type ? T_973 : T_983;
  assign T_988 = T_963 & T_986;
  assign T_993 = tl_cnt_in + GEN_6;
  assign T_994 = T_993[2:0];
  assign GEN_5 = T_988 ? T_994 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_1056_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_1056_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_1056_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_1056_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_1056_g_type;
  assign gnt_arb_io_in_0_bits_data = T_1056_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_12;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1127_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1127_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1127_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1127_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1127_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1127_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_14;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_1026 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_1028 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_1056_addr_beat = T_1028;
  assign T_1056_client_xact_id = get_id_mapper_io_resp_tl_id;
  assign T_1056_manager_xact_id = 1'h0;
  assign T_1056_is_builtin_type = 1'h1;
  assign T_1056_g_type = {{1'd0}, T_1026};
  assign T_1056_data = io_nasti_r_bits_data;
  assign T_1084 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_1085 = T_1084 | roq_io_deq_matches;
  assign T_1086 = T_1085 | reset;
  assign T_1088 = T_1086 == 1'h0;
  assign T_1091 = T_1084 | get_id_mapper_io_resp_matches;
  assign T_1092 = T_1091 | reset;
  assign T_1094 = T_1092 == 1'h0;
  assign T_1127_addr_beat = {{2'd0}, 1'h0};
  assign T_1127_client_xact_id = put_id_mapper_io_resp_tl_id;
  assign T_1127_manager_xact_id = 1'h0;
  assign T_1127_is_builtin_type = 1'h1;
  assign T_1127_g_type = {{1'd0}, 3'h3};
  assign T_1127_data = {{63'd0}, 1'h0};
  assign T_1155 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1156 = T_1155 | put_id_mapper_io_resp_matches;
  assign T_1157 = T_1156 | reset;
  assign T_1159 = T_1157 == 1'h0;
  assign T_1161 = io_nasti_r_valid == 1'h0;
  assign GEN_13 = {{1'd0}, 1'h0};
  assign T_1163 = io_nasti_r_bits_resp == GEN_13;
  assign T_1164 = T_1161 | T_1163;
  assign T_1165 = T_1164 | reset;
  assign T_1167 = T_1165 == 1'h0;
  assign T_1169 = io_nasti_b_valid == 1'h0;
  assign T_1171 = io_nasti_b_bits_resp == GEN_13;
  assign T_1172 = T_1169 | T_1171;
  assign T_1173 = T_1172 | reset;
  assign T_1175 = T_1173 == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  tl_cnt_out = GEN_15[2:0];
  GEN_16 = {1{$random}};
  w_inflight = GEN_16[0:0];
  GEN_17 = {1{$random}};
  nasti_cnt_out = GEN_17[2:0];
  GEN_18 = {1{$random}};
  tl_cnt_in = GEN_18[2:0];
  GEN_19 = {1{$random}};
  GEN_8 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  GEN_12 = GEN_20[0:0];
  GEN_21 = {1{$random}};
  GEN_14 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      tl_cnt_out <= GEN_0;
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      w_inflight <= GEN_4;
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      nasti_cnt_out <= GEN_1;
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      tl_cnt_in <= GEN_5;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1088) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:609 assert(!gnt_arb.io.in(0).valid || roq.io.deq.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1088) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1094) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:610 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1094) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1159) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:621 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1159) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1167) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at converters.scala:623 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1167) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1175) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at converters.scala:624 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1175) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_39(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [7:0] io_enq_bits_len,
  input  [2:0] io_enq_bits_size,
  input  [1:0] io_enq_bits_burst,
  input   io_enq_bits_lock,
  input  [3:0] io_enq_bits_cache,
  input  [2:0] io_enq_bits_prot,
  input  [3:0] io_enq_bits_qos,
  input  [3:0] io_enq_bits_region,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [7:0] io_deq_bits_len,
  output [2:0] io_deq_bits_size,
  output [1:0] io_deq_bits_burst,
  output  io_deq_bits_lock,
  output [3:0] io_deq_bits_cache,
  output [2:0] io_deq_bits_prot,
  output [3:0] io_deq_bits_qos,
  output [3:0] io_deq_bits_region,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [31:0] ram_addr [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_addr_T_144_data;
  wire  ram_addr_T_144_addr;
  wire  ram_addr_T_144_en;
  wire [31:0] ram_addr_T_125_data;
  wire  ram_addr_T_125_addr;
  wire  ram_addr_T_125_mask;
  wire  ram_addr_T_125_en;
  reg [7:0] ram_len [0:0];
  reg [31:0] GEN_1;
  wire [7:0] ram_len_T_144_data;
  wire  ram_len_T_144_addr;
  wire  ram_len_T_144_en;
  wire [7:0] ram_len_T_125_data;
  wire  ram_len_T_125_addr;
  wire  ram_len_T_125_mask;
  wire  ram_len_T_125_en;
  reg [2:0] ram_size [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_size_T_144_data;
  wire  ram_size_T_144_addr;
  wire  ram_size_T_144_en;
  wire [2:0] ram_size_T_125_data;
  wire  ram_size_T_125_addr;
  wire  ram_size_T_125_mask;
  wire  ram_size_T_125_en;
  reg [1:0] ram_burst [0:0];
  reg [31:0] GEN_3;
  wire [1:0] ram_burst_T_144_data;
  wire  ram_burst_T_144_addr;
  wire  ram_burst_T_144_en;
  wire [1:0] ram_burst_T_125_data;
  wire  ram_burst_T_125_addr;
  wire  ram_burst_T_125_mask;
  wire  ram_burst_T_125_en;
  reg  ram_lock [0:0];
  reg [31:0] GEN_4;
  wire  ram_lock_T_144_data;
  wire  ram_lock_T_144_addr;
  wire  ram_lock_T_144_en;
  wire  ram_lock_T_125_data;
  wire  ram_lock_T_125_addr;
  wire  ram_lock_T_125_mask;
  wire  ram_lock_T_125_en;
  reg [3:0] ram_cache [0:0];
  reg [31:0] GEN_5;
  wire [3:0] ram_cache_T_144_data;
  wire  ram_cache_T_144_addr;
  wire  ram_cache_T_144_en;
  wire [3:0] ram_cache_T_125_data;
  wire  ram_cache_T_125_addr;
  wire  ram_cache_T_125_mask;
  wire  ram_cache_T_125_en;
  reg [2:0] ram_prot [0:0];
  reg [31:0] GEN_6;
  wire [2:0] ram_prot_T_144_data;
  wire  ram_prot_T_144_addr;
  wire  ram_prot_T_144_en;
  wire [2:0] ram_prot_T_125_data;
  wire  ram_prot_T_125_addr;
  wire  ram_prot_T_125_mask;
  wire  ram_prot_T_125_en;
  reg [3:0] ram_qos [0:0];
  reg [31:0] GEN_7;
  wire [3:0] ram_qos_T_144_data;
  wire  ram_qos_T_144_addr;
  wire  ram_qos_T_144_en;
  wire [3:0] ram_qos_T_125_data;
  wire  ram_qos_T_125_addr;
  wire  ram_qos_T_125_mask;
  wire  ram_qos_T_125_en;
  reg [3:0] ram_region [0:0];
  reg [31:0] GEN_8;
  wire [3:0] ram_region_T_144_data;
  wire  ram_region_T_144_addr;
  wire  ram_region_T_144_en;
  wire [3:0] ram_region_T_125_data;
  wire  ram_region_T_125_addr;
  wire  ram_region_T_125_mask;
  wire  ram_region_T_125_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_9;
  wire [4:0] ram_id_T_144_data;
  wire  ram_id_T_144_addr;
  wire  ram_id_T_144_en;
  wire [4:0] ram_id_T_125_data;
  wire  ram_id_T_125_addr;
  wire  ram_id_T_125_mask;
  wire  ram_id_T_125_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_10;
  wire  ram_user_T_144_data;
  wire  ram_user_T_144_addr;
  wire  ram_user_T_144_en;
  wire  ram_user_T_125_data;
  wire  ram_user_T_125_addr;
  wire  ram_user_T_125_mask;
  wire  ram_user_T_125_en;
  reg  maybe_full;
  reg [31:0] GEN_11;
  wire  T_122;
  wire  T_123;
  wire  do_enq;
  wire  T_124;
  wire  do_deq;
  wire  T_139;
  wire  GEN_25;
  wire  T_141;
  wire [1:0] T_156;
  wire  ptr_diff;
  wire [1:0] T_158;
  assign io_enq_ready = T_122;
  assign io_deq_valid = T_141;
  assign io_deq_bits_addr = ram_addr_T_144_data;
  assign io_deq_bits_len = ram_len_T_144_data;
  assign io_deq_bits_size = ram_size_T_144_data;
  assign io_deq_bits_burst = ram_burst_T_144_data;
  assign io_deq_bits_lock = ram_lock_T_144_data;
  assign io_deq_bits_cache = ram_cache_T_144_data;
  assign io_deq_bits_prot = ram_prot_T_144_data;
  assign io_deq_bits_qos = ram_qos_T_144_data;
  assign io_deq_bits_region = ram_region_T_144_data;
  assign io_deq_bits_id = ram_id_T_144_data;
  assign io_deq_bits_user = ram_user_T_144_data;
  assign io_count = T_158[0];
  assign ram_addr_T_144_addr = 1'h0;
  assign ram_addr_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_T_144_data = ram_addr[ram_addr_T_144_addr];
  `else
  assign ram_addr_T_144_data = ram_addr_T_144_addr >= 1'h1 ? $random : ram_addr[ram_addr_T_144_addr];
  `endif
  assign ram_addr_T_125_data = io_enq_bits_addr;
  assign ram_addr_T_125_addr = 1'h0;
  assign ram_addr_T_125_mask = do_enq;
  assign ram_addr_T_125_en = do_enq;
  assign ram_len_T_144_addr = 1'h0;
  assign ram_len_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_len_T_144_data = ram_len[ram_len_T_144_addr];
  `else
  assign ram_len_T_144_data = ram_len_T_144_addr >= 1'h1 ? $random : ram_len[ram_len_T_144_addr];
  `endif
  assign ram_len_T_125_data = io_enq_bits_len;
  assign ram_len_T_125_addr = 1'h0;
  assign ram_len_T_125_mask = do_enq;
  assign ram_len_T_125_en = do_enq;
  assign ram_size_T_144_addr = 1'h0;
  assign ram_size_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_size_T_144_data = ram_size[ram_size_T_144_addr];
  `else
  assign ram_size_T_144_data = ram_size_T_144_addr >= 1'h1 ? $random : ram_size[ram_size_T_144_addr];
  `endif
  assign ram_size_T_125_data = io_enq_bits_size;
  assign ram_size_T_125_addr = 1'h0;
  assign ram_size_T_125_mask = do_enq;
  assign ram_size_T_125_en = do_enq;
  assign ram_burst_T_144_addr = 1'h0;
  assign ram_burst_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_burst_T_144_data = ram_burst[ram_burst_T_144_addr];
  `else
  assign ram_burst_T_144_data = ram_burst_T_144_addr >= 1'h1 ? $random : ram_burst[ram_burst_T_144_addr];
  `endif
  assign ram_burst_T_125_data = io_enq_bits_burst;
  assign ram_burst_T_125_addr = 1'h0;
  assign ram_burst_T_125_mask = do_enq;
  assign ram_burst_T_125_en = do_enq;
  assign ram_lock_T_144_addr = 1'h0;
  assign ram_lock_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_lock_T_144_data = ram_lock[ram_lock_T_144_addr];
  `else
  assign ram_lock_T_144_data = ram_lock_T_144_addr >= 1'h1 ? $random : ram_lock[ram_lock_T_144_addr];
  `endif
  assign ram_lock_T_125_data = io_enq_bits_lock;
  assign ram_lock_T_125_addr = 1'h0;
  assign ram_lock_T_125_mask = do_enq;
  assign ram_lock_T_125_en = do_enq;
  assign ram_cache_T_144_addr = 1'h0;
  assign ram_cache_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_cache_T_144_data = ram_cache[ram_cache_T_144_addr];
  `else
  assign ram_cache_T_144_data = ram_cache_T_144_addr >= 1'h1 ? $random : ram_cache[ram_cache_T_144_addr];
  `endif
  assign ram_cache_T_125_data = io_enq_bits_cache;
  assign ram_cache_T_125_addr = 1'h0;
  assign ram_cache_T_125_mask = do_enq;
  assign ram_cache_T_125_en = do_enq;
  assign ram_prot_T_144_addr = 1'h0;
  assign ram_prot_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_prot_T_144_data = ram_prot[ram_prot_T_144_addr];
  `else
  assign ram_prot_T_144_data = ram_prot_T_144_addr >= 1'h1 ? $random : ram_prot[ram_prot_T_144_addr];
  `endif
  assign ram_prot_T_125_data = io_enq_bits_prot;
  assign ram_prot_T_125_addr = 1'h0;
  assign ram_prot_T_125_mask = do_enq;
  assign ram_prot_T_125_en = do_enq;
  assign ram_qos_T_144_addr = 1'h0;
  assign ram_qos_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_qos_T_144_data = ram_qos[ram_qos_T_144_addr];
  `else
  assign ram_qos_T_144_data = ram_qos_T_144_addr >= 1'h1 ? $random : ram_qos[ram_qos_T_144_addr];
  `endif
  assign ram_qos_T_125_data = io_enq_bits_qos;
  assign ram_qos_T_125_addr = 1'h0;
  assign ram_qos_T_125_mask = do_enq;
  assign ram_qos_T_125_en = do_enq;
  assign ram_region_T_144_addr = 1'h0;
  assign ram_region_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_region_T_144_data = ram_region[ram_region_T_144_addr];
  `else
  assign ram_region_T_144_data = ram_region_T_144_addr >= 1'h1 ? $random : ram_region[ram_region_T_144_addr];
  `endif
  assign ram_region_T_125_data = io_enq_bits_region;
  assign ram_region_T_125_addr = 1'h0;
  assign ram_region_T_125_mask = do_enq;
  assign ram_region_T_125_en = do_enq;
  assign ram_id_T_144_addr = 1'h0;
  assign ram_id_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_144_data = ram_id[ram_id_T_144_addr];
  `else
  assign ram_id_T_144_data = ram_id_T_144_addr >= 1'h1 ? $random : ram_id[ram_id_T_144_addr];
  `endif
  assign ram_id_T_125_data = io_enq_bits_id;
  assign ram_id_T_125_addr = 1'h0;
  assign ram_id_T_125_mask = do_enq;
  assign ram_id_T_125_en = do_enq;
  assign ram_user_T_144_addr = 1'h0;
  assign ram_user_T_144_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_144_data = ram_user[ram_user_T_144_addr];
  `else
  assign ram_user_T_144_data = ram_user_T_144_addr >= 1'h1 ? $random : ram_user[ram_user_T_144_addr];
  `endif
  assign ram_user_T_125_data = io_enq_bits_user;
  assign ram_user_T_125_addr = 1'h0;
  assign ram_user_T_125_mask = do_enq;
  assign ram_user_T_125_en = do_enq;
  assign T_122 = maybe_full == 1'h0;
  assign T_123 = io_enq_ready & io_enq_valid;
  assign do_enq = T_123;
  assign T_124 = io_deq_ready & io_deq_valid;
  assign do_deq = T_124;
  assign T_139 = do_enq != do_deq;
  assign GEN_25 = T_139 ? do_enq : maybe_full;
  assign T_141 = T_122 == 1'h0;
  assign T_156 = 1'h0 - 1'h0;
  assign ptr_diff = T_156[0:0];
  assign T_158 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[31:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = GEN_1[7:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_size[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_burst[initvar] = GEN_3[1:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_lock[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_cache[initvar] = GEN_5[3:0];
  GEN_6 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_prot[initvar] = GEN_6[2:0];
  GEN_7 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_qos[initvar] = GEN_7[3:0];
  GEN_8 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_region[initvar] = GEN_8[3:0];
  GEN_9 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_9[4:0];
  GEN_10 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_10[0:0];
  GEN_11 = {1{$random}};
  maybe_full = GEN_11[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_125_en & ram_addr_T_125_mask) begin
      ram_addr[ram_addr_T_125_addr] <= ram_addr_T_125_data;
    end
    if(ram_len_T_125_en & ram_len_T_125_mask) begin
      ram_len[ram_len_T_125_addr] <= ram_len_T_125_data;
    end
    if(ram_size_T_125_en & ram_size_T_125_mask) begin
      ram_size[ram_size_T_125_addr] <= ram_size_T_125_data;
    end
    if(ram_burst_T_125_en & ram_burst_T_125_mask) begin
      ram_burst[ram_burst_T_125_addr] <= ram_burst_T_125_data;
    end
    if(ram_lock_T_125_en & ram_lock_T_125_mask) begin
      ram_lock[ram_lock_T_125_addr] <= ram_lock_T_125_data;
    end
    if(ram_cache_T_125_en & ram_cache_T_125_mask) begin
      ram_cache[ram_cache_T_125_addr] <= ram_cache_T_125_data;
    end
    if(ram_prot_T_125_en & ram_prot_T_125_mask) begin
      ram_prot[ram_prot_T_125_addr] <= ram_prot_T_125_data;
    end
    if(ram_qos_T_125_en & ram_qos_T_125_mask) begin
      ram_qos[ram_qos_T_125_addr] <= ram_qos_T_125_data;
    end
    if(ram_region_T_125_en & ram_region_T_125_mask) begin
      ram_region[ram_region_T_125_addr] <= ram_region_T_125_data;
    end
    if(ram_id_T_125_en & ram_id_T_125_mask) begin
      ram_id[ram_id_T_125_addr] <= ram_id_T_125_data;
    end
    if(ram_user_T_125_en & ram_user_T_125_mask) begin
      ram_user[ram_user_T_125_addr] <= ram_user_T_125_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_25;
    end
  end
endmodule
module Queue_41(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input  [7:0] io_enq_bits_strb,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output [7:0] io_deq_bits_strb,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_0;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_1;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_2;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg [7:0] ram_strb [0:1];
  reg [31:0] GEN_3;
  wire [7:0] ram_strb_T_94_data;
  wire  ram_strb_T_94_addr;
  wire  ram_strb_T_94_en;
  wire [7:0] ram_strb_T_73_data;
  wire  ram_strb_T_73_addr;
  wire  ram_strb_T_73_mask;
  wire  ram_strb_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_strb = ram_strb_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  `else
  assign ram_data_T_94_data = ram_data_T_94_addr >= 2'h2 ? $random : ram_data[ram_data_T_94_addr];
  `endif
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  `else
  assign ram_last_T_94_data = ram_last_T_94_addr >= 2'h2 ? $random : ram_last[ram_last_T_94_addr];
  `endif
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  `else
  assign ram_id_T_94_data = ram_id_T_94_addr >= 2'h2 ? $random : ram_id[ram_id_T_94_addr];
  `endif
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_strb_T_94_addr = T_67;
  assign ram_strb_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_strb_T_94_data = ram_strb[ram_strb_T_94_addr];
  `else
  assign ram_strb_T_94_data = ram_strb_T_94_addr >= 2'h2 ? $random : ram_strb[ram_strb_T_94_addr];
  `endif
  assign ram_strb_T_73_data = io_enq_bits_strb;
  assign ram_strb_T_73_addr = T_65;
  assign ram_strb_T_73_mask = do_enq;
  assign ram_strb_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  `else
  assign ram_user_T_94_data = ram_user_T_94_addr >= 2'h2 ? $random : ram_user[ram_user_T_94_addr];
  `endif
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_0[63:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_2[4:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_strb[initvar] = GEN_3[7:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_strb_T_73_en & ram_strb_T_73_mask) begin
      ram_strb[ram_strb_T_73_addr] <= ram_strb_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      T_65 <= GEN_13;
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      T_67 <= GEN_14;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_15;
    end
  end
endmodule
module Queue_42(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [63:0] io_enq_bits_data,
  input   io_enq_bits_last,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [63:0] io_deq_bits_data,
  output  io_deq_bits_last,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output [1:0] io_count
);
  reg [1:0] ram_resp [0:1];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_94_data;
  wire  ram_resp_T_94_addr;
  wire  ram_resp_T_94_en;
  wire [1:0] ram_resp_T_73_data;
  wire  ram_resp_T_73_addr;
  wire  ram_resp_T_73_mask;
  wire  ram_resp_T_73_en;
  reg [63:0] ram_data [0:1];
  reg [63:0] GEN_1;
  wire [63:0] ram_data_T_94_data;
  wire  ram_data_T_94_addr;
  wire  ram_data_T_94_en;
  wire [63:0] ram_data_T_73_data;
  wire  ram_data_T_73_addr;
  wire  ram_data_T_73_mask;
  wire  ram_data_T_73_en;
  reg  ram_last [0:1];
  reg [31:0] GEN_2;
  wire  ram_last_T_94_data;
  wire  ram_last_T_94_addr;
  wire  ram_last_T_94_en;
  wire  ram_last_T_73_data;
  wire  ram_last_T_73_addr;
  wire  ram_last_T_73_mask;
  wire  ram_last_T_73_en;
  reg [4:0] ram_id [0:1];
  reg [31:0] GEN_3;
  wire [4:0] ram_id_T_94_data;
  wire  ram_id_T_94_addr;
  wire  ram_id_T_94_en;
  wire [4:0] ram_id_T_73_data;
  wire  ram_id_T_73_addr;
  wire  ram_id_T_73_mask;
  wire  ram_id_T_73_en;
  reg  ram_user [0:1];
  reg [31:0] GEN_4;
  wire  ram_user_T_94_data;
  wire  ram_user_T_94_addr;
  wire  ram_user_T_94_en;
  wire  ram_user_T_73_data;
  wire  ram_user_T_73_addr;
  wire  ram_user_T_73_mask;
  wire  ram_user_T_73_en;
  reg  T_65;
  reg [31:0] GEN_5;
  reg  T_67;
  reg [31:0] GEN_6;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  ptr_match;
  wire  T_70;
  wire  empty;
  wire  full;
  wire  T_71;
  wire  do_enq;
  wire  T_72;
  wire  do_deq;
  wire [1:0] T_82;
  wire  T_83;
  wire  GEN_13;
  wire [1:0] T_87;
  wire  T_88;
  wire  GEN_14;
  wire  T_89;
  wire  GEN_15;
  wire  T_91;
  wire  T_93;
  wire [1:0] T_100;
  wire  ptr_diff;
  wire  T_101;
  wire [1:0] T_102;
  assign io_enq_ready = T_93;
  assign io_deq_valid = T_91;
  assign io_deq_bits_resp = ram_resp_T_94_data;
  assign io_deq_bits_data = ram_data_T_94_data;
  assign io_deq_bits_last = ram_last_T_94_data;
  assign io_deq_bits_id = ram_id_T_94_data;
  assign io_deq_bits_user = ram_user_T_94_data;
  assign io_count = T_102;
  assign ram_resp_T_94_addr = T_67;
  assign ram_resp_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_resp_T_94_data = ram_resp[ram_resp_T_94_addr];
  `else
  assign ram_resp_T_94_data = ram_resp_T_94_addr >= 2'h2 ? $random : ram_resp[ram_resp_T_94_addr];
  `endif
  assign ram_resp_T_73_data = io_enq_bits_resp;
  assign ram_resp_T_73_addr = T_65;
  assign ram_resp_T_73_mask = do_enq;
  assign ram_resp_T_73_en = do_enq;
  assign ram_data_T_94_addr = T_67;
  assign ram_data_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_94_data = ram_data[ram_data_T_94_addr];
  `else
  assign ram_data_T_94_data = ram_data_T_94_addr >= 2'h2 ? $random : ram_data[ram_data_T_94_addr];
  `endif
  assign ram_data_T_73_data = io_enq_bits_data;
  assign ram_data_T_73_addr = T_65;
  assign ram_data_T_73_mask = do_enq;
  assign ram_data_T_73_en = do_enq;
  assign ram_last_T_94_addr = T_67;
  assign ram_last_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_last_T_94_data = ram_last[ram_last_T_94_addr];
  `else
  assign ram_last_T_94_data = ram_last_T_94_addr >= 2'h2 ? $random : ram_last[ram_last_T_94_addr];
  `endif
  assign ram_last_T_73_data = io_enq_bits_last;
  assign ram_last_T_73_addr = T_65;
  assign ram_last_T_73_mask = do_enq;
  assign ram_last_T_73_en = do_enq;
  assign ram_id_T_94_addr = T_67;
  assign ram_id_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_94_data = ram_id[ram_id_T_94_addr];
  `else
  assign ram_id_T_94_data = ram_id_T_94_addr >= 2'h2 ? $random : ram_id[ram_id_T_94_addr];
  `endif
  assign ram_id_T_73_data = io_enq_bits_id;
  assign ram_id_T_73_addr = T_65;
  assign ram_id_T_73_mask = do_enq;
  assign ram_id_T_73_en = do_enq;
  assign ram_user_T_94_addr = T_67;
  assign ram_user_T_94_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_94_data = ram_user[ram_user_T_94_addr];
  `else
  assign ram_user_T_94_data = ram_user_T_94_addr >= 2'h2 ? $random : ram_user[ram_user_T_94_addr];
  `endif
  assign ram_user_T_73_data = io_enq_bits_user;
  assign ram_user_T_73_addr = T_65;
  assign ram_user_T_73_mask = do_enq;
  assign ram_user_T_73_en = do_enq;
  assign ptr_match = T_65 == T_67;
  assign T_70 = maybe_full == 1'h0;
  assign empty = ptr_match & T_70;
  assign full = ptr_match & maybe_full;
  assign T_71 = io_enq_ready & io_enq_valid;
  assign do_enq = T_71;
  assign T_72 = io_deq_ready & io_deq_valid;
  assign do_deq = T_72;
  assign T_82 = T_65 + 1'h1;
  assign T_83 = T_82[0:0];
  assign GEN_13 = do_enq ? T_83 : T_65;
  assign T_87 = T_67 + 1'h1;
  assign T_88 = T_87[0:0];
  assign GEN_14 = do_deq ? T_88 : T_67;
  assign T_89 = do_enq != do_deq;
  assign GEN_15 = T_89 ? do_enq : maybe_full;
  assign T_91 = empty == 1'h0;
  assign T_93 = full == 1'h0;
  assign T_100 = T_65 - T_67;
  assign ptr_diff = T_100[0:0];
  assign T_101 = maybe_full & ptr_match;
  assign T_102 = {T_101,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_data[initvar] = GEN_1[63:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_last[initvar] = GEN_2[0:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_id[initvar] = GEN_3[4:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 2; initvar = initvar+1)
    ram_user[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  T_65 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  T_67 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_73_en & ram_resp_T_73_mask) begin
      ram_resp[ram_resp_T_73_addr] <= ram_resp_T_73_data;
    end
    if(ram_data_T_73_en & ram_data_T_73_mask) begin
      ram_data[ram_data_T_73_addr] <= ram_data_T_73_data;
    end
    if(ram_last_T_73_en & ram_last_T_73_mask) begin
      ram_last[ram_last_T_73_addr] <= ram_last_T_73_data;
    end
    if(ram_id_T_73_en & ram_id_T_73_mask) begin
      ram_id[ram_id_T_73_addr] <= ram_id_T_73_data;
    end
    if(ram_user_T_73_en & ram_user_T_73_mask) begin
      ram_user[ram_user_T_73_addr] <= ram_user_T_73_data;
    end
    if(reset) begin
      T_65 <= 1'h0;
    end else begin
      T_65 <= GEN_13;
    end
    if(reset) begin
      T_67 <= 1'h0;
    end else begin
      T_67 <= GEN_14;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_15;
    end
  end
endmodule
module Queue_43(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [1:0] io_enq_bits_resp,
  input  [4:0] io_enq_bits_id,
  input   io_enq_bits_user,
  input   io_deq_ready,
  output  io_deq_valid,
  output [1:0] io_deq_bits_resp,
  output [4:0] io_deq_bits_id,
  output  io_deq_bits_user,
  output  io_count
);
  reg [1:0] ram_resp [0:0];
  reg [31:0] GEN_0;
  wire [1:0] ram_resp_T_64_data;
  wire  ram_resp_T_64_addr;
  wire  ram_resp_T_64_en;
  wire [1:0] ram_resp_T_53_data;
  wire  ram_resp_T_53_addr;
  wire  ram_resp_T_53_mask;
  wire  ram_resp_T_53_en;
  reg [4:0] ram_id [0:0];
  reg [31:0] GEN_1;
  wire [4:0] ram_id_T_64_data;
  wire  ram_id_T_64_addr;
  wire  ram_id_T_64_en;
  wire [4:0] ram_id_T_53_data;
  wire  ram_id_T_53_addr;
  wire  ram_id_T_53_mask;
  wire  ram_id_T_53_en;
  reg  ram_user [0:0];
  reg [31:0] GEN_2;
  wire  ram_user_T_64_data;
  wire  ram_user_T_64_addr;
  wire  ram_user_T_64_en;
  wire  ram_user_T_53_data;
  wire  ram_user_T_53_addr;
  wire  ram_user_T_53_mask;
  wire  ram_user_T_53_en;
  reg  maybe_full;
  reg [31:0] GEN_3;
  wire  T_50;
  wire  T_51;
  wire  do_enq;
  wire  T_52;
  wire  do_deq;
  wire  T_59;
  wire  GEN_9;
  wire  T_61;
  wire [1:0] T_68;
  wire  ptr_diff;
  wire [1:0] T_70;
  assign io_enq_ready = T_50;
  assign io_deq_valid = T_61;
  assign io_deq_bits_resp = ram_resp_T_64_data;
  assign io_deq_bits_id = ram_id_T_64_data;
  assign io_deq_bits_user = ram_user_T_64_data;
  assign io_count = T_70[0];
  assign ram_resp_T_64_addr = 1'h0;
  assign ram_resp_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_resp_T_64_data = ram_resp[ram_resp_T_64_addr];
  `else
  assign ram_resp_T_64_data = ram_resp_T_64_addr >= 1'h1 ? $random : ram_resp[ram_resp_T_64_addr];
  `endif
  assign ram_resp_T_53_data = io_enq_bits_resp;
  assign ram_resp_T_53_addr = 1'h0;
  assign ram_resp_T_53_mask = do_enq;
  assign ram_resp_T_53_en = do_enq;
  assign ram_id_T_64_addr = 1'h0;
  assign ram_id_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_id_T_64_data = ram_id[ram_id_T_64_addr];
  `else
  assign ram_id_T_64_data = ram_id_T_64_addr >= 1'h1 ? $random : ram_id[ram_id_T_64_addr];
  `endif
  assign ram_id_T_53_data = io_enq_bits_id;
  assign ram_id_T_53_addr = 1'h0;
  assign ram_id_T_53_mask = do_enq;
  assign ram_id_T_53_en = do_enq;
  assign ram_user_T_64_addr = 1'h0;
  assign ram_user_T_64_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_user_T_64_data = ram_user[ram_user_T_64_addr];
  `else
  assign ram_user_T_64_data = ram_user_T_64_addr >= 1'h1 ? $random : ram_user[ram_user_T_64_addr];
  `endif
  assign ram_user_T_53_data = io_enq_bits_user;
  assign ram_user_T_53_addr = 1'h0;
  assign ram_user_T_53_mask = do_enq;
  assign ram_user_T_53_en = do_enq;
  assign T_50 = maybe_full == 1'h0;
  assign T_51 = io_enq_ready & io_enq_valid;
  assign do_enq = T_51;
  assign T_52 = io_deq_ready & io_deq_valid;
  assign do_deq = T_52;
  assign T_59 = do_enq != do_deq;
  assign GEN_9 = T_59 ? do_enq : maybe_full;
  assign T_61 = T_50 == 1'h0;
  assign T_68 = 1'h0 - 1'h0;
  assign ptr_diff = T_68[0:0];
  assign T_70 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_resp[initvar] = GEN_0[1:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_id[initvar] = GEN_1[4:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_user[initvar] = GEN_2[0:0];
  GEN_3 = {1{$random}};
  maybe_full = GEN_3[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_resp_T_53_en & ram_resp_T_53_mask) begin
      ram_resp[ram_resp_T_53_addr] <= ram_resp_T_53_data;
    end
    if(ram_id_T_53_en & ram_id_T_53_mask) begin
      ram_id[ram_id_T_53_addr] <= ram_id_T_53_data;
    end
    if(ram_user_T_53_en & ram_user_T_53_mask) begin
      ram_user[ram_user_T_53_addr] <= ram_user_T_53_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_9;
    end
  end
endmodule
module OuterMemorySystem(
  input   clk,
  input   reset,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input  [1:0] io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_cached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [2:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  output  io_htif_uncached_acquire_ready,
  input   io_htif_uncached_acquire_valid,
  input  [25:0] io_htif_uncached_acquire_bits_addr_block,
  input  [1:0] io_htif_uncached_acquire_bits_client_xact_id,
  input  [2:0] io_htif_uncached_acquire_bits_addr_beat,
  input   io_htif_uncached_acquire_bits_is_builtin_type,
  input  [2:0] io_htif_uncached_acquire_bits_a_type,
  input  [11:0] io_htif_uncached_acquire_bits_union,
  input  [63:0] io_htif_uncached_acquire_bits_data,
  input   io_htif_uncached_grant_ready,
  output  io_htif_uncached_grant_valid,
  output [2:0] io_htif_uncached_grant_bits_addr_beat,
  output [1:0] io_htif_uncached_grant_bits_client_xact_id,
  output [2:0] io_htif_uncached_grant_bits_manager_xact_id,
  output  io_htif_uncached_grant_bits_is_builtin_type,
  output [3:0] io_htif_uncached_grant_bits_g_type,
  output [63:0] io_htif_uncached_grant_bits_data,
  input   io_incoherent_0,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_mmio_acquire_ready,
  output  io_mmio_acquire_valid,
  output [25:0] io_mmio_acquire_bits_addr_block,
  output [1:0] io_mmio_acquire_bits_client_xact_id,
  output [2:0] io_mmio_acquire_bits_addr_beat,
  output  io_mmio_acquire_bits_is_builtin_type,
  output [2:0] io_mmio_acquire_bits_a_type,
  output [11:0] io_mmio_acquire_bits_union,
  output [63:0] io_mmio_acquire_bits_data,
  output  io_mmio_grant_ready,
  input   io_mmio_grant_valid,
  input  [2:0] io_mmio_grant_bits_addr_beat,
  input  [1:0] io_mmio_grant_bits_client_xact_id,
  input   io_mmio_grant_bits_manager_xact_id,
  input   io_mmio_grant_bits_is_builtin_type,
  input  [3:0] io_mmio_grant_bits_g_type,
  input  [63:0] io_mmio_grant_bits_data
);
  wire  l1tol2net_clk;
  wire  l1tol2net_reset;
  wire  l1tol2net_io_clients_cached_0_acquire_ready;
  wire  l1tol2net_io_clients_cached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_cached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_cached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_cached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_cached_0_probe_ready;
  wire  l1tol2net_io_clients_cached_0_probe_valid;
  wire [25:0] l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_probe_bits_p_type;
  wire  l1tol2net_io_clients_cached_0_release_ready;
  wire  l1tol2net_io_clients_cached_0_release_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_clients_cached_0_release_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_cached_0_release_bits_client_xact_id;
  wire  l1tol2net_io_clients_cached_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_clients_cached_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_clients_cached_0_release_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_ready;
  wire  l1tol2net_io_clients_cached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_cached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_cached_0_grant_bits_data;
  wire  l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  wire  l1tol2net_io_clients_cached_0_finish_ready;
  wire  l1tol2net_io_clients_cached_0_finish_valid;
  wire [2:0] l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_clients_cached_0_finish_bits_manager_id;
  wire  l1tol2net_io_clients_uncached_0_acquire_ready;
  wire  l1tol2net_io_clients_uncached_0_acquire_valid;
  wire [25:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_uncached_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_uncached_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_uncached_0_acquire_bits_data;
  wire  l1tol2net_io_clients_uncached_0_grant_ready;
  wire  l1tol2net_io_clients_uncached_0_grant_valid;
  wire [2:0] l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_uncached_0_grant_bits_data;
  wire  l1tol2net_io_clients_uncached_1_acquire_ready;
  wire  l1tol2net_io_clients_uncached_1_acquire_valid;
  wire [25:0] l1tol2net_io_clients_uncached_1_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_clients_uncached_1_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_1_acquire_bits_addr_beat;
  wire  l1tol2net_io_clients_uncached_1_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_clients_uncached_1_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_clients_uncached_1_acquire_bits_union;
  wire [63:0] l1tol2net_io_clients_uncached_1_acquire_bits_data;
  wire  l1tol2net_io_clients_uncached_1_grant_ready;
  wire  l1tol2net_io_clients_uncached_1_grant_valid;
  wire [2:0] l1tol2net_io_clients_uncached_1_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_clients_uncached_1_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_clients_uncached_1_grant_bits_manager_xact_id;
  wire  l1tol2net_io_clients_uncached_1_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_clients_uncached_1_grant_bits_g_type;
  wire [63:0] l1tol2net_io_clients_uncached_1_grant_bits_data;
  wire  l1tol2net_io_managers_0_acquire_ready;
  wire  l1tol2net_io_managers_0_acquire_valid;
  wire [25:0] l1tol2net_io_managers_0_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_0_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_0_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_0_acquire_bits_data;
  wire [1:0] l1tol2net_io_managers_0_acquire_bits_client_id;
  wire  l1tol2net_io_managers_0_grant_ready;
  wire  l1tol2net_io_managers_0_grant_valid;
  wire [2:0] l1tol2net_io_managers_0_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_managers_0_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_0_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_0_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_0_grant_bits_data;
  wire [1:0] l1tol2net_io_managers_0_grant_bits_client_id;
  wire  l1tol2net_io_managers_0_finish_ready;
  wire  l1tol2net_io_managers_0_finish_valid;
  wire [2:0] l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_0_probe_ready;
  wire  l1tol2net_io_managers_0_probe_valid;
  wire [25:0] l1tol2net_io_managers_0_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_probe_bits_p_type;
  wire [1:0] l1tol2net_io_managers_0_probe_bits_client_id;
  wire  l1tol2net_io_managers_0_release_ready;
  wire  l1tol2net_io_managers_0_release_valid;
  wire [2:0] l1tol2net_io_managers_0_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_0_release_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_0_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_0_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_0_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_0_release_bits_data;
  wire [1:0] l1tol2net_io_managers_0_release_bits_client_id;
  wire  l1tol2net_io_managers_1_acquire_ready;
  wire  l1tol2net_io_managers_1_acquire_valid;
  wire [25:0] l1tol2net_io_managers_1_acquire_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_addr_beat;
  wire  l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  wire [2:0] l1tol2net_io_managers_1_acquire_bits_a_type;
  wire [11:0] l1tol2net_io_managers_1_acquire_bits_union;
  wire [63:0] l1tol2net_io_managers_1_acquire_bits_data;
  wire [1:0] l1tol2net_io_managers_1_acquire_bits_client_id;
  wire  l1tol2net_io_managers_1_grant_ready;
  wire  l1tol2net_io_managers_1_grant_valid;
  wire [2:0] l1tol2net_io_managers_1_grant_bits_addr_beat;
  wire [1:0] l1tol2net_io_managers_1_grant_bits_client_xact_id;
  wire [2:0] l1tol2net_io_managers_1_grant_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_grant_bits_is_builtin_type;
  wire [3:0] l1tol2net_io_managers_1_grant_bits_g_type;
  wire [63:0] l1tol2net_io_managers_1_grant_bits_data;
  wire [1:0] l1tol2net_io_managers_1_grant_bits_client_id;
  wire  l1tol2net_io_managers_1_finish_ready;
  wire  l1tol2net_io_managers_1_finish_valid;
  wire [2:0] l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  wire  l1tol2net_io_managers_1_probe_ready;
  wire  l1tol2net_io_managers_1_probe_valid;
  wire [25:0] l1tol2net_io_managers_1_probe_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_probe_bits_p_type;
  wire [1:0] l1tol2net_io_managers_1_probe_bits_client_id;
  wire  l1tol2net_io_managers_1_release_ready;
  wire  l1tol2net_io_managers_1_release_valid;
  wire [2:0] l1tol2net_io_managers_1_release_bits_addr_beat;
  wire [25:0] l1tol2net_io_managers_1_release_bits_addr_block;
  wire [1:0] l1tol2net_io_managers_1_release_bits_client_xact_id;
  wire  l1tol2net_io_managers_1_release_bits_voluntary;
  wire [2:0] l1tol2net_io_managers_1_release_bits_r_type;
  wire [63:0] l1tol2net_io_managers_1_release_bits_data;
  wire [1:0] l1tol2net_io_managers_1_release_bits_client_id;
  wire  L2BroadcastHub_8569_clk;
  wire  L2BroadcastHub_8569_reset;
  wire  L2BroadcastHub_8569_io_inner_acquire_ready;
  wire  L2BroadcastHub_8569_io_inner_acquire_valid;
  wire [25:0] L2BroadcastHub_8569_io_inner_acquire_bits_addr_block;
  wire [1:0] L2BroadcastHub_8569_io_inner_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_8569_io_inner_acquire_bits_addr_beat;
  wire  L2BroadcastHub_8569_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_8569_io_inner_acquire_bits_a_type;
  wire [11:0] L2BroadcastHub_8569_io_inner_acquire_bits_union;
  wire [63:0] L2BroadcastHub_8569_io_inner_acquire_bits_data;
  wire [1:0] L2BroadcastHub_8569_io_inner_acquire_bits_client_id;
  wire  L2BroadcastHub_8569_io_inner_grant_ready;
  wire  L2BroadcastHub_8569_io_inner_grant_valid;
  wire [2:0] L2BroadcastHub_8569_io_inner_grant_bits_addr_beat;
  wire [1:0] L2BroadcastHub_8569_io_inner_grant_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_8569_io_inner_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_8569_io_inner_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_8569_io_inner_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_8569_io_inner_grant_bits_data;
  wire [1:0] L2BroadcastHub_8569_io_inner_grant_bits_client_id;
  wire  L2BroadcastHub_8569_io_inner_finish_ready;
  wire  L2BroadcastHub_8569_io_inner_finish_valid;
  wire [2:0] L2BroadcastHub_8569_io_inner_finish_bits_manager_xact_id;
  wire  L2BroadcastHub_8569_io_inner_probe_ready;
  wire  L2BroadcastHub_8569_io_inner_probe_valid;
  wire [25:0] L2BroadcastHub_8569_io_inner_probe_bits_addr_block;
  wire [1:0] L2BroadcastHub_8569_io_inner_probe_bits_p_type;
  wire [1:0] L2BroadcastHub_8569_io_inner_probe_bits_client_id;
  wire  L2BroadcastHub_8569_io_inner_release_ready;
  wire  L2BroadcastHub_8569_io_inner_release_valid;
  wire [2:0] L2BroadcastHub_8569_io_inner_release_bits_addr_beat;
  wire [25:0] L2BroadcastHub_8569_io_inner_release_bits_addr_block;
  wire [1:0] L2BroadcastHub_8569_io_inner_release_bits_client_xact_id;
  wire  L2BroadcastHub_8569_io_inner_release_bits_voluntary;
  wire [2:0] L2BroadcastHub_8569_io_inner_release_bits_r_type;
  wire [63:0] L2BroadcastHub_8569_io_inner_release_bits_data;
  wire [1:0] L2BroadcastHub_8569_io_inner_release_bits_client_id;
  wire  L2BroadcastHub_8569_io_incoherent_0;
  wire  L2BroadcastHub_8569_io_outer_acquire_ready;
  wire  L2BroadcastHub_8569_io_outer_acquire_valid;
  wire [25:0] L2BroadcastHub_8569_io_outer_acquire_bits_addr_block;
  wire [2:0] L2BroadcastHub_8569_io_outer_acquire_bits_client_xact_id;
  wire [2:0] L2BroadcastHub_8569_io_outer_acquire_bits_addr_beat;
  wire  L2BroadcastHub_8569_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] L2BroadcastHub_8569_io_outer_acquire_bits_a_type;
  wire [11:0] L2BroadcastHub_8569_io_outer_acquire_bits_union;
  wire [63:0] L2BroadcastHub_8569_io_outer_acquire_bits_data;
  wire  L2BroadcastHub_8569_io_outer_grant_ready;
  wire  L2BroadcastHub_8569_io_outer_grant_valid;
  wire [2:0] L2BroadcastHub_8569_io_outer_grant_bits_addr_beat;
  wire [2:0] L2BroadcastHub_8569_io_outer_grant_bits_client_xact_id;
  wire  L2BroadcastHub_8569_io_outer_grant_bits_manager_xact_id;
  wire  L2BroadcastHub_8569_io_outer_grant_bits_is_builtin_type;
  wire [3:0] L2BroadcastHub_8569_io_outer_grant_bits_g_type;
  wire [63:0] L2BroadcastHub_8569_io_outer_grant_bits_data;
  wire  mmioManager_clk;
  wire  mmioManager_reset;
  wire  mmioManager_io_inner_acquire_ready;
  wire  mmioManager_io_inner_acquire_valid;
  wire [25:0] mmioManager_io_inner_acquire_bits_addr_block;
  wire [1:0] mmioManager_io_inner_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_inner_acquire_bits_addr_beat;
  wire  mmioManager_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_inner_acquire_bits_a_type;
  wire [11:0] mmioManager_io_inner_acquire_bits_union;
  wire [63:0] mmioManager_io_inner_acquire_bits_data;
  wire [1:0] mmioManager_io_inner_acquire_bits_client_id;
  wire  mmioManager_io_inner_grant_ready;
  wire  mmioManager_io_inner_grant_valid;
  wire [2:0] mmioManager_io_inner_grant_bits_addr_beat;
  wire [1:0] mmioManager_io_inner_grant_bits_client_xact_id;
  wire [2:0] mmioManager_io_inner_grant_bits_manager_xact_id;
  wire  mmioManager_io_inner_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_inner_grant_bits_g_type;
  wire [63:0] mmioManager_io_inner_grant_bits_data;
  wire [1:0] mmioManager_io_inner_grant_bits_client_id;
  wire  mmioManager_io_inner_finish_ready;
  wire  mmioManager_io_inner_finish_valid;
  wire [2:0] mmioManager_io_inner_finish_bits_manager_xact_id;
  wire  mmioManager_io_inner_probe_ready;
  wire  mmioManager_io_inner_probe_valid;
  wire [25:0] mmioManager_io_inner_probe_bits_addr_block;
  wire [1:0] mmioManager_io_inner_probe_bits_p_type;
  wire [1:0] mmioManager_io_inner_probe_bits_client_id;
  wire  mmioManager_io_inner_release_ready;
  wire  mmioManager_io_inner_release_valid;
  wire [2:0] mmioManager_io_inner_release_bits_addr_beat;
  wire [25:0] mmioManager_io_inner_release_bits_addr_block;
  wire [1:0] mmioManager_io_inner_release_bits_client_xact_id;
  wire  mmioManager_io_inner_release_bits_voluntary;
  wire [2:0] mmioManager_io_inner_release_bits_r_type;
  wire [63:0] mmioManager_io_inner_release_bits_data;
  wire [1:0] mmioManager_io_inner_release_bits_client_id;
  wire  mmioManager_io_incoherent_0;
  wire  mmioManager_io_outer_acquire_ready;
  wire  mmioManager_io_outer_acquire_valid;
  wire [25:0] mmioManager_io_outer_acquire_bits_addr_block;
  wire [1:0] mmioManager_io_outer_acquire_bits_client_xact_id;
  wire [2:0] mmioManager_io_outer_acquire_bits_addr_beat;
  wire  mmioManager_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] mmioManager_io_outer_acquire_bits_a_type;
  wire [11:0] mmioManager_io_outer_acquire_bits_union;
  wire [63:0] mmioManager_io_outer_acquire_bits_data;
  wire  mmioManager_io_outer_grant_ready;
  wire  mmioManager_io_outer_grant_valid;
  wire [2:0] mmioManager_io_outer_grant_bits_addr_beat;
  wire [1:0] mmioManager_io_outer_grant_bits_client_xact_id;
  wire  mmioManager_io_outer_grant_bits_manager_xact_id;
  wire  mmioManager_io_outer_grant_bits_is_builtin_type;
  wire [3:0] mmioManager_io_outer_grant_bits_g_type;
  wire [63:0] mmioManager_io_outer_grant_bits_data;
  wire  mem_ic_clk;
  wire  mem_ic_reset;
  wire  mem_ic_io_in_0_acquire_ready;
  wire  mem_ic_io_in_0_acquire_valid;
  wire [25:0] mem_ic_io_in_0_acquire_bits_addr_block;
  wire [2:0] mem_ic_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_in_0_acquire_bits_addr_beat;
  wire  mem_ic_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_in_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_in_0_acquire_bits_union;
  wire [63:0] mem_ic_io_in_0_acquire_bits_data;
  wire  mem_ic_io_in_0_grant_ready;
  wire  mem_ic_io_in_0_grant_valid;
  wire [2:0] mem_ic_io_in_0_grant_bits_addr_beat;
  wire [2:0] mem_ic_io_in_0_grant_bits_client_xact_id;
  wire  mem_ic_io_in_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_in_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_in_0_grant_bits_data;
  wire  mem_ic_io_out_0_acquire_ready;
  wire  mem_ic_io_out_0_acquire_valid;
  wire [25:0] mem_ic_io_out_0_acquire_bits_addr_block;
  wire [2:0] mem_ic_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] mem_ic_io_out_0_acquire_bits_addr_beat;
  wire  mem_ic_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] mem_ic_io_out_0_acquire_bits_a_type;
  wire [11:0] mem_ic_io_out_0_acquire_bits_union;
  wire [63:0] mem_ic_io_out_0_acquire_bits_data;
  wire  mem_ic_io_out_0_grant_ready;
  wire  mem_ic_io_out_0_grant_valid;
  wire [2:0] mem_ic_io_out_0_grant_bits_addr_beat;
  wire [2:0] mem_ic_io_out_0_grant_bits_client_xact_id;
  wire  mem_ic_io_out_0_grant_bits_manager_xact_id;
  wire  mem_ic_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] mem_ic_io_out_0_grant_bits_g_type;
  wire [63:0] mem_ic_io_out_0_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_8570_clk;
  wire  ClientTileLinkIOUnwrapper_8570_reset;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_probe_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_probe_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_p_type;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_release_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_release_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_release_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_release_bits_r_type;
  wire [63:0] ClientTileLinkIOUnwrapper_8570_io_in_release_bits_data;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_grant_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_data;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_finish_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_finish_valid;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_acquire_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_data;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_grant_ready;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_data;
  wire  ClientTileLinkIOWrapper_8571_clk;
  wire  ClientTileLinkIOWrapper_8571_reset;
  wire  ClientTileLinkIOWrapper_8571_io_in_acquire_ready;
  wire  ClientTileLinkIOWrapper_8571_io_in_acquire_valid;
  wire [25:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_beat;
  wire  ClientTileLinkIOWrapper_8571_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_union;
  wire [63:0] ClientTileLinkIOWrapper_8571_io_in_acquire_bits_data;
  wire  ClientTileLinkIOWrapper_8571_io_in_grant_ready;
  wire  ClientTileLinkIOWrapper_8571_io_in_grant_valid;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_in_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_in_grant_bits_client_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_in_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOWrapper_8571_io_in_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOWrapper_8571_io_in_grant_bits_data;
  wire  ClientTileLinkIOWrapper_8571_io_out_acquire_ready;
  wire  ClientTileLinkIOWrapper_8571_io_out_acquire_valid;
  wire [25:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_beat;
  wire  ClientTileLinkIOWrapper_8571_io_out_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_a_type;
  wire [11:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_union;
  wire [63:0] ClientTileLinkIOWrapper_8571_io_out_acquire_bits_data;
  wire  ClientTileLinkIOWrapper_8571_io_out_probe_ready;
  wire  ClientTileLinkIOWrapper_8571_io_out_probe_valid;
  wire [25:0] ClientTileLinkIOWrapper_8571_io_out_probe_bits_addr_block;
  wire [1:0] ClientTileLinkIOWrapper_8571_io_out_probe_bits_p_type;
  wire  ClientTileLinkIOWrapper_8571_io_out_release_ready;
  wire  ClientTileLinkIOWrapper_8571_io_out_release_valid;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_beat;
  wire [25:0] ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_block;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_release_bits_client_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_out_release_bits_voluntary;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_release_bits_r_type;
  wire [63:0] ClientTileLinkIOWrapper_8571_io_out_release_bits_data;
  wire  ClientTileLinkIOWrapper_8571_io_out_grant_ready;
  wire  ClientTileLinkIOWrapper_8571_io_out_grant_valid;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkIOWrapper_8571_io_out_grant_bits_client_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_out_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkIOWrapper_8571_io_out_grant_bits_g_type;
  wire [63:0] ClientTileLinkIOWrapper_8571_io_out_grant_bits_data;
  wire  ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_id;
  wire  ClientTileLinkIOWrapper_8571_io_out_finish_ready;
  wire  ClientTileLinkIOWrapper_8571_io_out_finish_valid;
  wire  ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_xact_id;
  wire  ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_8572_clk;
  wire  ClientTileLinkEnqueuer_8572_reset;
  wire  ClientTileLinkEnqueuer_8572_io_inner_acquire_ready;
  wire  ClientTileLinkEnqueuer_8572_io_inner_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_inner_probe_ready;
  wire  ClientTileLinkEnqueuer_8572_io_inner_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_inner_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_8572_io_inner_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_8572_io_inner_release_ready;
  wire  ClientTileLinkEnqueuer_8572_io_inner_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_inner_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_inner_release_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_inner_grant_ready;
  wire  ClientTileLinkEnqueuer_8572_io_inner_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_inner_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_inner_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_8572_io_inner_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_inner_grant_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_8572_io_inner_finish_ready;
  wire  ClientTileLinkEnqueuer_8572_io_inner_finish_valid;
  wire  ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_acquire_ready;
  wire  ClientTileLinkEnqueuer_8572_io_outer_acquire_valid;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_client_xact_id;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_beat;
  wire  ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_is_builtin_type;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_a_type;
  wire [11:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_union;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_outer_probe_ready;
  wire  ClientTileLinkEnqueuer_8572_io_outer_probe_valid;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_outer_probe_bits_addr_block;
  wire [1:0] ClientTileLinkEnqueuer_8572_io_outer_probe_bits_p_type;
  wire  ClientTileLinkEnqueuer_8572_io_outer_release_ready;
  wire  ClientTileLinkEnqueuer_8572_io_outer_release_valid;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_beat;
  wire [25:0] ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_block;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_release_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_release_bits_voluntary;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_release_bits_r_type;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_outer_release_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_outer_grant_ready;
  wire  ClientTileLinkEnqueuer_8572_io_outer_grant_valid;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_grant_bits_addr_beat;
  wire [2:0] ClientTileLinkEnqueuer_8572_io_outer_grant_bits_client_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_grant_bits_is_builtin_type;
  wire [3:0] ClientTileLinkEnqueuer_8572_io_outer_grant_bits_g_type;
  wire [63:0] ClientTileLinkEnqueuer_8572_io_outer_grant_bits_data;
  wire  ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_finish_ready;
  wire  ClientTileLinkEnqueuer_8572_io_outer_finish_valid;
  wire  ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_xact_id;
  wire  ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_id;
  wire  NastiIOTileLinkIOConverter_8573_clk;
  wire  NastiIOTileLinkIOConverter_8573_reset;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_block;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_addr_beat;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_user;
  wire  Queue_39_8586_clk;
  wire  Queue_39_8586_reset;
  wire  Queue_39_8586_io_enq_ready;
  wire  Queue_39_8586_io_enq_valid;
  wire [31:0] Queue_39_8586_io_enq_bits_addr;
  wire [7:0] Queue_39_8586_io_enq_bits_len;
  wire [2:0] Queue_39_8586_io_enq_bits_size;
  wire [1:0] Queue_39_8586_io_enq_bits_burst;
  wire  Queue_39_8586_io_enq_bits_lock;
  wire [3:0] Queue_39_8586_io_enq_bits_cache;
  wire [2:0] Queue_39_8586_io_enq_bits_prot;
  wire [3:0] Queue_39_8586_io_enq_bits_qos;
  wire [3:0] Queue_39_8586_io_enq_bits_region;
  wire [4:0] Queue_39_8586_io_enq_bits_id;
  wire  Queue_39_8586_io_enq_bits_user;
  wire  Queue_39_8586_io_deq_ready;
  wire  Queue_39_8586_io_deq_valid;
  wire [31:0] Queue_39_8586_io_deq_bits_addr;
  wire [7:0] Queue_39_8586_io_deq_bits_len;
  wire [2:0] Queue_39_8586_io_deq_bits_size;
  wire [1:0] Queue_39_8586_io_deq_bits_burst;
  wire  Queue_39_8586_io_deq_bits_lock;
  wire [3:0] Queue_39_8586_io_deq_bits_cache;
  wire [2:0] Queue_39_8586_io_deq_bits_prot;
  wire [3:0] Queue_39_8586_io_deq_bits_qos;
  wire [3:0] Queue_39_8586_io_deq_bits_region;
  wire [4:0] Queue_39_8586_io_deq_bits_id;
  wire  Queue_39_8586_io_deq_bits_user;
  wire  Queue_39_8586_io_count;
  wire  Queue_40_8599_clk;
  wire  Queue_40_8599_reset;
  wire  Queue_40_8599_io_enq_ready;
  wire  Queue_40_8599_io_enq_valid;
  wire [31:0] Queue_40_8599_io_enq_bits_addr;
  wire [7:0] Queue_40_8599_io_enq_bits_len;
  wire [2:0] Queue_40_8599_io_enq_bits_size;
  wire [1:0] Queue_40_8599_io_enq_bits_burst;
  wire  Queue_40_8599_io_enq_bits_lock;
  wire [3:0] Queue_40_8599_io_enq_bits_cache;
  wire [2:0] Queue_40_8599_io_enq_bits_prot;
  wire [3:0] Queue_40_8599_io_enq_bits_qos;
  wire [3:0] Queue_40_8599_io_enq_bits_region;
  wire [4:0] Queue_40_8599_io_enq_bits_id;
  wire  Queue_40_8599_io_enq_bits_user;
  wire  Queue_40_8599_io_deq_ready;
  wire  Queue_40_8599_io_deq_valid;
  wire [31:0] Queue_40_8599_io_deq_bits_addr;
  wire [7:0] Queue_40_8599_io_deq_bits_len;
  wire [2:0] Queue_40_8599_io_deq_bits_size;
  wire [1:0] Queue_40_8599_io_deq_bits_burst;
  wire  Queue_40_8599_io_deq_bits_lock;
  wire [3:0] Queue_40_8599_io_deq_bits_cache;
  wire [2:0] Queue_40_8599_io_deq_bits_prot;
  wire [3:0] Queue_40_8599_io_deq_bits_qos;
  wire [3:0] Queue_40_8599_io_deq_bits_region;
  wire [4:0] Queue_40_8599_io_deq_bits_id;
  wire  Queue_40_8599_io_deq_bits_user;
  wire  Queue_40_8599_io_count;
  wire  Queue_41_8606_clk;
  wire  Queue_41_8606_reset;
  wire  Queue_41_8606_io_enq_ready;
  wire  Queue_41_8606_io_enq_valid;
  wire [63:0] Queue_41_8606_io_enq_bits_data;
  wire  Queue_41_8606_io_enq_bits_last;
  wire [4:0] Queue_41_8606_io_enq_bits_id;
  wire [7:0] Queue_41_8606_io_enq_bits_strb;
  wire  Queue_41_8606_io_enq_bits_user;
  wire  Queue_41_8606_io_deq_ready;
  wire  Queue_41_8606_io_deq_valid;
  wire [63:0] Queue_41_8606_io_deq_bits_data;
  wire  Queue_41_8606_io_deq_bits_last;
  wire [4:0] Queue_41_8606_io_deq_bits_id;
  wire [7:0] Queue_41_8606_io_deq_bits_strb;
  wire  Queue_41_8606_io_deq_bits_user;
  wire [1:0] Queue_41_8606_io_count;
  wire  Queue_42_8613_clk;
  wire  Queue_42_8613_reset;
  wire  Queue_42_8613_io_enq_ready;
  wire  Queue_42_8613_io_enq_valid;
  wire [1:0] Queue_42_8613_io_enq_bits_resp;
  wire [63:0] Queue_42_8613_io_enq_bits_data;
  wire  Queue_42_8613_io_enq_bits_last;
  wire [4:0] Queue_42_8613_io_enq_bits_id;
  wire  Queue_42_8613_io_enq_bits_user;
  wire  Queue_42_8613_io_deq_ready;
  wire  Queue_42_8613_io_deq_valid;
  wire [1:0] Queue_42_8613_io_deq_bits_resp;
  wire [63:0] Queue_42_8613_io_deq_bits_data;
  wire  Queue_42_8613_io_deq_bits_last;
  wire [4:0] Queue_42_8613_io_deq_bits_id;
  wire  Queue_42_8613_io_deq_bits_user;
  wire [1:0] Queue_42_8613_io_count;
  wire  Queue_43_8618_clk;
  wire  Queue_43_8618_reset;
  wire  Queue_43_8618_io_enq_ready;
  wire  Queue_43_8618_io_enq_valid;
  wire [1:0] Queue_43_8618_io_enq_bits_resp;
  wire [4:0] Queue_43_8618_io_enq_bits_id;
  wire  Queue_43_8618_io_enq_bits_user;
  wire  Queue_43_8618_io_deq_ready;
  wire  Queue_43_8618_io_deq_valid;
  wire [1:0] Queue_43_8618_io_deq_bits_resp;
  wire [4:0] Queue_43_8618_io_deq_bits_id;
  wire  Queue_43_8618_io_deq_bits_user;
  wire  Queue_43_8618_io_count;
  reg  GEN_0;
  reg [31:0] GEN_1;
  PortedTileLinkCrossbar l1tol2net (
    .clk(l1tol2net_clk),
    .reset(l1tol2net_reset),
    .io_clients_cached_0_acquire_ready(l1tol2net_io_clients_cached_0_acquire_ready),
    .io_clients_cached_0_acquire_valid(l1tol2net_io_clients_cached_0_acquire_valid),
    .io_clients_cached_0_acquire_bits_addr_block(l1tol2net_io_clients_cached_0_acquire_bits_addr_block),
    .io_clients_cached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id),
    .io_clients_cached_0_acquire_bits_addr_beat(l1tol2net_io_clients_cached_0_acquire_bits_addr_beat),
    .io_clients_cached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type),
    .io_clients_cached_0_acquire_bits_a_type(l1tol2net_io_clients_cached_0_acquire_bits_a_type),
    .io_clients_cached_0_acquire_bits_union(l1tol2net_io_clients_cached_0_acquire_bits_union),
    .io_clients_cached_0_acquire_bits_data(l1tol2net_io_clients_cached_0_acquire_bits_data),
    .io_clients_cached_0_probe_ready(l1tol2net_io_clients_cached_0_probe_ready),
    .io_clients_cached_0_probe_valid(l1tol2net_io_clients_cached_0_probe_valid),
    .io_clients_cached_0_probe_bits_addr_block(l1tol2net_io_clients_cached_0_probe_bits_addr_block),
    .io_clients_cached_0_probe_bits_p_type(l1tol2net_io_clients_cached_0_probe_bits_p_type),
    .io_clients_cached_0_release_ready(l1tol2net_io_clients_cached_0_release_ready),
    .io_clients_cached_0_release_valid(l1tol2net_io_clients_cached_0_release_valid),
    .io_clients_cached_0_release_bits_addr_beat(l1tol2net_io_clients_cached_0_release_bits_addr_beat),
    .io_clients_cached_0_release_bits_addr_block(l1tol2net_io_clients_cached_0_release_bits_addr_block),
    .io_clients_cached_0_release_bits_client_xact_id(l1tol2net_io_clients_cached_0_release_bits_client_xact_id),
    .io_clients_cached_0_release_bits_voluntary(l1tol2net_io_clients_cached_0_release_bits_voluntary),
    .io_clients_cached_0_release_bits_r_type(l1tol2net_io_clients_cached_0_release_bits_r_type),
    .io_clients_cached_0_release_bits_data(l1tol2net_io_clients_cached_0_release_bits_data),
    .io_clients_cached_0_grant_ready(l1tol2net_io_clients_cached_0_grant_ready),
    .io_clients_cached_0_grant_valid(l1tol2net_io_clients_cached_0_grant_valid),
    .io_clients_cached_0_grant_bits_addr_beat(l1tol2net_io_clients_cached_0_grant_bits_addr_beat),
    .io_clients_cached_0_grant_bits_client_xact_id(l1tol2net_io_clients_cached_0_grant_bits_client_xact_id),
    .io_clients_cached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id),
    .io_clients_cached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type),
    .io_clients_cached_0_grant_bits_g_type(l1tol2net_io_clients_cached_0_grant_bits_g_type),
    .io_clients_cached_0_grant_bits_data(l1tol2net_io_clients_cached_0_grant_bits_data),
    .io_clients_cached_0_grant_bits_manager_id(l1tol2net_io_clients_cached_0_grant_bits_manager_id),
    .io_clients_cached_0_finish_ready(l1tol2net_io_clients_cached_0_finish_ready),
    .io_clients_cached_0_finish_valid(l1tol2net_io_clients_cached_0_finish_valid),
    .io_clients_cached_0_finish_bits_manager_xact_id(l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id),
    .io_clients_cached_0_finish_bits_manager_id(l1tol2net_io_clients_cached_0_finish_bits_manager_id),
    .io_clients_uncached_0_acquire_ready(l1tol2net_io_clients_uncached_0_acquire_ready),
    .io_clients_uncached_0_acquire_valid(l1tol2net_io_clients_uncached_0_acquire_valid),
    .io_clients_uncached_0_acquire_bits_addr_block(l1tol2net_io_clients_uncached_0_acquire_bits_addr_block),
    .io_clients_uncached_0_acquire_bits_client_xact_id(l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id),
    .io_clients_uncached_0_acquire_bits_addr_beat(l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat),
    .io_clients_uncached_0_acquire_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type),
    .io_clients_uncached_0_acquire_bits_a_type(l1tol2net_io_clients_uncached_0_acquire_bits_a_type),
    .io_clients_uncached_0_acquire_bits_union(l1tol2net_io_clients_uncached_0_acquire_bits_union),
    .io_clients_uncached_0_acquire_bits_data(l1tol2net_io_clients_uncached_0_acquire_bits_data),
    .io_clients_uncached_0_grant_ready(l1tol2net_io_clients_uncached_0_grant_ready),
    .io_clients_uncached_0_grant_valid(l1tol2net_io_clients_uncached_0_grant_valid),
    .io_clients_uncached_0_grant_bits_addr_beat(l1tol2net_io_clients_uncached_0_grant_bits_addr_beat),
    .io_clients_uncached_0_grant_bits_client_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id),
    .io_clients_uncached_0_grant_bits_manager_xact_id(l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id),
    .io_clients_uncached_0_grant_bits_is_builtin_type(l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type),
    .io_clients_uncached_0_grant_bits_g_type(l1tol2net_io_clients_uncached_0_grant_bits_g_type),
    .io_clients_uncached_0_grant_bits_data(l1tol2net_io_clients_uncached_0_grant_bits_data),
    .io_clients_uncached_1_acquire_ready(l1tol2net_io_clients_uncached_1_acquire_ready),
    .io_clients_uncached_1_acquire_valid(l1tol2net_io_clients_uncached_1_acquire_valid),
    .io_clients_uncached_1_acquire_bits_addr_block(l1tol2net_io_clients_uncached_1_acquire_bits_addr_block),
    .io_clients_uncached_1_acquire_bits_client_xact_id(l1tol2net_io_clients_uncached_1_acquire_bits_client_xact_id),
    .io_clients_uncached_1_acquire_bits_addr_beat(l1tol2net_io_clients_uncached_1_acquire_bits_addr_beat),
    .io_clients_uncached_1_acquire_bits_is_builtin_type(l1tol2net_io_clients_uncached_1_acquire_bits_is_builtin_type),
    .io_clients_uncached_1_acquire_bits_a_type(l1tol2net_io_clients_uncached_1_acquire_bits_a_type),
    .io_clients_uncached_1_acquire_bits_union(l1tol2net_io_clients_uncached_1_acquire_bits_union),
    .io_clients_uncached_1_acquire_bits_data(l1tol2net_io_clients_uncached_1_acquire_bits_data),
    .io_clients_uncached_1_grant_ready(l1tol2net_io_clients_uncached_1_grant_ready),
    .io_clients_uncached_1_grant_valid(l1tol2net_io_clients_uncached_1_grant_valid),
    .io_clients_uncached_1_grant_bits_addr_beat(l1tol2net_io_clients_uncached_1_grant_bits_addr_beat),
    .io_clients_uncached_1_grant_bits_client_xact_id(l1tol2net_io_clients_uncached_1_grant_bits_client_xact_id),
    .io_clients_uncached_1_grant_bits_manager_xact_id(l1tol2net_io_clients_uncached_1_grant_bits_manager_xact_id),
    .io_clients_uncached_1_grant_bits_is_builtin_type(l1tol2net_io_clients_uncached_1_grant_bits_is_builtin_type),
    .io_clients_uncached_1_grant_bits_g_type(l1tol2net_io_clients_uncached_1_grant_bits_g_type),
    .io_clients_uncached_1_grant_bits_data(l1tol2net_io_clients_uncached_1_grant_bits_data),
    .io_managers_0_acquire_ready(l1tol2net_io_managers_0_acquire_ready),
    .io_managers_0_acquire_valid(l1tol2net_io_managers_0_acquire_valid),
    .io_managers_0_acquire_bits_addr_block(l1tol2net_io_managers_0_acquire_bits_addr_block),
    .io_managers_0_acquire_bits_client_xact_id(l1tol2net_io_managers_0_acquire_bits_client_xact_id),
    .io_managers_0_acquire_bits_addr_beat(l1tol2net_io_managers_0_acquire_bits_addr_beat),
    .io_managers_0_acquire_bits_is_builtin_type(l1tol2net_io_managers_0_acquire_bits_is_builtin_type),
    .io_managers_0_acquire_bits_a_type(l1tol2net_io_managers_0_acquire_bits_a_type),
    .io_managers_0_acquire_bits_union(l1tol2net_io_managers_0_acquire_bits_union),
    .io_managers_0_acquire_bits_data(l1tol2net_io_managers_0_acquire_bits_data),
    .io_managers_0_acquire_bits_client_id(l1tol2net_io_managers_0_acquire_bits_client_id),
    .io_managers_0_grant_ready(l1tol2net_io_managers_0_grant_ready),
    .io_managers_0_grant_valid(l1tol2net_io_managers_0_grant_valid),
    .io_managers_0_grant_bits_addr_beat(l1tol2net_io_managers_0_grant_bits_addr_beat),
    .io_managers_0_grant_bits_client_xact_id(l1tol2net_io_managers_0_grant_bits_client_xact_id),
    .io_managers_0_grant_bits_manager_xact_id(l1tol2net_io_managers_0_grant_bits_manager_xact_id),
    .io_managers_0_grant_bits_is_builtin_type(l1tol2net_io_managers_0_grant_bits_is_builtin_type),
    .io_managers_0_grant_bits_g_type(l1tol2net_io_managers_0_grant_bits_g_type),
    .io_managers_0_grant_bits_data(l1tol2net_io_managers_0_grant_bits_data),
    .io_managers_0_grant_bits_client_id(l1tol2net_io_managers_0_grant_bits_client_id),
    .io_managers_0_finish_ready(l1tol2net_io_managers_0_finish_ready),
    .io_managers_0_finish_valid(l1tol2net_io_managers_0_finish_valid),
    .io_managers_0_finish_bits_manager_xact_id(l1tol2net_io_managers_0_finish_bits_manager_xact_id),
    .io_managers_0_probe_ready(l1tol2net_io_managers_0_probe_ready),
    .io_managers_0_probe_valid(l1tol2net_io_managers_0_probe_valid),
    .io_managers_0_probe_bits_addr_block(l1tol2net_io_managers_0_probe_bits_addr_block),
    .io_managers_0_probe_bits_p_type(l1tol2net_io_managers_0_probe_bits_p_type),
    .io_managers_0_probe_bits_client_id(l1tol2net_io_managers_0_probe_bits_client_id),
    .io_managers_0_release_ready(l1tol2net_io_managers_0_release_ready),
    .io_managers_0_release_valid(l1tol2net_io_managers_0_release_valid),
    .io_managers_0_release_bits_addr_beat(l1tol2net_io_managers_0_release_bits_addr_beat),
    .io_managers_0_release_bits_addr_block(l1tol2net_io_managers_0_release_bits_addr_block),
    .io_managers_0_release_bits_client_xact_id(l1tol2net_io_managers_0_release_bits_client_xact_id),
    .io_managers_0_release_bits_voluntary(l1tol2net_io_managers_0_release_bits_voluntary),
    .io_managers_0_release_bits_r_type(l1tol2net_io_managers_0_release_bits_r_type),
    .io_managers_0_release_bits_data(l1tol2net_io_managers_0_release_bits_data),
    .io_managers_0_release_bits_client_id(l1tol2net_io_managers_0_release_bits_client_id),
    .io_managers_1_acquire_ready(l1tol2net_io_managers_1_acquire_ready),
    .io_managers_1_acquire_valid(l1tol2net_io_managers_1_acquire_valid),
    .io_managers_1_acquire_bits_addr_block(l1tol2net_io_managers_1_acquire_bits_addr_block),
    .io_managers_1_acquire_bits_client_xact_id(l1tol2net_io_managers_1_acquire_bits_client_xact_id),
    .io_managers_1_acquire_bits_addr_beat(l1tol2net_io_managers_1_acquire_bits_addr_beat),
    .io_managers_1_acquire_bits_is_builtin_type(l1tol2net_io_managers_1_acquire_bits_is_builtin_type),
    .io_managers_1_acquire_bits_a_type(l1tol2net_io_managers_1_acquire_bits_a_type),
    .io_managers_1_acquire_bits_union(l1tol2net_io_managers_1_acquire_bits_union),
    .io_managers_1_acquire_bits_data(l1tol2net_io_managers_1_acquire_bits_data),
    .io_managers_1_acquire_bits_client_id(l1tol2net_io_managers_1_acquire_bits_client_id),
    .io_managers_1_grant_ready(l1tol2net_io_managers_1_grant_ready),
    .io_managers_1_grant_valid(l1tol2net_io_managers_1_grant_valid),
    .io_managers_1_grant_bits_addr_beat(l1tol2net_io_managers_1_grant_bits_addr_beat),
    .io_managers_1_grant_bits_client_xact_id(l1tol2net_io_managers_1_grant_bits_client_xact_id),
    .io_managers_1_grant_bits_manager_xact_id(l1tol2net_io_managers_1_grant_bits_manager_xact_id),
    .io_managers_1_grant_bits_is_builtin_type(l1tol2net_io_managers_1_grant_bits_is_builtin_type),
    .io_managers_1_grant_bits_g_type(l1tol2net_io_managers_1_grant_bits_g_type),
    .io_managers_1_grant_bits_data(l1tol2net_io_managers_1_grant_bits_data),
    .io_managers_1_grant_bits_client_id(l1tol2net_io_managers_1_grant_bits_client_id),
    .io_managers_1_finish_ready(l1tol2net_io_managers_1_finish_ready),
    .io_managers_1_finish_valid(l1tol2net_io_managers_1_finish_valid),
    .io_managers_1_finish_bits_manager_xact_id(l1tol2net_io_managers_1_finish_bits_manager_xact_id),
    .io_managers_1_probe_ready(l1tol2net_io_managers_1_probe_ready),
    .io_managers_1_probe_valid(l1tol2net_io_managers_1_probe_valid),
    .io_managers_1_probe_bits_addr_block(l1tol2net_io_managers_1_probe_bits_addr_block),
    .io_managers_1_probe_bits_p_type(l1tol2net_io_managers_1_probe_bits_p_type),
    .io_managers_1_probe_bits_client_id(l1tol2net_io_managers_1_probe_bits_client_id),
    .io_managers_1_release_ready(l1tol2net_io_managers_1_release_ready),
    .io_managers_1_release_valid(l1tol2net_io_managers_1_release_valid),
    .io_managers_1_release_bits_addr_beat(l1tol2net_io_managers_1_release_bits_addr_beat),
    .io_managers_1_release_bits_addr_block(l1tol2net_io_managers_1_release_bits_addr_block),
    .io_managers_1_release_bits_client_xact_id(l1tol2net_io_managers_1_release_bits_client_xact_id),
    .io_managers_1_release_bits_voluntary(l1tol2net_io_managers_1_release_bits_voluntary),
    .io_managers_1_release_bits_r_type(l1tol2net_io_managers_1_release_bits_r_type),
    .io_managers_1_release_bits_data(l1tol2net_io_managers_1_release_bits_data),
    .io_managers_1_release_bits_client_id(l1tol2net_io_managers_1_release_bits_client_id)
  );
  L2BroadcastHub L2BroadcastHub_8569 (
    .clk(L2BroadcastHub_8569_clk),
    .reset(L2BroadcastHub_8569_reset),
    .io_inner_acquire_ready(L2BroadcastHub_8569_io_inner_acquire_ready),
    .io_inner_acquire_valid(L2BroadcastHub_8569_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(L2BroadcastHub_8569_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(L2BroadcastHub_8569_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(L2BroadcastHub_8569_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(L2BroadcastHub_8569_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(L2BroadcastHub_8569_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(L2BroadcastHub_8569_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(L2BroadcastHub_8569_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(L2BroadcastHub_8569_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(L2BroadcastHub_8569_io_inner_grant_ready),
    .io_inner_grant_valid(L2BroadcastHub_8569_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(L2BroadcastHub_8569_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(L2BroadcastHub_8569_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(L2BroadcastHub_8569_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(L2BroadcastHub_8569_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(L2BroadcastHub_8569_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(L2BroadcastHub_8569_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(L2BroadcastHub_8569_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(L2BroadcastHub_8569_io_inner_finish_ready),
    .io_inner_finish_valid(L2BroadcastHub_8569_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(L2BroadcastHub_8569_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(L2BroadcastHub_8569_io_inner_probe_ready),
    .io_inner_probe_valid(L2BroadcastHub_8569_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(L2BroadcastHub_8569_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(L2BroadcastHub_8569_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(L2BroadcastHub_8569_io_inner_probe_bits_client_id),
    .io_inner_release_ready(L2BroadcastHub_8569_io_inner_release_ready),
    .io_inner_release_valid(L2BroadcastHub_8569_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(L2BroadcastHub_8569_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(L2BroadcastHub_8569_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(L2BroadcastHub_8569_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(L2BroadcastHub_8569_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(L2BroadcastHub_8569_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(L2BroadcastHub_8569_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(L2BroadcastHub_8569_io_inner_release_bits_client_id),
    .io_incoherent_0(L2BroadcastHub_8569_io_incoherent_0),
    .io_outer_acquire_ready(L2BroadcastHub_8569_io_outer_acquire_ready),
    .io_outer_acquire_valid(L2BroadcastHub_8569_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(L2BroadcastHub_8569_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(L2BroadcastHub_8569_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(L2BroadcastHub_8569_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(L2BroadcastHub_8569_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(L2BroadcastHub_8569_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(L2BroadcastHub_8569_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(L2BroadcastHub_8569_io_outer_acquire_bits_data),
    .io_outer_grant_ready(L2BroadcastHub_8569_io_outer_grant_ready),
    .io_outer_grant_valid(L2BroadcastHub_8569_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(L2BroadcastHub_8569_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(L2BroadcastHub_8569_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(L2BroadcastHub_8569_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(L2BroadcastHub_8569_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(L2BroadcastHub_8569_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(L2BroadcastHub_8569_io_outer_grant_bits_data)
  );
  MMIOTileLinkManager mmioManager (
    .clk(mmioManager_clk),
    .reset(mmioManager_reset),
    .io_inner_acquire_ready(mmioManager_io_inner_acquire_ready),
    .io_inner_acquire_valid(mmioManager_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(mmioManager_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(mmioManager_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(mmioManager_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(mmioManager_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(mmioManager_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(mmioManager_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(mmioManager_io_inner_acquire_bits_data),
    .io_inner_acquire_bits_client_id(mmioManager_io_inner_acquire_bits_client_id),
    .io_inner_grant_ready(mmioManager_io_inner_grant_ready),
    .io_inner_grant_valid(mmioManager_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(mmioManager_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(mmioManager_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(mmioManager_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(mmioManager_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(mmioManager_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(mmioManager_io_inner_grant_bits_data),
    .io_inner_grant_bits_client_id(mmioManager_io_inner_grant_bits_client_id),
    .io_inner_finish_ready(mmioManager_io_inner_finish_ready),
    .io_inner_finish_valid(mmioManager_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(mmioManager_io_inner_finish_bits_manager_xact_id),
    .io_inner_probe_ready(mmioManager_io_inner_probe_ready),
    .io_inner_probe_valid(mmioManager_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(mmioManager_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(mmioManager_io_inner_probe_bits_p_type),
    .io_inner_probe_bits_client_id(mmioManager_io_inner_probe_bits_client_id),
    .io_inner_release_ready(mmioManager_io_inner_release_ready),
    .io_inner_release_valid(mmioManager_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(mmioManager_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(mmioManager_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(mmioManager_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(mmioManager_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(mmioManager_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(mmioManager_io_inner_release_bits_data),
    .io_inner_release_bits_client_id(mmioManager_io_inner_release_bits_client_id),
    .io_incoherent_0(mmioManager_io_incoherent_0),
    .io_outer_acquire_ready(mmioManager_io_outer_acquire_ready),
    .io_outer_acquire_valid(mmioManager_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(mmioManager_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(mmioManager_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(mmioManager_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(mmioManager_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(mmioManager_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(mmioManager_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(mmioManager_io_outer_acquire_bits_data),
    .io_outer_grant_ready(mmioManager_io_outer_grant_ready),
    .io_outer_grant_valid(mmioManager_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(mmioManager_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(mmioManager_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(mmioManager_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(mmioManager_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(mmioManager_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(mmioManager_io_outer_grant_bits_data)
  );
  TileLinkMemoryInterconnect mem_ic (
    .clk(mem_ic_clk),
    .reset(mem_ic_reset),
    .io_in_0_acquire_ready(mem_ic_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(mem_ic_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(mem_ic_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(mem_ic_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(mem_ic_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(mem_ic_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(mem_ic_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(mem_ic_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(mem_ic_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(mem_ic_io_in_0_grant_ready),
    .io_in_0_grant_valid(mem_ic_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(mem_ic_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(mem_ic_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(mem_ic_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(mem_ic_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(mem_ic_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(mem_ic_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(mem_ic_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(mem_ic_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(mem_ic_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(mem_ic_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(mem_ic_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(mem_ic_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(mem_ic_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(mem_ic_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(mem_ic_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(mem_ic_io_out_0_grant_ready),
    .io_out_0_grant_valid(mem_ic_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(mem_ic_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(mem_ic_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(mem_ic_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(mem_ic_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(mem_ic_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(mem_ic_io_out_0_grant_bits_data)
  );
  ClientTileLinkIOUnwrapper ClientTileLinkIOUnwrapper_8570 (
    .clk(ClientTileLinkIOUnwrapper_8570_clk),
    .reset(ClientTileLinkIOUnwrapper_8570_reset),
    .io_in_acquire_ready(ClientTileLinkIOUnwrapper_8570_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOUnwrapper_8570_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_data),
    .io_in_probe_ready(ClientTileLinkIOUnwrapper_8570_io_in_probe_ready),
    .io_in_probe_valid(ClientTileLinkIOUnwrapper_8570_io_in_probe_valid),
    .io_in_probe_bits_addr_block(ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_addr_block),
    .io_in_probe_bits_p_type(ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_p_type),
    .io_in_release_ready(ClientTileLinkIOUnwrapper_8570_io_in_release_ready),
    .io_in_release_valid(ClientTileLinkIOUnwrapper_8570_io_in_release_valid),
    .io_in_release_bits_addr_beat(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_beat),
    .io_in_release_bits_addr_block(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_block),
    .io_in_release_bits_client_xact_id(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_client_xact_id),
    .io_in_release_bits_voluntary(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_voluntary),
    .io_in_release_bits_r_type(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_r_type),
    .io_in_release_bits_data(ClientTileLinkIOUnwrapper_8570_io_in_release_bits_data),
    .io_in_grant_ready(ClientTileLinkIOUnwrapper_8570_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOUnwrapper_8570_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_data),
    .io_in_grant_bits_manager_id(ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_id),
    .io_in_finish_ready(ClientTileLinkIOUnwrapper_8570_io_in_finish_ready),
    .io_in_finish_valid(ClientTileLinkIOUnwrapper_8570_io_in_finish_valid),
    .io_in_finish_bits_manager_xact_id(ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_xact_id),
    .io_in_finish_bits_manager_id(ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_id),
    .io_out_acquire_ready(ClientTileLinkIOUnwrapper_8570_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOUnwrapper_8570_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_data),
    .io_out_grant_ready(ClientTileLinkIOUnwrapper_8570_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOUnwrapper_8570_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_data)
  );
  ClientTileLinkIOWrapper ClientTileLinkIOWrapper_8571 (
    .clk(ClientTileLinkIOWrapper_8571_clk),
    .reset(ClientTileLinkIOWrapper_8571_reset),
    .io_in_acquire_ready(ClientTileLinkIOWrapper_8571_io_in_acquire_ready),
    .io_in_acquire_valid(ClientTileLinkIOWrapper_8571_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientTileLinkIOWrapper_8571_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientTileLinkIOWrapper_8571_io_in_grant_ready),
    .io_in_grant_valid(ClientTileLinkIOWrapper_8571_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientTileLinkIOWrapper_8571_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientTileLinkIOWrapper_8571_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientTileLinkIOWrapper_8571_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientTileLinkIOWrapper_8571_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientTileLinkIOWrapper_8571_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientTileLinkIOWrapper_8571_io_in_grant_bits_data),
    .io_out_acquire_ready(ClientTileLinkIOWrapper_8571_io_out_acquire_ready),
    .io_out_acquire_valid(ClientTileLinkIOWrapper_8571_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(ClientTileLinkIOWrapper_8571_io_out_acquire_bits_data),
    .io_out_probe_ready(ClientTileLinkIOWrapper_8571_io_out_probe_ready),
    .io_out_probe_valid(ClientTileLinkIOWrapper_8571_io_out_probe_valid),
    .io_out_probe_bits_addr_block(ClientTileLinkIOWrapper_8571_io_out_probe_bits_addr_block),
    .io_out_probe_bits_p_type(ClientTileLinkIOWrapper_8571_io_out_probe_bits_p_type),
    .io_out_release_ready(ClientTileLinkIOWrapper_8571_io_out_release_ready),
    .io_out_release_valid(ClientTileLinkIOWrapper_8571_io_out_release_valid),
    .io_out_release_bits_addr_beat(ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_beat),
    .io_out_release_bits_addr_block(ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_block),
    .io_out_release_bits_client_xact_id(ClientTileLinkIOWrapper_8571_io_out_release_bits_client_xact_id),
    .io_out_release_bits_voluntary(ClientTileLinkIOWrapper_8571_io_out_release_bits_voluntary),
    .io_out_release_bits_r_type(ClientTileLinkIOWrapper_8571_io_out_release_bits_r_type),
    .io_out_release_bits_data(ClientTileLinkIOWrapper_8571_io_out_release_bits_data),
    .io_out_grant_ready(ClientTileLinkIOWrapper_8571_io_out_grant_ready),
    .io_out_grant_valid(ClientTileLinkIOWrapper_8571_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(ClientTileLinkIOWrapper_8571_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(ClientTileLinkIOWrapper_8571_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(ClientTileLinkIOWrapper_8571_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(ClientTileLinkIOWrapper_8571_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(ClientTileLinkIOWrapper_8571_io_out_grant_bits_data),
    .io_out_grant_bits_manager_id(ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_id),
    .io_out_finish_ready(ClientTileLinkIOWrapper_8571_io_out_finish_ready),
    .io_out_finish_valid(ClientTileLinkIOWrapper_8571_io_out_finish_valid),
    .io_out_finish_bits_manager_xact_id(ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_xact_id),
    .io_out_finish_bits_manager_id(ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_id)
  );
  ClientTileLinkEnqueuer ClientTileLinkEnqueuer_8572 (
    .clk(ClientTileLinkEnqueuer_8572_clk),
    .reset(ClientTileLinkEnqueuer_8572_reset),
    .io_inner_acquire_ready(ClientTileLinkEnqueuer_8572_io_inner_acquire_ready),
    .io_inner_acquire_valid(ClientTileLinkEnqueuer_8572_io_inner_acquire_valid),
    .io_inner_acquire_bits_addr_block(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_block),
    .io_inner_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_client_xact_id),
    .io_inner_acquire_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_beat),
    .io_inner_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_is_builtin_type),
    .io_inner_acquire_bits_a_type(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_a_type),
    .io_inner_acquire_bits_union(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_union),
    .io_inner_acquire_bits_data(ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_data),
    .io_inner_probe_ready(ClientTileLinkEnqueuer_8572_io_inner_probe_ready),
    .io_inner_probe_valid(ClientTileLinkEnqueuer_8572_io_inner_probe_valid),
    .io_inner_probe_bits_addr_block(ClientTileLinkEnqueuer_8572_io_inner_probe_bits_addr_block),
    .io_inner_probe_bits_p_type(ClientTileLinkEnqueuer_8572_io_inner_probe_bits_p_type),
    .io_inner_release_ready(ClientTileLinkEnqueuer_8572_io_inner_release_ready),
    .io_inner_release_valid(ClientTileLinkEnqueuer_8572_io_inner_release_valid),
    .io_inner_release_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_beat),
    .io_inner_release_bits_addr_block(ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_block),
    .io_inner_release_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_inner_release_bits_client_xact_id),
    .io_inner_release_bits_voluntary(ClientTileLinkEnqueuer_8572_io_inner_release_bits_voluntary),
    .io_inner_release_bits_r_type(ClientTileLinkEnqueuer_8572_io_inner_release_bits_r_type),
    .io_inner_release_bits_data(ClientTileLinkEnqueuer_8572_io_inner_release_bits_data),
    .io_inner_grant_ready(ClientTileLinkEnqueuer_8572_io_inner_grant_ready),
    .io_inner_grant_valid(ClientTileLinkEnqueuer_8572_io_inner_grant_valid),
    .io_inner_grant_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_addr_beat),
    .io_inner_grant_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_client_xact_id),
    .io_inner_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_xact_id),
    .io_inner_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_is_builtin_type),
    .io_inner_grant_bits_g_type(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_g_type),
    .io_inner_grant_bits_data(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_data),
    .io_inner_grant_bits_manager_id(ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_id),
    .io_inner_finish_ready(ClientTileLinkEnqueuer_8572_io_inner_finish_ready),
    .io_inner_finish_valid(ClientTileLinkEnqueuer_8572_io_inner_finish_valid),
    .io_inner_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_xact_id),
    .io_inner_finish_bits_manager_id(ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_id),
    .io_outer_acquire_ready(ClientTileLinkEnqueuer_8572_io_outer_acquire_ready),
    .io_outer_acquire_valid(ClientTileLinkEnqueuer_8572_io_outer_acquire_valid),
    .io_outer_acquire_bits_addr_block(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_block),
    .io_outer_acquire_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_client_xact_id),
    .io_outer_acquire_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_beat),
    .io_outer_acquire_bits_is_builtin_type(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_is_builtin_type),
    .io_outer_acquire_bits_a_type(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_a_type),
    .io_outer_acquire_bits_union(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_union),
    .io_outer_acquire_bits_data(ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_data),
    .io_outer_probe_ready(ClientTileLinkEnqueuer_8572_io_outer_probe_ready),
    .io_outer_probe_valid(ClientTileLinkEnqueuer_8572_io_outer_probe_valid),
    .io_outer_probe_bits_addr_block(ClientTileLinkEnqueuer_8572_io_outer_probe_bits_addr_block),
    .io_outer_probe_bits_p_type(ClientTileLinkEnqueuer_8572_io_outer_probe_bits_p_type),
    .io_outer_release_ready(ClientTileLinkEnqueuer_8572_io_outer_release_ready),
    .io_outer_release_valid(ClientTileLinkEnqueuer_8572_io_outer_release_valid),
    .io_outer_release_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_beat),
    .io_outer_release_bits_addr_block(ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_block),
    .io_outer_release_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_outer_release_bits_client_xact_id),
    .io_outer_release_bits_voluntary(ClientTileLinkEnqueuer_8572_io_outer_release_bits_voluntary),
    .io_outer_release_bits_r_type(ClientTileLinkEnqueuer_8572_io_outer_release_bits_r_type),
    .io_outer_release_bits_data(ClientTileLinkEnqueuer_8572_io_outer_release_bits_data),
    .io_outer_grant_ready(ClientTileLinkEnqueuer_8572_io_outer_grant_ready),
    .io_outer_grant_valid(ClientTileLinkEnqueuer_8572_io_outer_grant_valid),
    .io_outer_grant_bits_addr_beat(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_addr_beat),
    .io_outer_grant_bits_client_xact_id(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_client_xact_id),
    .io_outer_grant_bits_manager_xact_id(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_xact_id),
    .io_outer_grant_bits_is_builtin_type(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_is_builtin_type),
    .io_outer_grant_bits_g_type(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_g_type),
    .io_outer_grant_bits_data(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_data),
    .io_outer_grant_bits_manager_id(ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_id),
    .io_outer_finish_ready(ClientTileLinkEnqueuer_8572_io_outer_finish_ready),
    .io_outer_finish_valid(ClientTileLinkEnqueuer_8572_io_outer_finish_valid),
    .io_outer_finish_bits_manager_xact_id(ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_xact_id),
    .io_outer_finish_bits_manager_id(ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_id)
  );
  NastiIOTileLinkIOConverter NastiIOTileLinkIOConverter_8573 (
    .clk(NastiIOTileLinkIOConverter_8573_clk),
    .reset(NastiIOTileLinkIOConverter_8573_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_8573_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_8573_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_8573_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_8573_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_8573_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_8573_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_8573_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_8573_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_8573_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_8573_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_8573_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_8573_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_8573_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_8573_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_user)
  );
  Queue_39 Queue_39_8586 (
    .clk(Queue_39_8586_clk),
    .reset(Queue_39_8586_reset),
    .io_enq_ready(Queue_39_8586_io_enq_ready),
    .io_enq_valid(Queue_39_8586_io_enq_valid),
    .io_enq_bits_addr(Queue_39_8586_io_enq_bits_addr),
    .io_enq_bits_len(Queue_39_8586_io_enq_bits_len),
    .io_enq_bits_size(Queue_39_8586_io_enq_bits_size),
    .io_enq_bits_burst(Queue_39_8586_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_39_8586_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_39_8586_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_39_8586_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_39_8586_io_enq_bits_qos),
    .io_enq_bits_region(Queue_39_8586_io_enq_bits_region),
    .io_enq_bits_id(Queue_39_8586_io_enq_bits_id),
    .io_enq_bits_user(Queue_39_8586_io_enq_bits_user),
    .io_deq_ready(Queue_39_8586_io_deq_ready),
    .io_deq_valid(Queue_39_8586_io_deq_valid),
    .io_deq_bits_addr(Queue_39_8586_io_deq_bits_addr),
    .io_deq_bits_len(Queue_39_8586_io_deq_bits_len),
    .io_deq_bits_size(Queue_39_8586_io_deq_bits_size),
    .io_deq_bits_burst(Queue_39_8586_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_39_8586_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_39_8586_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_39_8586_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_39_8586_io_deq_bits_qos),
    .io_deq_bits_region(Queue_39_8586_io_deq_bits_region),
    .io_deq_bits_id(Queue_39_8586_io_deq_bits_id),
    .io_deq_bits_user(Queue_39_8586_io_deq_bits_user),
    .io_count(Queue_39_8586_io_count)
  );
  Queue_39 Queue_40_8599 (
    .clk(Queue_40_8599_clk),
    .reset(Queue_40_8599_reset),
    .io_enq_ready(Queue_40_8599_io_enq_ready),
    .io_enq_valid(Queue_40_8599_io_enq_valid),
    .io_enq_bits_addr(Queue_40_8599_io_enq_bits_addr),
    .io_enq_bits_len(Queue_40_8599_io_enq_bits_len),
    .io_enq_bits_size(Queue_40_8599_io_enq_bits_size),
    .io_enq_bits_burst(Queue_40_8599_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_40_8599_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_40_8599_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_40_8599_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_40_8599_io_enq_bits_qos),
    .io_enq_bits_region(Queue_40_8599_io_enq_bits_region),
    .io_enq_bits_id(Queue_40_8599_io_enq_bits_id),
    .io_enq_bits_user(Queue_40_8599_io_enq_bits_user),
    .io_deq_ready(Queue_40_8599_io_deq_ready),
    .io_deq_valid(Queue_40_8599_io_deq_valid),
    .io_deq_bits_addr(Queue_40_8599_io_deq_bits_addr),
    .io_deq_bits_len(Queue_40_8599_io_deq_bits_len),
    .io_deq_bits_size(Queue_40_8599_io_deq_bits_size),
    .io_deq_bits_burst(Queue_40_8599_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_40_8599_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_40_8599_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_40_8599_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_40_8599_io_deq_bits_qos),
    .io_deq_bits_region(Queue_40_8599_io_deq_bits_region),
    .io_deq_bits_id(Queue_40_8599_io_deq_bits_id),
    .io_deq_bits_user(Queue_40_8599_io_deq_bits_user),
    .io_count(Queue_40_8599_io_count)
  );
  Queue_41 Queue_41_8606 (
    .clk(Queue_41_8606_clk),
    .reset(Queue_41_8606_reset),
    .io_enq_ready(Queue_41_8606_io_enq_ready),
    .io_enq_valid(Queue_41_8606_io_enq_valid),
    .io_enq_bits_data(Queue_41_8606_io_enq_bits_data),
    .io_enq_bits_last(Queue_41_8606_io_enq_bits_last),
    .io_enq_bits_id(Queue_41_8606_io_enq_bits_id),
    .io_enq_bits_strb(Queue_41_8606_io_enq_bits_strb),
    .io_enq_bits_user(Queue_41_8606_io_enq_bits_user),
    .io_deq_ready(Queue_41_8606_io_deq_ready),
    .io_deq_valid(Queue_41_8606_io_deq_valid),
    .io_deq_bits_data(Queue_41_8606_io_deq_bits_data),
    .io_deq_bits_last(Queue_41_8606_io_deq_bits_last),
    .io_deq_bits_id(Queue_41_8606_io_deq_bits_id),
    .io_deq_bits_strb(Queue_41_8606_io_deq_bits_strb),
    .io_deq_bits_user(Queue_41_8606_io_deq_bits_user),
    .io_count(Queue_41_8606_io_count)
  );
  Queue_42 Queue_42_8613 (
    .clk(Queue_42_8613_clk),
    .reset(Queue_42_8613_reset),
    .io_enq_ready(Queue_42_8613_io_enq_ready),
    .io_enq_valid(Queue_42_8613_io_enq_valid),
    .io_enq_bits_resp(Queue_42_8613_io_enq_bits_resp),
    .io_enq_bits_data(Queue_42_8613_io_enq_bits_data),
    .io_enq_bits_last(Queue_42_8613_io_enq_bits_last),
    .io_enq_bits_id(Queue_42_8613_io_enq_bits_id),
    .io_enq_bits_user(Queue_42_8613_io_enq_bits_user),
    .io_deq_ready(Queue_42_8613_io_deq_ready),
    .io_deq_valid(Queue_42_8613_io_deq_valid),
    .io_deq_bits_resp(Queue_42_8613_io_deq_bits_resp),
    .io_deq_bits_data(Queue_42_8613_io_deq_bits_data),
    .io_deq_bits_last(Queue_42_8613_io_deq_bits_last),
    .io_deq_bits_id(Queue_42_8613_io_deq_bits_id),
    .io_deq_bits_user(Queue_42_8613_io_deq_bits_user),
    .io_count(Queue_42_8613_io_count)
  );
  Queue_43 Queue_43_8618 (
    .clk(Queue_43_8618_clk),
    .reset(Queue_43_8618_reset),
    .io_enq_ready(Queue_43_8618_io_enq_ready),
    .io_enq_valid(Queue_43_8618_io_enq_valid),
    .io_enq_bits_resp(Queue_43_8618_io_enq_bits_resp),
    .io_enq_bits_id(Queue_43_8618_io_enq_bits_id),
    .io_enq_bits_user(Queue_43_8618_io_enq_bits_user),
    .io_deq_ready(Queue_43_8618_io_deq_ready),
    .io_deq_valid(Queue_43_8618_io_deq_valid),
    .io_deq_bits_resp(Queue_43_8618_io_deq_bits_resp),
    .io_deq_bits_id(Queue_43_8618_io_deq_bits_id),
    .io_deq_bits_user(Queue_43_8618_io_deq_bits_user),
    .io_count(Queue_43_8618_io_count)
  );
  assign io_tiles_cached_0_acquire_ready = l1tol2net_io_clients_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = l1tol2net_io_clients_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = l1tol2net_io_clients_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = l1tol2net_io_clients_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = l1tol2net_io_clients_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = l1tol2net_io_clients_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = l1tol2net_io_clients_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = l1tol2net_io_clients_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = l1tol2net_io_clients_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = l1tol2net_io_clients_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = l1tol2net_io_clients_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = l1tol2net_io_clients_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = l1tol2net_io_clients_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = l1tol2net_io_clients_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = l1tol2net_io_clients_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = l1tol2net_io_clients_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = l1tol2net_io_clients_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = l1tol2net_io_clients_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = l1tol2net_io_clients_uncached_0_grant_bits_data;
  assign io_htif_uncached_acquire_ready = l1tol2net_io_clients_uncached_1_acquire_ready;
  assign io_htif_uncached_grant_valid = l1tol2net_io_clients_uncached_1_grant_valid;
  assign io_htif_uncached_grant_bits_addr_beat = l1tol2net_io_clients_uncached_1_grant_bits_addr_beat;
  assign io_htif_uncached_grant_bits_client_xact_id = l1tol2net_io_clients_uncached_1_grant_bits_client_xact_id;
  assign io_htif_uncached_grant_bits_manager_xact_id = l1tol2net_io_clients_uncached_1_grant_bits_manager_xact_id;
  assign io_htif_uncached_grant_bits_is_builtin_type = l1tol2net_io_clients_uncached_1_grant_bits_is_builtin_type;
  assign io_htif_uncached_grant_bits_g_type = l1tol2net_io_clients_uncached_1_grant_bits_g_type;
  assign io_htif_uncached_grant_bits_data = l1tol2net_io_clients_uncached_1_grant_bits_data;
  assign io_mem_axi_0_aw_valid = Queue_40_8599_io_deq_valid;
  assign io_mem_axi_0_aw_bits_addr = Queue_40_8599_io_deq_bits_addr;
  assign io_mem_axi_0_aw_bits_len = Queue_40_8599_io_deq_bits_len;
  assign io_mem_axi_0_aw_bits_size = Queue_40_8599_io_deq_bits_size;
  assign io_mem_axi_0_aw_bits_burst = Queue_40_8599_io_deq_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = Queue_40_8599_io_deq_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = 4'h3;
  assign io_mem_axi_0_aw_bits_prot = Queue_40_8599_io_deq_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = Queue_40_8599_io_deq_bits_qos;
  assign io_mem_axi_0_aw_bits_region = Queue_40_8599_io_deq_bits_region;
  assign io_mem_axi_0_aw_bits_id = Queue_40_8599_io_deq_bits_id;
  assign io_mem_axi_0_aw_bits_user = Queue_40_8599_io_deq_bits_user;
  assign io_mem_axi_0_w_valid = Queue_41_8606_io_deq_valid;
  assign io_mem_axi_0_w_bits_data = Queue_41_8606_io_deq_bits_data;
  assign io_mem_axi_0_w_bits_last = Queue_41_8606_io_deq_bits_last;
  assign io_mem_axi_0_w_bits_id = Queue_41_8606_io_deq_bits_id;
  assign io_mem_axi_0_w_bits_strb = Queue_41_8606_io_deq_bits_strb;
  assign io_mem_axi_0_w_bits_user = Queue_41_8606_io_deq_bits_user;
  assign io_mem_axi_0_b_ready = Queue_43_8618_io_enq_ready;
  assign io_mem_axi_0_ar_valid = Queue_39_8586_io_deq_valid;
  assign io_mem_axi_0_ar_bits_addr = Queue_39_8586_io_deq_bits_addr;
  assign io_mem_axi_0_ar_bits_len = Queue_39_8586_io_deq_bits_len;
  assign io_mem_axi_0_ar_bits_size = Queue_39_8586_io_deq_bits_size;
  assign io_mem_axi_0_ar_bits_burst = Queue_39_8586_io_deq_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = Queue_39_8586_io_deq_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = 4'h3;
  assign io_mem_axi_0_ar_bits_prot = Queue_39_8586_io_deq_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = Queue_39_8586_io_deq_bits_qos;
  assign io_mem_axi_0_ar_bits_region = Queue_39_8586_io_deq_bits_region;
  assign io_mem_axi_0_ar_bits_id = Queue_39_8586_io_deq_bits_id;
  assign io_mem_axi_0_ar_bits_user = Queue_39_8586_io_deq_bits_user;
  assign io_mem_axi_0_r_ready = Queue_42_8613_io_enq_ready;
  assign io_mmio_acquire_valid = mmioManager_io_outer_acquire_valid;
  assign io_mmio_acquire_bits_addr_block = mmioManager_io_outer_acquire_bits_addr_block;
  assign io_mmio_acquire_bits_client_xact_id = mmioManager_io_outer_acquire_bits_client_xact_id;
  assign io_mmio_acquire_bits_addr_beat = mmioManager_io_outer_acquire_bits_addr_beat;
  assign io_mmio_acquire_bits_is_builtin_type = mmioManager_io_outer_acquire_bits_is_builtin_type;
  assign io_mmio_acquire_bits_a_type = mmioManager_io_outer_acquire_bits_a_type;
  assign io_mmio_acquire_bits_union = mmioManager_io_outer_acquire_bits_union;
  assign io_mmio_acquire_bits_data = mmioManager_io_outer_acquire_bits_data;
  assign io_mmio_grant_ready = mmioManager_io_outer_grant_ready;
  assign l1tol2net_clk = clk;
  assign l1tol2net_reset = reset;
  assign l1tol2net_io_clients_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign l1tol2net_io_clients_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign l1tol2net_io_clients_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign l1tol2net_io_clients_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign l1tol2net_io_clients_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign l1tol2net_io_clients_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign l1tol2net_io_clients_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign l1tol2net_io_clients_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign l1tol2net_io_clients_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign l1tol2net_io_clients_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign l1tol2net_io_clients_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign l1tol2net_io_clients_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign l1tol2net_io_clients_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign l1tol2net_io_clients_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign l1tol2net_io_clients_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign l1tol2net_io_clients_uncached_1_acquire_valid = io_htif_uncached_acquire_valid;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_addr_block = io_htif_uncached_acquire_bits_addr_block;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_client_xact_id = io_htif_uncached_acquire_bits_client_xact_id;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_addr_beat = io_htif_uncached_acquire_bits_addr_beat;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_is_builtin_type = io_htif_uncached_acquire_bits_is_builtin_type;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_a_type = io_htif_uncached_acquire_bits_a_type;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_union = io_htif_uncached_acquire_bits_union;
  assign l1tol2net_io_clients_uncached_1_acquire_bits_data = io_htif_uncached_acquire_bits_data;
  assign l1tol2net_io_clients_uncached_1_grant_ready = io_htif_uncached_grant_ready;
  assign l1tol2net_io_managers_0_acquire_ready = L2BroadcastHub_8569_io_inner_acquire_ready;
  assign l1tol2net_io_managers_0_grant_valid = L2BroadcastHub_8569_io_inner_grant_valid;
  assign l1tol2net_io_managers_0_grant_bits_addr_beat = L2BroadcastHub_8569_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_0_grant_bits_client_xact_id = L2BroadcastHub_8569_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_manager_xact_id = L2BroadcastHub_8569_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_0_grant_bits_is_builtin_type = L2BroadcastHub_8569_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_0_grant_bits_g_type = L2BroadcastHub_8569_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_0_grant_bits_data = L2BroadcastHub_8569_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_0_grant_bits_client_id = L2BroadcastHub_8569_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_0_finish_ready = L2BroadcastHub_8569_io_inner_finish_ready;
  assign l1tol2net_io_managers_0_probe_valid = L2BroadcastHub_8569_io_inner_probe_valid;
  assign l1tol2net_io_managers_0_probe_bits_addr_block = L2BroadcastHub_8569_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_0_probe_bits_p_type = L2BroadcastHub_8569_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_0_probe_bits_client_id = L2BroadcastHub_8569_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_0_release_ready = L2BroadcastHub_8569_io_inner_release_ready;
  assign l1tol2net_io_managers_1_acquire_ready = mmioManager_io_inner_acquire_ready;
  assign l1tol2net_io_managers_1_grant_valid = mmioManager_io_inner_grant_valid;
  assign l1tol2net_io_managers_1_grant_bits_addr_beat = mmioManager_io_inner_grant_bits_addr_beat;
  assign l1tol2net_io_managers_1_grant_bits_client_xact_id = mmioManager_io_inner_grant_bits_client_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_manager_xact_id = mmioManager_io_inner_grant_bits_manager_xact_id;
  assign l1tol2net_io_managers_1_grant_bits_is_builtin_type = mmioManager_io_inner_grant_bits_is_builtin_type;
  assign l1tol2net_io_managers_1_grant_bits_g_type = mmioManager_io_inner_grant_bits_g_type;
  assign l1tol2net_io_managers_1_grant_bits_data = mmioManager_io_inner_grant_bits_data;
  assign l1tol2net_io_managers_1_grant_bits_client_id = mmioManager_io_inner_grant_bits_client_id;
  assign l1tol2net_io_managers_1_finish_ready = mmioManager_io_inner_finish_ready;
  assign l1tol2net_io_managers_1_probe_valid = mmioManager_io_inner_probe_valid;
  assign l1tol2net_io_managers_1_probe_bits_addr_block = mmioManager_io_inner_probe_bits_addr_block;
  assign l1tol2net_io_managers_1_probe_bits_p_type = mmioManager_io_inner_probe_bits_p_type;
  assign l1tol2net_io_managers_1_probe_bits_client_id = mmioManager_io_inner_probe_bits_client_id;
  assign l1tol2net_io_managers_1_release_ready = mmioManager_io_inner_release_ready;
  assign L2BroadcastHub_8569_clk = clk;
  assign L2BroadcastHub_8569_reset = reset;
  assign L2BroadcastHub_8569_io_inner_acquire_valid = l1tol2net_io_managers_0_acquire_valid;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_0_acquire_bits_addr_block;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_0_acquire_bits_client_xact_id;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_0_acquire_bits_addr_beat;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_0_acquire_bits_is_builtin_type;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_a_type = l1tol2net_io_managers_0_acquire_bits_a_type;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_union = l1tol2net_io_managers_0_acquire_bits_union;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_data = l1tol2net_io_managers_0_acquire_bits_data;
  assign L2BroadcastHub_8569_io_inner_acquire_bits_client_id = l1tol2net_io_managers_0_acquire_bits_client_id;
  assign L2BroadcastHub_8569_io_inner_grant_ready = l1tol2net_io_managers_0_grant_ready;
  assign L2BroadcastHub_8569_io_inner_finish_valid = l1tol2net_io_managers_0_finish_valid;
  assign L2BroadcastHub_8569_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_0_finish_bits_manager_xact_id;
  assign L2BroadcastHub_8569_io_inner_probe_ready = l1tol2net_io_managers_0_probe_ready;
  assign L2BroadcastHub_8569_io_inner_release_valid = l1tol2net_io_managers_0_release_valid;
  assign L2BroadcastHub_8569_io_inner_release_bits_addr_beat = l1tol2net_io_managers_0_release_bits_addr_beat;
  assign L2BroadcastHub_8569_io_inner_release_bits_addr_block = l1tol2net_io_managers_0_release_bits_addr_block;
  assign L2BroadcastHub_8569_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_0_release_bits_client_xact_id;
  assign L2BroadcastHub_8569_io_inner_release_bits_voluntary = l1tol2net_io_managers_0_release_bits_voluntary;
  assign L2BroadcastHub_8569_io_inner_release_bits_r_type = l1tol2net_io_managers_0_release_bits_r_type;
  assign L2BroadcastHub_8569_io_inner_release_bits_data = l1tol2net_io_managers_0_release_bits_data;
  assign L2BroadcastHub_8569_io_inner_release_bits_client_id = l1tol2net_io_managers_0_release_bits_client_id;
  assign L2BroadcastHub_8569_io_incoherent_0 = io_incoherent_0;
  assign L2BroadcastHub_8569_io_outer_acquire_ready = ClientTileLinkIOWrapper_8571_io_in_acquire_ready;
  assign L2BroadcastHub_8569_io_outer_grant_valid = ClientTileLinkIOWrapper_8571_io_in_grant_valid;
  assign L2BroadcastHub_8569_io_outer_grant_bits_addr_beat = ClientTileLinkIOWrapper_8571_io_in_grant_bits_addr_beat;
  assign L2BroadcastHub_8569_io_outer_grant_bits_client_xact_id = ClientTileLinkIOWrapper_8571_io_in_grant_bits_client_xact_id;
  assign L2BroadcastHub_8569_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOWrapper_8571_io_in_grant_bits_manager_xact_id;
  assign L2BroadcastHub_8569_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOWrapper_8571_io_in_grant_bits_is_builtin_type;
  assign L2BroadcastHub_8569_io_outer_grant_bits_g_type = ClientTileLinkIOWrapper_8571_io_in_grant_bits_g_type;
  assign L2BroadcastHub_8569_io_outer_grant_bits_data = ClientTileLinkIOWrapper_8571_io_in_grant_bits_data;
  assign mmioManager_clk = clk;
  assign mmioManager_reset = reset;
  assign mmioManager_io_inner_acquire_valid = l1tol2net_io_managers_1_acquire_valid;
  assign mmioManager_io_inner_acquire_bits_addr_block = l1tol2net_io_managers_1_acquire_bits_addr_block;
  assign mmioManager_io_inner_acquire_bits_client_xact_id = l1tol2net_io_managers_1_acquire_bits_client_xact_id;
  assign mmioManager_io_inner_acquire_bits_addr_beat = l1tol2net_io_managers_1_acquire_bits_addr_beat;
  assign mmioManager_io_inner_acquire_bits_is_builtin_type = l1tol2net_io_managers_1_acquire_bits_is_builtin_type;
  assign mmioManager_io_inner_acquire_bits_a_type = l1tol2net_io_managers_1_acquire_bits_a_type;
  assign mmioManager_io_inner_acquire_bits_union = l1tol2net_io_managers_1_acquire_bits_union;
  assign mmioManager_io_inner_acquire_bits_data = l1tol2net_io_managers_1_acquire_bits_data;
  assign mmioManager_io_inner_acquire_bits_client_id = l1tol2net_io_managers_1_acquire_bits_client_id;
  assign mmioManager_io_inner_grant_ready = l1tol2net_io_managers_1_grant_ready;
  assign mmioManager_io_inner_finish_valid = l1tol2net_io_managers_1_finish_valid;
  assign mmioManager_io_inner_finish_bits_manager_xact_id = l1tol2net_io_managers_1_finish_bits_manager_xact_id;
  assign mmioManager_io_inner_probe_ready = l1tol2net_io_managers_1_probe_ready;
  assign mmioManager_io_inner_release_valid = l1tol2net_io_managers_1_release_valid;
  assign mmioManager_io_inner_release_bits_addr_beat = l1tol2net_io_managers_1_release_bits_addr_beat;
  assign mmioManager_io_inner_release_bits_addr_block = l1tol2net_io_managers_1_release_bits_addr_block;
  assign mmioManager_io_inner_release_bits_client_xact_id = l1tol2net_io_managers_1_release_bits_client_xact_id;
  assign mmioManager_io_inner_release_bits_voluntary = l1tol2net_io_managers_1_release_bits_voluntary;
  assign mmioManager_io_inner_release_bits_r_type = l1tol2net_io_managers_1_release_bits_r_type;
  assign mmioManager_io_inner_release_bits_data = l1tol2net_io_managers_1_release_bits_data;
  assign mmioManager_io_inner_release_bits_client_id = l1tol2net_io_managers_1_release_bits_client_id;
  assign mmioManager_io_incoherent_0 = GEN_0;
  assign mmioManager_io_outer_acquire_ready = io_mmio_acquire_ready;
  assign mmioManager_io_outer_grant_valid = io_mmio_grant_valid;
  assign mmioManager_io_outer_grant_bits_addr_beat = io_mmio_grant_bits_addr_beat;
  assign mmioManager_io_outer_grant_bits_client_xact_id = io_mmio_grant_bits_client_xact_id;
  assign mmioManager_io_outer_grant_bits_manager_xact_id = io_mmio_grant_bits_manager_xact_id;
  assign mmioManager_io_outer_grant_bits_is_builtin_type = io_mmio_grant_bits_is_builtin_type;
  assign mmioManager_io_outer_grant_bits_g_type = io_mmio_grant_bits_g_type;
  assign mmioManager_io_outer_grant_bits_data = io_mmio_grant_bits_data;
  assign mem_ic_clk = clk;
  assign mem_ic_reset = reset;
  assign mem_ic_io_in_0_acquire_valid = ClientTileLinkIOUnwrapper_8570_io_out_acquire_valid;
  assign mem_ic_io_in_0_acquire_bits_addr_block = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_block;
  assign mem_ic_io_in_0_acquire_bits_client_xact_id = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_client_xact_id;
  assign mem_ic_io_in_0_acquire_bits_addr_beat = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_addr_beat;
  assign mem_ic_io_in_0_acquire_bits_is_builtin_type = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_is_builtin_type;
  assign mem_ic_io_in_0_acquire_bits_a_type = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_a_type;
  assign mem_ic_io_in_0_acquire_bits_union = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_union;
  assign mem_ic_io_in_0_acquire_bits_data = ClientTileLinkIOUnwrapper_8570_io_out_acquire_bits_data;
  assign mem_ic_io_in_0_grant_ready = ClientTileLinkIOUnwrapper_8570_io_out_grant_ready;
  assign mem_ic_io_out_0_acquire_ready = NastiIOTileLinkIOConverter_8573_io_tl_acquire_ready;
  assign mem_ic_io_out_0_grant_valid = NastiIOTileLinkIOConverter_8573_io_tl_grant_valid;
  assign mem_ic_io_out_0_grant_bits_addr_beat = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_addr_beat;
  assign mem_ic_io_out_0_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_client_xact_id;
  assign mem_ic_io_out_0_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_manager_xact_id;
  assign mem_ic_io_out_0_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_is_builtin_type;
  assign mem_ic_io_out_0_grant_bits_g_type = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_g_type;
  assign mem_ic_io_out_0_grant_bits_data = NastiIOTileLinkIOConverter_8573_io_tl_grant_bits_data;
  assign ClientTileLinkIOUnwrapper_8570_clk = clk;
  assign ClientTileLinkIOUnwrapper_8570_reset = reset;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_valid = ClientTileLinkEnqueuer_8572_io_outer_acquire_valid;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_block = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_client_xact_id = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_addr_beat = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_is_builtin_type = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_a_type = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_union = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_union;
  assign ClientTileLinkIOUnwrapper_8570_io_in_acquire_bits_data = ClientTileLinkEnqueuer_8572_io_outer_acquire_bits_data;
  assign ClientTileLinkIOUnwrapper_8570_io_in_probe_ready = ClientTileLinkEnqueuer_8572_io_outer_probe_ready;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_valid = ClientTileLinkEnqueuer_8572_io_outer_release_valid;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_beat = ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_addr_block = ClientTileLinkEnqueuer_8572_io_outer_release_bits_addr_block;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_client_xact_id = ClientTileLinkEnqueuer_8572_io_outer_release_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_voluntary = ClientTileLinkEnqueuer_8572_io_outer_release_bits_voluntary;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_r_type = ClientTileLinkEnqueuer_8572_io_outer_release_bits_r_type;
  assign ClientTileLinkIOUnwrapper_8570_io_in_release_bits_data = ClientTileLinkEnqueuer_8572_io_outer_release_bits_data;
  assign ClientTileLinkIOUnwrapper_8570_io_in_grant_ready = ClientTileLinkEnqueuer_8572_io_outer_grant_ready;
  assign ClientTileLinkIOUnwrapper_8570_io_in_finish_valid = ClientTileLinkEnqueuer_8572_io_outer_finish_valid;
  assign ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_xact_id = ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_8570_io_in_finish_bits_manager_id = ClientTileLinkEnqueuer_8572_io_outer_finish_bits_manager_id;
  assign ClientTileLinkIOUnwrapper_8570_io_out_acquire_ready = mem_ic_io_in_0_acquire_ready;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_valid = mem_ic_io_in_0_grant_valid;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_addr_beat = mem_ic_io_in_0_grant_bits_addr_beat;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_client_xact_id = mem_ic_io_in_0_grant_bits_client_xact_id;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_manager_xact_id = mem_ic_io_in_0_grant_bits_manager_xact_id;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_is_builtin_type = mem_ic_io_in_0_grant_bits_is_builtin_type;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_g_type = mem_ic_io_in_0_grant_bits_g_type;
  assign ClientTileLinkIOUnwrapper_8570_io_out_grant_bits_data = mem_ic_io_in_0_grant_bits_data;
  assign ClientTileLinkIOWrapper_8571_clk = clk;
  assign ClientTileLinkIOWrapper_8571_reset = reset;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_valid = L2BroadcastHub_8569_io_outer_acquire_valid;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_block = L2BroadcastHub_8569_io_outer_acquire_bits_addr_block;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_client_xact_id = L2BroadcastHub_8569_io_outer_acquire_bits_client_xact_id;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_addr_beat = L2BroadcastHub_8569_io_outer_acquire_bits_addr_beat;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_is_builtin_type = L2BroadcastHub_8569_io_outer_acquire_bits_is_builtin_type;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_a_type = L2BroadcastHub_8569_io_outer_acquire_bits_a_type;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_union = L2BroadcastHub_8569_io_outer_acquire_bits_union;
  assign ClientTileLinkIOWrapper_8571_io_in_acquire_bits_data = L2BroadcastHub_8569_io_outer_acquire_bits_data;
  assign ClientTileLinkIOWrapper_8571_io_in_grant_ready = L2BroadcastHub_8569_io_outer_grant_ready;
  assign ClientTileLinkIOWrapper_8571_io_out_acquire_ready = ClientTileLinkEnqueuer_8572_io_inner_acquire_ready;
  assign ClientTileLinkIOWrapper_8571_io_out_probe_valid = ClientTileLinkEnqueuer_8572_io_inner_probe_valid;
  assign ClientTileLinkIOWrapper_8571_io_out_probe_bits_addr_block = ClientTileLinkEnqueuer_8572_io_inner_probe_bits_addr_block;
  assign ClientTileLinkIOWrapper_8571_io_out_probe_bits_p_type = ClientTileLinkEnqueuer_8572_io_inner_probe_bits_p_type;
  assign ClientTileLinkIOWrapper_8571_io_out_release_ready = ClientTileLinkEnqueuer_8572_io_inner_release_ready;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_valid = ClientTileLinkEnqueuer_8572_io_inner_grant_valid;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_addr_beat = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_addr_beat;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_client_xact_id = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_client_xact_id;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_xact_id = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_xact_id;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_is_builtin_type = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_is_builtin_type;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_g_type = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_g_type;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_data = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_data;
  assign ClientTileLinkIOWrapper_8571_io_out_grant_bits_manager_id = ClientTileLinkEnqueuer_8572_io_inner_grant_bits_manager_id;
  assign ClientTileLinkIOWrapper_8571_io_out_finish_ready = ClientTileLinkEnqueuer_8572_io_inner_finish_ready;
  assign ClientTileLinkEnqueuer_8572_clk = clk;
  assign ClientTileLinkEnqueuer_8572_reset = reset;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_valid = ClientTileLinkIOWrapper_8571_io_out_acquire_valid;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_block = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_block;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_client_xact_id = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_addr_beat = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_addr_beat;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_is_builtin_type = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_a_type = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_a_type;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_union = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_union;
  assign ClientTileLinkEnqueuer_8572_io_inner_acquire_bits_data = ClientTileLinkIOWrapper_8571_io_out_acquire_bits_data;
  assign ClientTileLinkEnqueuer_8572_io_inner_probe_ready = ClientTileLinkIOWrapper_8571_io_out_probe_ready;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_valid = ClientTileLinkIOWrapper_8571_io_out_release_valid;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_beat = ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_beat;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_addr_block = ClientTileLinkIOWrapper_8571_io_out_release_bits_addr_block;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_client_xact_id = ClientTileLinkIOWrapper_8571_io_out_release_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_voluntary = ClientTileLinkIOWrapper_8571_io_out_release_bits_voluntary;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_r_type = ClientTileLinkIOWrapper_8571_io_out_release_bits_r_type;
  assign ClientTileLinkEnqueuer_8572_io_inner_release_bits_data = ClientTileLinkIOWrapper_8571_io_out_release_bits_data;
  assign ClientTileLinkEnqueuer_8572_io_inner_grant_ready = ClientTileLinkIOWrapper_8571_io_out_grant_ready;
  assign ClientTileLinkEnqueuer_8572_io_inner_finish_valid = ClientTileLinkIOWrapper_8571_io_out_finish_valid;
  assign ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_xact_id = ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_8572_io_inner_finish_bits_manager_id = ClientTileLinkIOWrapper_8571_io_out_finish_bits_manager_id;
  assign ClientTileLinkEnqueuer_8572_io_outer_acquire_ready = ClientTileLinkIOUnwrapper_8570_io_in_acquire_ready;
  assign ClientTileLinkEnqueuer_8572_io_outer_probe_valid = ClientTileLinkIOUnwrapper_8570_io_in_probe_valid;
  assign ClientTileLinkEnqueuer_8572_io_outer_probe_bits_addr_block = ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_addr_block;
  assign ClientTileLinkEnqueuer_8572_io_outer_probe_bits_p_type = ClientTileLinkIOUnwrapper_8570_io_in_probe_bits_p_type;
  assign ClientTileLinkEnqueuer_8572_io_outer_release_ready = ClientTileLinkIOUnwrapper_8570_io_in_release_ready;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_valid = ClientTileLinkIOUnwrapper_8570_io_in_grant_valid;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_addr_beat = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_addr_beat;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_client_xact_id = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_client_xact_id;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_xact_id = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_xact_id;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_is_builtin_type = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_is_builtin_type;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_g_type = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_g_type;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_data = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_data;
  assign ClientTileLinkEnqueuer_8572_io_outer_grant_bits_manager_id = ClientTileLinkIOUnwrapper_8570_io_in_grant_bits_manager_id;
  assign ClientTileLinkEnqueuer_8572_io_outer_finish_ready = ClientTileLinkIOUnwrapper_8570_io_in_finish_ready;
  assign NastiIOTileLinkIOConverter_8573_clk = clk;
  assign NastiIOTileLinkIOConverter_8573_reset = reset;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_valid = mem_ic_io_out_0_acquire_valid;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_block = mem_ic_io_out_0_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_client_xact_id = mem_ic_io_out_0_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_addr_beat = mem_ic_io_out_0_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_is_builtin_type = mem_ic_io_out_0_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_a_type = mem_ic_io_out_0_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_union = mem_ic_io_out_0_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_8573_io_tl_acquire_bits_data = mem_ic_io_out_0_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_8573_io_tl_grant_ready = mem_ic_io_out_0_grant_ready;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_aw_ready = Queue_40_8599_io_enq_ready;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_w_ready = Queue_41_8606_io_enq_ready;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_b_valid = Queue_43_8618_io_deq_valid;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_resp = Queue_43_8618_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_id = Queue_43_8618_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_b_bits_user = Queue_43_8618_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_ar_ready = Queue_39_8586_io_enq_ready;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_valid = Queue_42_8613_io_deq_valid;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_resp = Queue_42_8613_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_data = Queue_42_8613_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_last = Queue_42_8613_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_id = Queue_42_8613_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_8573_io_nasti_r_bits_user = Queue_42_8613_io_deq_bits_user;
  assign Queue_39_8586_clk = clk;
  assign Queue_39_8586_reset = reset;
  assign Queue_39_8586_io_enq_valid = NastiIOTileLinkIOConverter_8573_io_nasti_ar_valid;
  assign Queue_39_8586_io_enq_bits_addr = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_addr;
  assign Queue_39_8586_io_enq_bits_len = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_len;
  assign Queue_39_8586_io_enq_bits_size = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_size;
  assign Queue_39_8586_io_enq_bits_burst = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_burst;
  assign Queue_39_8586_io_enq_bits_lock = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_lock;
  assign Queue_39_8586_io_enq_bits_cache = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_cache;
  assign Queue_39_8586_io_enq_bits_prot = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_prot;
  assign Queue_39_8586_io_enq_bits_qos = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_qos;
  assign Queue_39_8586_io_enq_bits_region = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_region;
  assign Queue_39_8586_io_enq_bits_id = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_id;
  assign Queue_39_8586_io_enq_bits_user = NastiIOTileLinkIOConverter_8573_io_nasti_ar_bits_user;
  assign Queue_39_8586_io_deq_ready = io_mem_axi_0_ar_ready;
  assign Queue_40_8599_clk = clk;
  assign Queue_40_8599_reset = reset;
  assign Queue_40_8599_io_enq_valid = NastiIOTileLinkIOConverter_8573_io_nasti_aw_valid;
  assign Queue_40_8599_io_enq_bits_addr = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_addr;
  assign Queue_40_8599_io_enq_bits_len = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_len;
  assign Queue_40_8599_io_enq_bits_size = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_size;
  assign Queue_40_8599_io_enq_bits_burst = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_burst;
  assign Queue_40_8599_io_enq_bits_lock = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_lock;
  assign Queue_40_8599_io_enq_bits_cache = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_cache;
  assign Queue_40_8599_io_enq_bits_prot = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_prot;
  assign Queue_40_8599_io_enq_bits_qos = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_qos;
  assign Queue_40_8599_io_enq_bits_region = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_region;
  assign Queue_40_8599_io_enq_bits_id = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_id;
  assign Queue_40_8599_io_enq_bits_user = NastiIOTileLinkIOConverter_8573_io_nasti_aw_bits_user;
  assign Queue_40_8599_io_deq_ready = io_mem_axi_0_aw_ready;
  assign Queue_41_8606_clk = clk;
  assign Queue_41_8606_reset = reset;
  assign Queue_41_8606_io_enq_valid = NastiIOTileLinkIOConverter_8573_io_nasti_w_valid;
  assign Queue_41_8606_io_enq_bits_data = NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_data;
  assign Queue_41_8606_io_enq_bits_last = NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_last;
  assign Queue_41_8606_io_enq_bits_id = NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_id;
  assign Queue_41_8606_io_enq_bits_strb = NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_strb;
  assign Queue_41_8606_io_enq_bits_user = NastiIOTileLinkIOConverter_8573_io_nasti_w_bits_user;
  assign Queue_41_8606_io_deq_ready = io_mem_axi_0_w_ready;
  assign Queue_42_8613_clk = clk;
  assign Queue_42_8613_reset = reset;
  assign Queue_42_8613_io_enq_valid = io_mem_axi_0_r_valid;
  assign Queue_42_8613_io_enq_bits_resp = io_mem_axi_0_r_bits_resp;
  assign Queue_42_8613_io_enq_bits_data = io_mem_axi_0_r_bits_data;
  assign Queue_42_8613_io_enq_bits_last = io_mem_axi_0_r_bits_last;
  assign Queue_42_8613_io_enq_bits_id = io_mem_axi_0_r_bits_id;
  assign Queue_42_8613_io_enq_bits_user = io_mem_axi_0_r_bits_user;
  assign Queue_42_8613_io_deq_ready = NastiIOTileLinkIOConverter_8573_io_nasti_r_ready;
  assign Queue_43_8618_clk = clk;
  assign Queue_43_8618_reset = reset;
  assign Queue_43_8618_io_enq_valid = io_mem_axi_0_b_valid;
  assign Queue_43_8618_io_enq_bits_resp = io_mem_axi_0_b_bits_resp;
  assign Queue_43_8618_io_enq_bits_id = io_mem_axi_0_b_bits_id;
  assign Queue_43_8618_io_enq_bits_user = io_mem_axi_0_b_bits_user;
  assign Queue_43_8618_io_deq_ready = NastiIOTileLinkIOConverter_8573_io_nasti_b_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  GEN_0 = GEN_1[0:0];
  end
`endif
endmodule
module SCRFile(
  input   clk,
  input   reset,
  output  io_smi_req_ready,
  input   io_smi_req_valid,
  input   io_smi_req_bits_rw,
  input  [5:0] io_smi_req_bits_addr,
  input  [63:0] io_smi_req_bits_data,
  input   io_smi_resp_ready,
  output  io_smi_resp_valid,
  output [63:0] io_smi_resp_bits,
  input  [63:0] io_scr_rdata_0,
  input  [63:0] io_scr_rdata_1,
  input  [63:0] io_scr_rdata_2,
  input  [63:0] io_scr_rdata_3,
  input  [63:0] io_scr_rdata_4,
  input  [63:0] io_scr_rdata_5,
  input  [63:0] io_scr_rdata_6,
  input  [63:0] io_scr_rdata_7,
  input  [63:0] io_scr_rdata_8,
  input  [63:0] io_scr_rdata_9,
  input  [63:0] io_scr_rdata_10,
  input  [63:0] io_scr_rdata_11,
  input  [63:0] io_scr_rdata_12,
  input  [63:0] io_scr_rdata_13,
  input  [63:0] io_scr_rdata_14,
  input  [63:0] io_scr_rdata_15,
  input  [63:0] io_scr_rdata_16,
  input  [63:0] io_scr_rdata_17,
  input  [63:0] io_scr_rdata_18,
  input  [63:0] io_scr_rdata_19,
  input  [63:0] io_scr_rdata_20,
  input  [63:0] io_scr_rdata_21,
  input  [63:0] io_scr_rdata_22,
  input  [63:0] io_scr_rdata_23,
  input  [63:0] io_scr_rdata_24,
  input  [63:0] io_scr_rdata_25,
  input  [63:0] io_scr_rdata_26,
  input  [63:0] io_scr_rdata_27,
  input  [63:0] io_scr_rdata_28,
  input  [63:0] io_scr_rdata_29,
  input  [63:0] io_scr_rdata_30,
  input  [63:0] io_scr_rdata_31,
  input  [63:0] io_scr_rdata_32,
  input  [63:0] io_scr_rdata_33,
  input  [63:0] io_scr_rdata_34,
  input  [63:0] io_scr_rdata_35,
  input  [63:0] io_scr_rdata_36,
  input  [63:0] io_scr_rdata_37,
  input  [63:0] io_scr_rdata_38,
  input  [63:0] io_scr_rdata_39,
  input  [63:0] io_scr_rdata_40,
  input  [63:0] io_scr_rdata_41,
  input  [63:0] io_scr_rdata_42,
  input  [63:0] io_scr_rdata_43,
  input  [63:0] io_scr_rdata_44,
  input  [63:0] io_scr_rdata_45,
  input  [63:0] io_scr_rdata_46,
  input  [63:0] io_scr_rdata_47,
  input  [63:0] io_scr_rdata_48,
  input  [63:0] io_scr_rdata_49,
  input  [63:0] io_scr_rdata_50,
  input  [63:0] io_scr_rdata_51,
  input  [63:0] io_scr_rdata_52,
  input  [63:0] io_scr_rdata_53,
  input  [63:0] io_scr_rdata_54,
  input  [63:0] io_scr_rdata_55,
  input  [63:0] io_scr_rdata_56,
  input  [63:0] io_scr_rdata_57,
  input  [63:0] io_scr_rdata_58,
  input  [63:0] io_scr_rdata_59,
  input  [63:0] io_scr_rdata_60,
  input  [63:0] io_scr_rdata_61,
  input  [63:0] io_scr_rdata_62,
  input  [63:0] io_scr_rdata_63,
  output  io_scr_wen,
  output [5:0] io_scr_waddr,
  output [63:0] io_scr_wdata
);
  wire [63:0] scr_rdata_0;
  wire [63:0] scr_rdata_1;
  wire [63:0] scr_rdata_2;
  wire [63:0] scr_rdata_3;
  wire [63:0] scr_rdata_4;
  wire [63:0] scr_rdata_5;
  wire [63:0] scr_rdata_6;
  wire [63:0] scr_rdata_7;
  wire [63:0] scr_rdata_8;
  wire [63:0] scr_rdata_9;
  wire [63:0] scr_rdata_10;
  wire [63:0] scr_rdata_11;
  wire [63:0] scr_rdata_12;
  wire [63:0] scr_rdata_13;
  wire [63:0] scr_rdata_14;
  wire [63:0] scr_rdata_15;
  wire [63:0] scr_rdata_16;
  wire [63:0] scr_rdata_17;
  wire [63:0] scr_rdata_18;
  wire [63:0] scr_rdata_19;
  wire [63:0] scr_rdata_20;
  wire [63:0] scr_rdata_21;
  wire [63:0] scr_rdata_22;
  wire [63:0] scr_rdata_23;
  wire [63:0] scr_rdata_24;
  wire [63:0] scr_rdata_25;
  wire [63:0] scr_rdata_26;
  wire [63:0] scr_rdata_27;
  wire [63:0] scr_rdata_28;
  wire [63:0] scr_rdata_29;
  wire [63:0] scr_rdata_30;
  wire [63:0] scr_rdata_31;
  wire [63:0] scr_rdata_32;
  wire [63:0] scr_rdata_33;
  wire [63:0] scr_rdata_34;
  wire [63:0] scr_rdata_35;
  wire [63:0] scr_rdata_36;
  wire [63:0] scr_rdata_37;
  wire [63:0] scr_rdata_38;
  wire [63:0] scr_rdata_39;
  wire [63:0] scr_rdata_40;
  wire [63:0] scr_rdata_41;
  wire [63:0] scr_rdata_42;
  wire [63:0] scr_rdata_43;
  wire [63:0] scr_rdata_44;
  wire [63:0] scr_rdata_45;
  wire [63:0] scr_rdata_46;
  wire [63:0] scr_rdata_47;
  wire [63:0] scr_rdata_48;
  wire [63:0] scr_rdata_49;
  wire [63:0] scr_rdata_50;
  wire [63:0] scr_rdata_51;
  wire [63:0] scr_rdata_52;
  wire [63:0] scr_rdata_53;
  wire [63:0] scr_rdata_54;
  wire [63:0] scr_rdata_55;
  wire [63:0] scr_rdata_56;
  wire [63:0] scr_rdata_57;
  wire [63:0] scr_rdata_58;
  wire [63:0] scr_rdata_59;
  wire [63:0] scr_rdata_60;
  wire [63:0] scr_rdata_61;
  wire [63:0] scr_rdata_62;
  wire [63:0] scr_rdata_63;
  reg [5:0] read_addr;
  reg [31:0] GEN_98;
  reg  resp_valid;
  reg [31:0] GEN_99;
  wire  T_164;
  wire [63:0] GEN_0;
  wire [5:0] GEN_67;
  wire [63:0] GEN_1;
  wire [5:0] GEN_68;
  wire [63:0] GEN_2;
  wire [5:0] GEN_69;
  wire [63:0] GEN_3;
  wire [5:0] GEN_70;
  wire [63:0] GEN_4;
  wire [5:0] GEN_71;
  wire [63:0] GEN_5;
  wire [5:0] GEN_72;
  wire [63:0] GEN_6;
  wire [5:0] GEN_73;
  wire [63:0] GEN_7;
  wire [5:0] GEN_74;
  wire [63:0] GEN_8;
  wire [5:0] GEN_75;
  wire [63:0] GEN_9;
  wire [5:0] GEN_76;
  wire [63:0] GEN_10;
  wire [5:0] GEN_77;
  wire [63:0] GEN_11;
  wire [5:0] GEN_78;
  wire [63:0] GEN_12;
  wire [5:0] GEN_79;
  wire [63:0] GEN_13;
  wire [5:0] GEN_80;
  wire [63:0] GEN_14;
  wire [5:0] GEN_81;
  wire [63:0] GEN_15;
  wire [5:0] GEN_82;
  wire [63:0] GEN_16;
  wire [5:0] GEN_83;
  wire [63:0] GEN_17;
  wire [5:0] GEN_84;
  wire [63:0] GEN_18;
  wire [5:0] GEN_85;
  wire [63:0] GEN_19;
  wire [5:0] GEN_86;
  wire [63:0] GEN_20;
  wire [5:0] GEN_87;
  wire [63:0] GEN_21;
  wire [5:0] GEN_88;
  wire [63:0] GEN_22;
  wire [5:0] GEN_89;
  wire [63:0] GEN_23;
  wire [5:0] GEN_90;
  wire [63:0] GEN_24;
  wire [5:0] GEN_91;
  wire [63:0] GEN_25;
  wire [5:0] GEN_92;
  wire [63:0] GEN_26;
  wire [5:0] GEN_93;
  wire [63:0] GEN_27;
  wire [5:0] GEN_94;
  wire [63:0] GEN_28;
  wire [5:0] GEN_95;
  wire [63:0] GEN_29;
  wire [5:0] GEN_96;
  wire [63:0] GEN_30;
  wire [5:0] GEN_97;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  wire [63:0] GEN_35;
  wire [63:0] GEN_36;
  wire [63:0] GEN_37;
  wire [63:0] GEN_38;
  wire [63:0] GEN_39;
  wire [63:0] GEN_40;
  wire [63:0] GEN_41;
  wire [63:0] GEN_42;
  wire [63:0] GEN_43;
  wire [63:0] GEN_44;
  wire [63:0] GEN_45;
  wire [63:0] GEN_46;
  wire [63:0] GEN_47;
  wire [63:0] GEN_48;
  wire [63:0] GEN_49;
  wire [63:0] GEN_50;
  wire [63:0] GEN_51;
  wire [63:0] GEN_52;
  wire [63:0] GEN_53;
  wire [63:0] GEN_54;
  wire [63:0] GEN_55;
  wire [63:0] GEN_56;
  wire [63:0] GEN_57;
  wire [63:0] GEN_58;
  wire [63:0] GEN_59;
  wire [63:0] GEN_60;
  wire [63:0] GEN_61;
  wire [63:0] GEN_62;
  wire [63:0] GEN_63;
  wire  T_165;
  wire  T_166;
  wire [5:0] GEN_64;
  wire  GEN_65;
  wire  T_169;
  wire  GEN_66;
  assign io_smi_req_ready = T_164;
  assign io_smi_resp_valid = resp_valid;
  assign io_smi_resp_bits = GEN_0;
  assign io_scr_wen = T_166;
  assign io_scr_waddr = io_smi_req_bits_addr;
  assign io_scr_wdata = io_smi_req_bits_data;
  assign scr_rdata_0 = io_scr_rdata_0;
  assign scr_rdata_1 = io_scr_rdata_1;
  assign scr_rdata_2 = io_scr_rdata_2;
  assign scr_rdata_3 = io_scr_rdata_3;
  assign scr_rdata_4 = io_scr_rdata_4;
  assign scr_rdata_5 = io_scr_rdata_5;
  assign scr_rdata_6 = io_scr_rdata_6;
  assign scr_rdata_7 = io_scr_rdata_7;
  assign scr_rdata_8 = io_scr_rdata_8;
  assign scr_rdata_9 = io_scr_rdata_9;
  assign scr_rdata_10 = io_scr_rdata_10;
  assign scr_rdata_11 = io_scr_rdata_11;
  assign scr_rdata_12 = io_scr_rdata_12;
  assign scr_rdata_13 = io_scr_rdata_13;
  assign scr_rdata_14 = io_scr_rdata_14;
  assign scr_rdata_15 = io_scr_rdata_15;
  assign scr_rdata_16 = io_scr_rdata_16;
  assign scr_rdata_17 = io_scr_rdata_17;
  assign scr_rdata_18 = io_scr_rdata_18;
  assign scr_rdata_19 = io_scr_rdata_19;
  assign scr_rdata_20 = io_scr_rdata_20;
  assign scr_rdata_21 = io_scr_rdata_21;
  assign scr_rdata_22 = io_scr_rdata_22;
  assign scr_rdata_23 = io_scr_rdata_23;
  assign scr_rdata_24 = io_scr_rdata_24;
  assign scr_rdata_25 = io_scr_rdata_25;
  assign scr_rdata_26 = io_scr_rdata_26;
  assign scr_rdata_27 = io_scr_rdata_27;
  assign scr_rdata_28 = io_scr_rdata_28;
  assign scr_rdata_29 = io_scr_rdata_29;
  assign scr_rdata_30 = io_scr_rdata_30;
  assign scr_rdata_31 = io_scr_rdata_31;
  assign scr_rdata_32 = io_scr_rdata_32;
  assign scr_rdata_33 = io_scr_rdata_33;
  assign scr_rdata_34 = io_scr_rdata_34;
  assign scr_rdata_35 = io_scr_rdata_35;
  assign scr_rdata_36 = io_scr_rdata_36;
  assign scr_rdata_37 = io_scr_rdata_37;
  assign scr_rdata_38 = io_scr_rdata_38;
  assign scr_rdata_39 = io_scr_rdata_39;
  assign scr_rdata_40 = io_scr_rdata_40;
  assign scr_rdata_41 = io_scr_rdata_41;
  assign scr_rdata_42 = io_scr_rdata_42;
  assign scr_rdata_43 = io_scr_rdata_43;
  assign scr_rdata_44 = io_scr_rdata_44;
  assign scr_rdata_45 = io_scr_rdata_45;
  assign scr_rdata_46 = io_scr_rdata_46;
  assign scr_rdata_47 = io_scr_rdata_47;
  assign scr_rdata_48 = io_scr_rdata_48;
  assign scr_rdata_49 = io_scr_rdata_49;
  assign scr_rdata_50 = io_scr_rdata_50;
  assign scr_rdata_51 = io_scr_rdata_51;
  assign scr_rdata_52 = io_scr_rdata_52;
  assign scr_rdata_53 = io_scr_rdata_53;
  assign scr_rdata_54 = io_scr_rdata_54;
  assign scr_rdata_55 = io_scr_rdata_55;
  assign scr_rdata_56 = io_scr_rdata_56;
  assign scr_rdata_57 = io_scr_rdata_57;
  assign scr_rdata_58 = io_scr_rdata_58;
  assign scr_rdata_59 = io_scr_rdata_59;
  assign scr_rdata_60 = io_scr_rdata_60;
  assign scr_rdata_61 = io_scr_rdata_61;
  assign scr_rdata_62 = io_scr_rdata_62;
  assign scr_rdata_63 = io_scr_rdata_63;
  assign T_164 = resp_valid == 1'h0;
  assign GEN_0 = GEN_63;
  assign GEN_67 = {{5'd0}, 1'h1};
  assign GEN_1 = GEN_67 == read_addr ? scr_rdata_1 : scr_rdata_0;
  assign GEN_68 = {{4'd0}, 2'h2};
  assign GEN_2 = GEN_68 == read_addr ? scr_rdata_2 : GEN_1;
  assign GEN_69 = {{4'd0}, 2'h3};
  assign GEN_3 = GEN_69 == read_addr ? scr_rdata_3 : GEN_2;
  assign GEN_70 = {{3'd0}, 3'h4};
  assign GEN_4 = GEN_70 == read_addr ? scr_rdata_4 : GEN_3;
  assign GEN_71 = {{3'd0}, 3'h5};
  assign GEN_5 = GEN_71 == read_addr ? scr_rdata_5 : GEN_4;
  assign GEN_72 = {{3'd0}, 3'h6};
  assign GEN_6 = GEN_72 == read_addr ? scr_rdata_6 : GEN_5;
  assign GEN_73 = {{3'd0}, 3'h7};
  assign GEN_7 = GEN_73 == read_addr ? scr_rdata_7 : GEN_6;
  assign GEN_74 = {{2'd0}, 4'h8};
  assign GEN_8 = GEN_74 == read_addr ? scr_rdata_8 : GEN_7;
  assign GEN_75 = {{2'd0}, 4'h9};
  assign GEN_9 = GEN_75 == read_addr ? scr_rdata_9 : GEN_8;
  assign GEN_76 = {{2'd0}, 4'ha};
  assign GEN_10 = GEN_76 == read_addr ? scr_rdata_10 : GEN_9;
  assign GEN_77 = {{2'd0}, 4'hb};
  assign GEN_11 = GEN_77 == read_addr ? scr_rdata_11 : GEN_10;
  assign GEN_78 = {{2'd0}, 4'hc};
  assign GEN_12 = GEN_78 == read_addr ? scr_rdata_12 : GEN_11;
  assign GEN_79 = {{2'd0}, 4'hd};
  assign GEN_13 = GEN_79 == read_addr ? scr_rdata_13 : GEN_12;
  assign GEN_80 = {{2'd0}, 4'he};
  assign GEN_14 = GEN_80 == read_addr ? scr_rdata_14 : GEN_13;
  assign GEN_81 = {{2'd0}, 4'hf};
  assign GEN_15 = GEN_81 == read_addr ? scr_rdata_15 : GEN_14;
  assign GEN_82 = {{1'd0}, 5'h10};
  assign GEN_16 = GEN_82 == read_addr ? scr_rdata_16 : GEN_15;
  assign GEN_83 = {{1'd0}, 5'h11};
  assign GEN_17 = GEN_83 == read_addr ? scr_rdata_17 : GEN_16;
  assign GEN_84 = {{1'd0}, 5'h12};
  assign GEN_18 = GEN_84 == read_addr ? scr_rdata_18 : GEN_17;
  assign GEN_85 = {{1'd0}, 5'h13};
  assign GEN_19 = GEN_85 == read_addr ? scr_rdata_19 : GEN_18;
  assign GEN_86 = {{1'd0}, 5'h14};
  assign GEN_20 = GEN_86 == read_addr ? scr_rdata_20 : GEN_19;
  assign GEN_87 = {{1'd0}, 5'h15};
  assign GEN_21 = GEN_87 == read_addr ? scr_rdata_21 : GEN_20;
  assign GEN_88 = {{1'd0}, 5'h16};
  assign GEN_22 = GEN_88 == read_addr ? scr_rdata_22 : GEN_21;
  assign GEN_89 = {{1'd0}, 5'h17};
  assign GEN_23 = GEN_89 == read_addr ? scr_rdata_23 : GEN_22;
  assign GEN_90 = {{1'd0}, 5'h18};
  assign GEN_24 = GEN_90 == read_addr ? scr_rdata_24 : GEN_23;
  assign GEN_91 = {{1'd0}, 5'h19};
  assign GEN_25 = GEN_91 == read_addr ? scr_rdata_25 : GEN_24;
  assign GEN_92 = {{1'd0}, 5'h1a};
  assign GEN_26 = GEN_92 == read_addr ? scr_rdata_26 : GEN_25;
  assign GEN_93 = {{1'd0}, 5'h1b};
  assign GEN_27 = GEN_93 == read_addr ? scr_rdata_27 : GEN_26;
  assign GEN_94 = {{1'd0}, 5'h1c};
  assign GEN_28 = GEN_94 == read_addr ? scr_rdata_28 : GEN_27;
  assign GEN_95 = {{1'd0}, 5'h1d};
  assign GEN_29 = GEN_95 == read_addr ? scr_rdata_29 : GEN_28;
  assign GEN_96 = {{1'd0}, 5'h1e};
  assign GEN_30 = GEN_96 == read_addr ? scr_rdata_30 : GEN_29;
  assign GEN_97 = {{1'd0}, 5'h1f};
  assign GEN_31 = GEN_97 == read_addr ? scr_rdata_31 : GEN_30;
  assign GEN_32 = 6'h20 == read_addr ? scr_rdata_32 : GEN_31;
  assign GEN_33 = 6'h21 == read_addr ? scr_rdata_33 : GEN_32;
  assign GEN_34 = 6'h22 == read_addr ? scr_rdata_34 : GEN_33;
  assign GEN_35 = 6'h23 == read_addr ? scr_rdata_35 : GEN_34;
  assign GEN_36 = 6'h24 == read_addr ? scr_rdata_36 : GEN_35;
  assign GEN_37 = 6'h25 == read_addr ? scr_rdata_37 : GEN_36;
  assign GEN_38 = 6'h26 == read_addr ? scr_rdata_38 : GEN_37;
  assign GEN_39 = 6'h27 == read_addr ? scr_rdata_39 : GEN_38;
  assign GEN_40 = 6'h28 == read_addr ? scr_rdata_40 : GEN_39;
  assign GEN_41 = 6'h29 == read_addr ? scr_rdata_41 : GEN_40;
  assign GEN_42 = 6'h2a == read_addr ? scr_rdata_42 : GEN_41;
  assign GEN_43 = 6'h2b == read_addr ? scr_rdata_43 : GEN_42;
  assign GEN_44 = 6'h2c == read_addr ? scr_rdata_44 : GEN_43;
  assign GEN_45 = 6'h2d == read_addr ? scr_rdata_45 : GEN_44;
  assign GEN_46 = 6'h2e == read_addr ? scr_rdata_46 : GEN_45;
  assign GEN_47 = 6'h2f == read_addr ? scr_rdata_47 : GEN_46;
  assign GEN_48 = 6'h30 == read_addr ? scr_rdata_48 : GEN_47;
  assign GEN_49 = 6'h31 == read_addr ? scr_rdata_49 : GEN_48;
  assign GEN_50 = 6'h32 == read_addr ? scr_rdata_50 : GEN_49;
  assign GEN_51 = 6'h33 == read_addr ? scr_rdata_51 : GEN_50;
  assign GEN_52 = 6'h34 == read_addr ? scr_rdata_52 : GEN_51;
  assign GEN_53 = 6'h35 == read_addr ? scr_rdata_53 : GEN_52;
  assign GEN_54 = 6'h36 == read_addr ? scr_rdata_54 : GEN_53;
  assign GEN_55 = 6'h37 == read_addr ? scr_rdata_55 : GEN_54;
  assign GEN_56 = 6'h38 == read_addr ? scr_rdata_56 : GEN_55;
  assign GEN_57 = 6'h39 == read_addr ? scr_rdata_57 : GEN_56;
  assign GEN_58 = 6'h3a == read_addr ? scr_rdata_58 : GEN_57;
  assign GEN_59 = 6'h3b == read_addr ? scr_rdata_59 : GEN_58;
  assign GEN_60 = 6'h3c == read_addr ? scr_rdata_60 : GEN_59;
  assign GEN_61 = 6'h3d == read_addr ? scr_rdata_61 : GEN_60;
  assign GEN_62 = 6'h3e == read_addr ? scr_rdata_62 : GEN_61;
  assign GEN_63 = 6'h3f == read_addr ? scr_rdata_63 : GEN_62;
  assign T_165 = io_smi_req_ready & io_smi_req_valid;
  assign T_166 = T_165 & io_smi_req_bits_rw;
  assign GEN_64 = T_165 ? io_smi_req_bits_addr : read_addr;
  assign GEN_65 = T_165 ? 1'h1 : resp_valid;
  assign T_169 = io_smi_resp_ready & io_smi_resp_valid;
  assign GEN_66 = T_169 ? 1'h0 : GEN_65;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_98 = {1{$random}};
  read_addr = GEN_98[5:0];
  GEN_99 = {1{$random}};
  resp_valid = GEN_99[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      read_addr <= 6'h0;
    end else begin
      read_addr <= GEN_64;
    end
    if(reset) begin
      resp_valid <= 1'h0;
    end else begin
      resp_valid <= GEN_66;
    end
  end
endmodule
module LockingRRArbiter_44(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [1:0] GEN_2;
  wire [1:0] GEN_9;
  wire  GEN_3;
  wire  GEN_10;
  wire  GEN_4;
  wire  GEN_11;
  wire [3:0] GEN_5;
  wire [3:0] GEN_12;
  wire [63:0] GEN_6;
  wire [63:0] GEN_13;
  reg [2:0] T_610;
  reg [31:0] GEN_24;
  reg  T_612;
  reg [31:0] GEN_25;
  wire [2:0] GEN_20;
  wire  T_614;
  wire [2:0] T_622_0;
  wire [3:0] GEN_21;
  wire  T_624;
  wire  T_632_0;
  wire [3:0] GEN_22;
  wire  T_634;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire [2:0] GEN_23;
  wire [3:0] T_644;
  wire [2:0] T_645;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  reg  lastGrant;
  reg [31:0] GEN_26;
  wire  GEN_17;
  wire  T_650;
  wire  T_652;
  wire  T_655;
  wire  T_659;
  wire  T_661;
  wire  T_665;
  wire  T_667;
  wire  T_668;
  wire  T_669;
  wire  T_672;
  wire  T_673;
  wire  GEN_18;
  wire  GEN_19;
  assign io_in_0_ready = T_669;
  assign io_in_1_ready = T_673;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_16;
  assign choice = GEN_19;
  assign GEN_0 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_3 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_4 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_5 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_6 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_20 = {{2'd0}, 1'h0};
  assign T_614 = T_610 != GEN_20;
  assign T_622_0 = 3'h5;
  assign GEN_21 = {{1'd0}, T_622_0};
  assign T_624 = GEN_21 == io_out_bits_g_type;
  assign T_632_0 = 1'h0;
  assign GEN_22 = {{3'd0}, T_632_0};
  assign T_634 = GEN_22 == io_out_bits_g_type;
  assign T_637 = io_out_bits_is_builtin_type ? T_624 : T_634;
  assign T_639 = io_out_ready & io_out_valid;
  assign T_640 = T_639 & T_637;
  assign GEN_23 = {{2'd0}, 1'h1};
  assign T_644 = T_610 + GEN_23;
  assign T_645 = T_644[2:0];
  assign GEN_14 = T_640 ? io_chosen : T_612;
  assign GEN_15 = T_640 ? T_645 : T_610;
  assign GEN_16 = T_614 ? T_612 : choice;
  assign GEN_17 = T_639 ? io_chosen : lastGrant;
  assign T_650 = 1'h1 > lastGrant;
  assign T_652 = io_in_1_valid & T_650;
  assign T_655 = T_652 | io_in_0_valid;
  assign T_659 = T_652 == 1'h0;
  assign T_661 = T_655 == 1'h0;
  assign T_665 = T_650 | T_661;
  assign T_667 = T_612 == 1'h0;
  assign T_668 = T_614 ? T_667 : T_659;
  assign T_669 = T_668 & io_out_ready;
  assign T_672 = T_614 ? T_612 : T_665;
  assign T_673 = T_672 & io_out_ready;
  assign GEN_18 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_19 = T_652 ? 1'h1 : GEN_18;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_24 = {1{$random}};
  T_610 = GEN_24[2:0];
  GEN_25 = {1{$random}};
  T_612 = GEN_25[0:0];
  GEN_26 = {1{$random}};
  lastGrant = GEN_26[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_610 <= 3'h0;
    end else begin
      T_610 <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_612 <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_17;
    end
  end
endmodule
module ClientUncachedTileLinkIORouter(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire [2:0] T_1442;
  wire [28:0] T_1443;
  wire [31:0] T_1444;
  wire [31:0] GEN_2;
  wire  T_1448;
  wire [31:0] GEN_3;
  wire  T_1451;
  wire  T_1453;
  wire  T_1454;
  wire [1:0] acq_route;
  wire  T_1456;
  wire  T_1457;
  wire  GEN_0;
  wire  T_1459;
  wire  T_1460;
  wire  GEN_1;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_chosen;
  wire  T_1485;
  wire [1:0] GEN_4;
  wire  T_1487;
  wire  T_1488;
  wire  T_1489;
  wire  T_1491;
  LockingRRArbiter_44 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_1;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_1457;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_1460;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign T_1442 = io_in_acquire_bits_union[11:9];
  assign T_1443 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_1444 = {T_1443,T_1442};
  assign GEN_2 = {{1'd0}, 31'h48000000};
  assign T_1448 = T_1444 < GEN_2;
  assign GEN_3 = {{1'd0}, 31'h60000000};
  assign T_1451 = GEN_3 <= T_1444;
  assign T_1453 = T_1444 < 32'h80000000;
  assign T_1454 = T_1451 & T_1453;
  assign acq_route = {T_1454,T_1448};
  assign T_1456 = acq_route[0];
  assign T_1457 = io_in_acquire_valid & T_1456;
  assign GEN_0 = T_1456 ? io_out_0_acquire_ready : 1'h0;
  assign T_1459 = acq_route[1];
  assign T_1460 = io_in_acquire_valid & T_1459;
  assign GEN_1 = T_1459 ? io_out_1_acquire_ready : GEN_0;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_1485 = io_in_acquire_valid == 1'h0;
  assign GEN_4 = {{1'd0}, 1'h0};
  assign T_1487 = acq_route != GEN_4;
  assign T_1488 = T_1485 | T_1487;
  assign T_1489 = T_1488 | reset;
  assign T_1491 = T_1489 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1491) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at interconnect.scala:218 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1491) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_2666_clk;
  wire  ClientUncachedTileLinkIORouter_2666_reset;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_data;
  ClientUncachedTileLinkIORouter ClientUncachedTileLinkIORouter_2666 (
    .clk(ClientUncachedTileLinkIORouter_2666_clk),
    .reset(ClientUncachedTileLinkIORouter_2666_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_2666_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_2666_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_2666_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_2666_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_2666_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_2666_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_2666_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_2666_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_2666_io_out_1_grant_ready;
  assign ClientUncachedTileLinkIORouter_2666_clk = clk;
  assign ClientUncachedTileLinkIORouter_2666_reset = reset;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_2666_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_2666_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_2666_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_2666_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
endmodule
module LockingRRArbiter_48(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_addr_beat,
  input  [1:0] io_in_2_bits_client_xact_id,
  input   io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_is_builtin_type,
  input  [3:0] io_in_2_bits_g_type,
  input  [63:0] io_in_2_bits_data,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [2:0] io_in_3_bits_addr_beat,
  input  [1:0] io_in_3_bits_client_xact_id,
  input   io_in_3_bits_manager_xact_id,
  input   io_in_3_bits_is_builtin_type,
  input  [3:0] io_in_3_bits_g_type,
  input  [63:0] io_in_3_bits_data,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [2:0] io_in_4_bits_addr_beat,
  input  [1:0] io_in_4_bits_client_xact_id,
  input   io_in_4_bits_manager_xact_id,
  input   io_in_4_bits_is_builtin_type,
  input  [3:0] io_in_4_bits_g_type,
  input  [63:0] io_in_4_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output [2:0] io_chosen
);
  wire [2:0] choice;
  wire  GEN_0;
  wire [2:0] GEN_47;
  wire  GEN_7;
  wire [2:0] GEN_48;
  wire  GEN_8;
  wire [2:0] GEN_49;
  wire  GEN_9;
  wire  GEN_10;
  wire [2:0] GEN_1;
  wire [2:0] GEN_11;
  wire [2:0] GEN_12;
  wire [2:0] GEN_13;
  wire [2:0] GEN_14;
  wire [1:0] GEN_2;
  wire [1:0] GEN_15;
  wire [1:0] GEN_16;
  wire [1:0] GEN_17;
  wire [1:0] GEN_18;
  wire  GEN_3;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_4;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [3:0] GEN_5;
  wire [3:0] GEN_27;
  wire [3:0] GEN_28;
  wire [3:0] GEN_29;
  wire [3:0] GEN_30;
  wire [63:0] GEN_6;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [63:0] GEN_33;
  wire [63:0] GEN_34;
  reg [2:0] T_886;
  reg [31:0] GEN_50;
  reg [2:0] T_888;
  reg [31:0] GEN_51;
  wire [2:0] GEN_68;
  wire  T_890;
  wire [2:0] T_898_0;
  wire [3:0] GEN_69;
  wire  T_900;
  wire  T_908_0;
  wire [3:0] GEN_70;
  wire  T_910;
  wire  T_913;
  wire  T_915;
  wire  T_916;
  wire [3:0] T_920;
  wire [2:0] T_921;
  wire [2:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  reg [2:0] lastGrant;
  reg [31:0] GEN_52;
  wire [2:0] GEN_38;
  wire  T_926;
  wire  T_928;
  wire  T_930;
  wire  T_932;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_950;
  wire  T_952;
  wire  T_954;
  wire  T_956;
  wire  T_958;
  wire  T_960;
  wire  T_962;
  wire  T_964;
  wire  T_968;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire  T_976;
  wire  T_977;
  wire  T_978;
  wire  T_980;
  wire  T_981;
  wire  T_982;
  wire  T_984;
  wire  T_985;
  wire  T_986;
  wire  T_988;
  wire  T_989;
  wire  T_990;
  wire  T_992;
  wire  T_993;
  wire  T_994;
  wire [2:0] GEN_39;
  wire [2:0] GEN_40;
  wire [2:0] GEN_41;
  wire [2:0] GEN_42;
  wire [2:0] GEN_43;
  wire [2:0] GEN_44;
  wire [2:0] GEN_45;
  wire [2:0] GEN_46;
  assign io_in_0_ready = T_978;
  assign io_in_1_ready = T_982;
  assign io_in_2_ready = T_986;
  assign io_in_3_ready = T_990;
  assign io_in_4_ready = T_994;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_37;
  assign choice = GEN_46;
  assign GEN_0 = GEN_10;
  assign GEN_47 = {{2'd0}, 1'h1};
  assign GEN_7 = GEN_47 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_48 = {{1'd0}, 2'h2};
  assign GEN_8 = GEN_48 == io_chosen ? io_in_2_valid : GEN_7;
  assign GEN_49 = {{1'd0}, 2'h3};
  assign GEN_9 = GEN_49 == io_chosen ? io_in_3_valid : GEN_8;
  assign GEN_10 = 3'h4 == io_chosen ? io_in_4_valid : GEN_9;
  assign GEN_1 = GEN_14;
  assign GEN_11 = GEN_47 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_12 = GEN_48 == io_chosen ? io_in_2_bits_addr_beat : GEN_11;
  assign GEN_13 = GEN_49 == io_chosen ? io_in_3_bits_addr_beat : GEN_12;
  assign GEN_14 = 3'h4 == io_chosen ? io_in_4_bits_addr_beat : GEN_13;
  assign GEN_2 = GEN_18;
  assign GEN_15 = GEN_47 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_16 = GEN_48 == io_chosen ? io_in_2_bits_client_xact_id : GEN_15;
  assign GEN_17 = GEN_49 == io_chosen ? io_in_3_bits_client_xact_id : GEN_16;
  assign GEN_18 = 3'h4 == io_chosen ? io_in_4_bits_client_xact_id : GEN_17;
  assign GEN_3 = GEN_22;
  assign GEN_19 = GEN_47 == io_chosen ? io_in_1_bits_manager_xact_id : io_in_0_bits_manager_xact_id;
  assign GEN_20 = GEN_48 == io_chosen ? io_in_2_bits_manager_xact_id : GEN_19;
  assign GEN_21 = GEN_49 == io_chosen ? io_in_3_bits_manager_xact_id : GEN_20;
  assign GEN_22 = 3'h4 == io_chosen ? io_in_4_bits_manager_xact_id : GEN_21;
  assign GEN_4 = GEN_26;
  assign GEN_23 = GEN_47 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_24 = GEN_48 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_23;
  assign GEN_25 = GEN_49 == io_chosen ? io_in_3_bits_is_builtin_type : GEN_24;
  assign GEN_26 = 3'h4 == io_chosen ? io_in_4_bits_is_builtin_type : GEN_25;
  assign GEN_5 = GEN_30;
  assign GEN_27 = GEN_47 == io_chosen ? io_in_1_bits_g_type : io_in_0_bits_g_type;
  assign GEN_28 = GEN_48 == io_chosen ? io_in_2_bits_g_type : GEN_27;
  assign GEN_29 = GEN_49 == io_chosen ? io_in_3_bits_g_type : GEN_28;
  assign GEN_30 = 3'h4 == io_chosen ? io_in_4_bits_g_type : GEN_29;
  assign GEN_6 = GEN_34;
  assign GEN_31 = GEN_47 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_32 = GEN_48 == io_chosen ? io_in_2_bits_data : GEN_31;
  assign GEN_33 = GEN_49 == io_chosen ? io_in_3_bits_data : GEN_32;
  assign GEN_34 = 3'h4 == io_chosen ? io_in_4_bits_data : GEN_33;
  assign GEN_68 = {{2'd0}, 1'h0};
  assign T_890 = T_886 != GEN_68;
  assign T_898_0 = 3'h5;
  assign GEN_69 = {{1'd0}, T_898_0};
  assign T_900 = GEN_69 == io_out_bits_g_type;
  assign T_908_0 = 1'h0;
  assign GEN_70 = {{3'd0}, T_908_0};
  assign T_910 = GEN_70 == io_out_bits_g_type;
  assign T_913 = io_out_bits_is_builtin_type ? T_900 : T_910;
  assign T_915 = io_out_ready & io_out_valid;
  assign T_916 = T_915 & T_913;
  assign T_920 = T_886 + GEN_47;
  assign T_921 = T_920[2:0];
  assign GEN_35 = T_916 ? io_chosen : T_888;
  assign GEN_36 = T_916 ? T_921 : T_886;
  assign GEN_37 = T_890 ? T_888 : choice;
  assign GEN_38 = T_915 ? io_chosen : lastGrant;
  assign T_926 = GEN_47 > lastGrant;
  assign T_928 = GEN_48 > lastGrant;
  assign T_930 = GEN_49 > lastGrant;
  assign T_932 = 3'h4 > lastGrant;
  assign T_934 = io_in_1_valid & T_926;
  assign T_935 = io_in_2_valid & T_928;
  assign T_936 = io_in_3_valid & T_930;
  assign T_937 = io_in_4_valid & T_932;
  assign T_940 = T_934 | T_935;
  assign T_941 = T_940 | T_936;
  assign T_942 = T_941 | T_937;
  assign T_943 = T_942 | io_in_0_valid;
  assign T_944 = T_943 | io_in_1_valid;
  assign T_945 = T_944 | io_in_2_valid;
  assign T_946 = T_945 | io_in_3_valid;
  assign T_950 = T_934 == 1'h0;
  assign T_952 = T_940 == 1'h0;
  assign T_954 = T_941 == 1'h0;
  assign T_956 = T_942 == 1'h0;
  assign T_958 = T_943 == 1'h0;
  assign T_960 = T_944 == 1'h0;
  assign T_962 = T_945 == 1'h0;
  assign T_964 = T_946 == 1'h0;
  assign T_968 = T_926 | T_958;
  assign T_969 = T_950 & T_928;
  assign T_970 = T_969 | T_960;
  assign T_971 = T_952 & T_930;
  assign T_972 = T_971 | T_962;
  assign T_973 = T_954 & T_932;
  assign T_974 = T_973 | T_964;
  assign T_976 = T_888 == GEN_68;
  assign T_977 = T_890 ? T_976 : T_956;
  assign T_978 = T_977 & io_out_ready;
  assign T_980 = T_888 == GEN_47;
  assign T_981 = T_890 ? T_980 : T_968;
  assign T_982 = T_981 & io_out_ready;
  assign T_984 = T_888 == GEN_48;
  assign T_985 = T_890 ? T_984 : T_970;
  assign T_986 = T_985 & io_out_ready;
  assign T_988 = T_888 == GEN_49;
  assign T_989 = T_890 ? T_988 : T_972;
  assign T_990 = T_989 & io_out_ready;
  assign T_992 = T_888 == 3'h4;
  assign T_993 = T_890 ? T_992 : T_974;
  assign T_994 = T_993 & io_out_ready;
  assign GEN_39 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_40 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_39;
  assign GEN_41 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_40;
  assign GEN_42 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_41;
  assign GEN_43 = T_937 ? 3'h4 : GEN_42;
  assign GEN_44 = T_936 ? {{1'd0}, 2'h3} : GEN_43;
  assign GEN_45 = T_935 ? {{1'd0}, 2'h2} : GEN_44;
  assign GEN_46 = T_934 ? {{2'd0}, 1'h1} : GEN_45;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_50 = {1{$random}};
  T_886 = GEN_50[2:0];
  GEN_51 = {1{$random}};
  T_888 = GEN_51[2:0];
  GEN_52 = {1{$random}};
  lastGrant = GEN_52[2:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_886 <= 3'h0;
    end else begin
      T_886 <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      T_888 <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      lastGrant <= GEN_38;
    end
  end
endmodule
module ClientUncachedTileLinkIORouter_47(
  input   clk,
  input   reset,
  output  io_in_acquire_ready,
  input   io_in_acquire_valid,
  input  [25:0] io_in_acquire_bits_addr_block,
  input  [1:0] io_in_acquire_bits_client_xact_id,
  input  [2:0] io_in_acquire_bits_addr_beat,
  input   io_in_acquire_bits_is_builtin_type,
  input  [2:0] io_in_acquire_bits_a_type,
  input  [11:0] io_in_acquire_bits_union,
  input  [63:0] io_in_acquire_bits_data,
  input   io_in_grant_ready,
  output  io_in_grant_valid,
  output [2:0] io_in_grant_bits_addr_beat,
  output [1:0] io_in_grant_bits_client_xact_id,
  output  io_in_grant_bits_manager_xact_id,
  output  io_in_grant_bits_is_builtin_type,
  output [3:0] io_in_grant_bits_g_type,
  output [63:0] io_in_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire [2:0] T_2051;
  wire [28:0] T_2052;
  wire [31:0] T_2053;
  wire [31:0] GEN_5;
  wire  T_2057;
  wire  T_2060;
  wire [31:0] GEN_7;
  wire  T_2062;
  wire  T_2063;
  wire  T_2065;
  wire [31:0] GEN_9;
  wire  T_2067;
  wire  T_2068;
  wire [31:0] GEN_10;
  wire  T_2070;
  wire [31:0] GEN_11;
  wire  T_2072;
  wire  T_2073;
  wire  T_2075;
  wire [31:0] GEN_13;
  wire  T_2077;
  wire  T_2078;
  wire [1:0] T_2079;
  wire [1:0] T_2080;
  wire [2:0] T_2081;
  wire [4:0] acq_route;
  wire  T_2083;
  wire  T_2084;
  wire  GEN_0;
  wire  T_2086;
  wire  T_2087;
  wire  GEN_1;
  wire  T_2089;
  wire  T_2090;
  wire  GEN_2;
  wire  T_2092;
  wire  T_2093;
  wire  GEN_3;
  wire  T_2095;
  wire  T_2096;
  wire  GEN_4;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_2_ready;
  wire  gnt_arb_io_in_2_valid;
  wire [2:0] gnt_arb_io_in_2_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_2_bits_client_xact_id;
  wire  gnt_arb_io_in_2_bits_manager_xact_id;
  wire  gnt_arb_io_in_2_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_2_bits_g_type;
  wire [63:0] gnt_arb_io_in_2_bits_data;
  wire  gnt_arb_io_in_3_ready;
  wire  gnt_arb_io_in_3_valid;
  wire [2:0] gnt_arb_io_in_3_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_3_bits_client_xact_id;
  wire  gnt_arb_io_in_3_bits_manager_xact_id;
  wire  gnt_arb_io_in_3_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_3_bits_g_type;
  wire [63:0] gnt_arb_io_in_3_bits_data;
  wire  gnt_arb_io_in_4_ready;
  wire  gnt_arb_io_in_4_valid;
  wire [2:0] gnt_arb_io_in_4_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_4_bits_client_xact_id;
  wire  gnt_arb_io_in_4_bits_manager_xact_id;
  wire  gnt_arb_io_in_4_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_4_bits_g_type;
  wire [63:0] gnt_arb_io_in_4_bits_data;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire [2:0] gnt_arb_io_chosen;
  wire  T_2121;
  wire [4:0] GEN_14;
  wire  T_2123;
  wire  T_2124;
  wire  T_2125;
  wire  T_2127;
  LockingRRArbiter_48 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_2_ready(gnt_arb_io_in_2_ready),
    .io_in_2_valid(gnt_arb_io_in_2_valid),
    .io_in_2_bits_addr_beat(gnt_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_client_xact_id(gnt_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_manager_xact_id(gnt_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_is_builtin_type(gnt_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_g_type(gnt_arb_io_in_2_bits_g_type),
    .io_in_2_bits_data(gnt_arb_io_in_2_bits_data),
    .io_in_3_ready(gnt_arb_io_in_3_ready),
    .io_in_3_valid(gnt_arb_io_in_3_valid),
    .io_in_3_bits_addr_beat(gnt_arb_io_in_3_bits_addr_beat),
    .io_in_3_bits_client_xact_id(gnt_arb_io_in_3_bits_client_xact_id),
    .io_in_3_bits_manager_xact_id(gnt_arb_io_in_3_bits_manager_xact_id),
    .io_in_3_bits_is_builtin_type(gnt_arb_io_in_3_bits_is_builtin_type),
    .io_in_3_bits_g_type(gnt_arb_io_in_3_bits_g_type),
    .io_in_3_bits_data(gnt_arb_io_in_3_bits_data),
    .io_in_4_ready(gnt_arb_io_in_4_ready),
    .io_in_4_valid(gnt_arb_io_in_4_valid),
    .io_in_4_bits_addr_beat(gnt_arb_io_in_4_bits_addr_beat),
    .io_in_4_bits_client_xact_id(gnt_arb_io_in_4_bits_client_xact_id),
    .io_in_4_bits_manager_xact_id(gnt_arb_io_in_4_bits_manager_xact_id),
    .io_in_4_bits_is_builtin_type(gnt_arb_io_in_4_bits_is_builtin_type),
    .io_in_4_bits_g_type(gnt_arb_io_in_4_bits_g_type),
    .io_in_4_bits_data(gnt_arb_io_in_4_bits_data),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_in_acquire_ready = GEN_4;
  assign io_in_grant_valid = gnt_arb_io_out_valid;
  assign io_in_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_in_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_in_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_in_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_in_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_in_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_out_0_acquire_valid = T_2084;
  assign io_out_0_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_0_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_0_grant_ready = gnt_arb_io_in_0_ready;
  assign io_out_1_acquire_valid = T_2087;
  assign io_out_1_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_1_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_1_grant_ready = gnt_arb_io_in_1_ready;
  assign io_out_2_acquire_valid = T_2090;
  assign io_out_2_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_2_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_2_grant_ready = gnt_arb_io_in_2_ready;
  assign io_out_3_acquire_valid = T_2093;
  assign io_out_3_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_3_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_3_grant_ready = gnt_arb_io_in_3_ready;
  assign io_out_4_acquire_valid = T_2096;
  assign io_out_4_acquire_bits_addr_block = io_in_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = io_in_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = io_in_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = io_in_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = io_in_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = io_in_acquire_bits_union;
  assign io_out_4_acquire_bits_data = io_in_acquire_bits_data;
  assign io_out_4_grant_ready = gnt_arb_io_in_4_ready;
  assign T_2051 = io_in_acquire_bits_union[11:9];
  assign T_2052 = {io_in_acquire_bits_addr_block,io_in_acquire_bits_addr_beat};
  assign T_2053 = {T_2052,T_2051};
  assign GEN_5 = {{19'd0}, 13'h1000};
  assign T_2057 = T_2053 < GEN_5;
  assign T_2060 = GEN_5 <= T_2053;
  assign GEN_7 = {{18'd0}, 14'h2000};
  assign T_2062 = T_2053 < GEN_7;
  assign T_2063 = T_2060 & T_2062;
  assign T_2065 = GEN_7 <= T_2053;
  assign GEN_9 = {{18'd0}, 14'h3000};
  assign T_2067 = T_2053 < GEN_9;
  assign T_2068 = T_2065 & T_2067;
  assign GEN_10 = {{1'd0}, 31'h40000000};
  assign T_2070 = GEN_10 <= T_2053;
  assign GEN_11 = {{1'd0}, 31'h44000000};
  assign T_2072 = T_2053 < GEN_11;
  assign T_2073 = T_2070 & T_2072;
  assign T_2075 = GEN_11 <= T_2053;
  assign GEN_13 = {{1'd0}, 31'h48000000};
  assign T_2077 = T_2053 < GEN_13;
  assign T_2078 = T_2075 & T_2077;
  assign T_2079 = {T_2063,T_2057};
  assign T_2080 = {T_2078,T_2073};
  assign T_2081 = {T_2080,T_2068};
  assign acq_route = {T_2081,T_2079};
  assign T_2083 = acq_route[0];
  assign T_2084 = io_in_acquire_valid & T_2083;
  assign GEN_0 = T_2083 ? io_out_0_acquire_ready : 1'h0;
  assign T_2086 = acq_route[1];
  assign T_2087 = io_in_acquire_valid & T_2086;
  assign GEN_1 = T_2086 ? io_out_1_acquire_ready : GEN_0;
  assign T_2089 = acq_route[2];
  assign T_2090 = io_in_acquire_valid & T_2089;
  assign GEN_2 = T_2089 ? io_out_2_acquire_ready : GEN_1;
  assign T_2092 = acq_route[3];
  assign T_2093 = io_in_acquire_valid & T_2092;
  assign GEN_3 = T_2092 ? io_out_3_acquire_ready : GEN_2;
  assign T_2095 = acq_route[4];
  assign T_2096 = io_in_acquire_valid & T_2095;
  assign GEN_4 = T_2095 ? io_out_4_acquire_ready : GEN_3;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_out_0_grant_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = io_out_0_grant_bits_g_type;
  assign gnt_arb_io_in_0_bits_data = io_out_0_grant_bits_data;
  assign gnt_arb_io_in_1_valid = io_out_1_grant_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = io_out_1_grant_bits_g_type;
  assign gnt_arb_io_in_1_bits_data = io_out_1_grant_bits_data;
  assign gnt_arb_io_in_2_valid = io_out_2_grant_valid;
  assign gnt_arb_io_in_2_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign gnt_arb_io_in_2_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign gnt_arb_io_in_2_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_2_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_2_bits_g_type = io_out_2_grant_bits_g_type;
  assign gnt_arb_io_in_2_bits_data = io_out_2_grant_bits_data;
  assign gnt_arb_io_in_3_valid = io_out_3_grant_valid;
  assign gnt_arb_io_in_3_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign gnt_arb_io_in_3_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign gnt_arb_io_in_3_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_3_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_3_bits_g_type = io_out_3_grant_bits_g_type;
  assign gnt_arb_io_in_3_bits_data = io_out_3_grant_bits_data;
  assign gnt_arb_io_in_4_valid = io_out_4_grant_valid;
  assign gnt_arb_io_in_4_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign gnt_arb_io_in_4_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign gnt_arb_io_in_4_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign gnt_arb_io_in_4_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign gnt_arb_io_in_4_bits_g_type = io_out_4_grant_bits_g_type;
  assign gnt_arb_io_in_4_bits_data = io_out_4_grant_bits_data;
  assign gnt_arb_io_out_ready = io_in_grant_ready;
  assign T_2121 = io_in_acquire_valid == 1'h0;
  assign GEN_14 = {{4'd0}, 1'h0};
  assign T_2123 = acq_route != GEN_14;
  assign T_2124 = T_2121 | T_2123;
  assign T_2125 = T_2124 | reset;
  assign T_2127 = T_2125 == 1'h0;
  always @(posedge clk) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2127) begin
          $fwrite(32'h80000002,"Assertion failed: No valid route\n    at interconnect.scala:218 assert(!io.in.acquire.valid || acq_route.orR, \"No valid route\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2127) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module ClientUncachedTileLinkIOCrossbar_46(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire  ClientUncachedTileLinkIORouter_47_3275_clk;
  wire  ClientUncachedTileLinkIORouter_47_3275_reset;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_valid;
  wire [25:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_block;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_beat;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_a_type;
  wire [11:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_union;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_data;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_ready;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_valid;
  wire [2:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_addr_beat;
  wire [1:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_client_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_manager_xact_id;
  wire  ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_g_type;
  wire [63:0] ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIORouter_47 ClientUncachedTileLinkIORouter_47_3275 (
    .clk(ClientUncachedTileLinkIORouter_47_3275_clk),
    .reset(ClientUncachedTileLinkIORouter_47_3275_reset),
    .io_in_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_ready),
    .io_in_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_valid),
    .io_in_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_block),
    .io_in_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_client_xact_id),
    .io_in_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_beat),
    .io_in_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_is_builtin_type),
    .io_in_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_a_type),
    .io_in_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_union),
    .io_in_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_data),
    .io_in_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_ready),
    .io_in_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_valid),
    .io_in_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_addr_beat),
    .io_in_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_client_xact_id),
    .io_in_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_manager_xact_id),
    .io_in_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_is_builtin_type),
    .io_in_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_g_type),
    .io_in_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_data),
    .io_out_0_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_ready),
    .io_out_0_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_ready),
    .io_out_1_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_ready),
    .io_out_2_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_ready),
    .io_out_3_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_ready),
    .io_out_4_grant_valid(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_ready;
  assign io_in_0_grant_valid = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_valid;
  assign io_in_0_grant_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_g_type;
  assign io_in_0_grant_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_in_grant_bits_data;
  assign io_out_0_acquire_valid = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_clk = clk;
  assign ClientUncachedTileLinkIORouter_47_3275_reset = reset;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_valid = io_in_0_acquire_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_union = io_in_0_acquire_bits_union;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_acquire_bits_data = io_in_0_acquire_bits_data;
  assign ClientUncachedTileLinkIORouter_47_3275_io_in_grant_ready = io_in_0_grant_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_valid = io_out_0_grant_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_valid = io_out_1_grant_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_valid = io_out_2_grant_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_valid = io_out_3_grant_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_valid = io_out_4_grant_valid;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign ClientUncachedTileLinkIORouter_47_3275_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect_45(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  xbar_io_out_2_acquire_ready;
  wire  xbar_io_out_2_acquire_valid;
  wire [25:0] xbar_io_out_2_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_2_acquire_bits_addr_beat;
  wire  xbar_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_2_acquire_bits_a_type;
  wire [11:0] xbar_io_out_2_acquire_bits_union;
  wire [63:0] xbar_io_out_2_acquire_bits_data;
  wire  xbar_io_out_2_grant_ready;
  wire  xbar_io_out_2_grant_valid;
  wire [2:0] xbar_io_out_2_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_2_grant_bits_client_xact_id;
  wire  xbar_io_out_2_grant_bits_manager_xact_id;
  wire  xbar_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_2_grant_bits_g_type;
  wire [63:0] xbar_io_out_2_grant_bits_data;
  wire  xbar_io_out_3_acquire_ready;
  wire  xbar_io_out_3_acquire_valid;
  wire [25:0] xbar_io_out_3_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_3_acquire_bits_addr_beat;
  wire  xbar_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_3_acquire_bits_a_type;
  wire [11:0] xbar_io_out_3_acquire_bits_union;
  wire [63:0] xbar_io_out_3_acquire_bits_data;
  wire  xbar_io_out_3_grant_ready;
  wire  xbar_io_out_3_grant_valid;
  wire [2:0] xbar_io_out_3_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_3_grant_bits_client_xact_id;
  wire  xbar_io_out_3_grant_bits_manager_xact_id;
  wire  xbar_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_3_grant_bits_g_type;
  wire [63:0] xbar_io_out_3_grant_bits_data;
  wire  xbar_io_out_4_acquire_ready;
  wire  xbar_io_out_4_acquire_valid;
  wire [25:0] xbar_io_out_4_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_4_acquire_bits_addr_beat;
  wire  xbar_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_4_acquire_bits_a_type;
  wire [11:0] xbar_io_out_4_acquire_bits_union;
  wire [63:0] xbar_io_out_4_acquire_bits_data;
  wire  xbar_io_out_4_grant_ready;
  wire  xbar_io_out_4_grant_valid;
  wire [2:0] xbar_io_out_4_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_4_grant_bits_client_xact_id;
  wire  xbar_io_out_4_grant_bits_manager_xact_id;
  wire  xbar_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_4_grant_bits_g_type;
  wire [63:0] xbar_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar_46 xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(xbar_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(xbar_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(xbar_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(xbar_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(xbar_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(xbar_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(xbar_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(xbar_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(xbar_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(xbar_io_out_2_grant_ready),
    .io_out_2_grant_valid(xbar_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(xbar_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(xbar_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(xbar_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(xbar_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(xbar_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(xbar_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(xbar_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(xbar_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(xbar_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(xbar_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(xbar_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(xbar_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(xbar_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(xbar_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(xbar_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(xbar_io_out_3_grant_ready),
    .io_out_3_grant_valid(xbar_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(xbar_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(xbar_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(xbar_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(xbar_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(xbar_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(xbar_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(xbar_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(xbar_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(xbar_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(xbar_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(xbar_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(xbar_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(xbar_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(xbar_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(xbar_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(xbar_io_out_4_grant_ready),
    .io_out_4_grant_valid(xbar_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(xbar_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(xbar_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(xbar_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(xbar_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(xbar_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(xbar_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = xbar_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = xbar_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = xbar_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = xbar_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = xbar_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = xbar_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = xbar_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = xbar_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = xbar_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = xbar_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = xbar_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = xbar_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = xbar_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = xbar_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = xbar_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = xbar_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = xbar_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = xbar_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = xbar_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = xbar_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = xbar_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = xbar_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = xbar_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = xbar_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = xbar_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = xbar_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = xbar_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = xbar_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = xbar_io_out_4_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = io_out_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_1_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign xbar_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign xbar_io_out_2_grant_valid = io_out_2_grant_valid;
  assign xbar_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign xbar_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign xbar_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign xbar_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign xbar_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign xbar_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign xbar_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign xbar_io_out_3_grant_valid = io_out_3_grant_valid;
  assign xbar_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign xbar_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign xbar_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign xbar_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign xbar_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign xbar_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign xbar_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign xbar_io_out_4_grant_valid = io_out_4_grant_valid;
  assign xbar_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign xbar_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign xbar_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign xbar_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign xbar_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign xbar_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module TileLinkRecursiveInterconnect(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output  io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_0_acquire_ready,
  output  io_out_0_acquire_valid,
  output [25:0] io_out_0_acquire_bits_addr_block,
  output [1:0] io_out_0_acquire_bits_client_xact_id,
  output [2:0] io_out_0_acquire_bits_addr_beat,
  output  io_out_0_acquire_bits_is_builtin_type,
  output [2:0] io_out_0_acquire_bits_a_type,
  output [11:0] io_out_0_acquire_bits_union,
  output [63:0] io_out_0_acquire_bits_data,
  output  io_out_0_grant_ready,
  input   io_out_0_grant_valid,
  input  [2:0] io_out_0_grant_bits_addr_beat,
  input  [1:0] io_out_0_grant_bits_client_xact_id,
  input   io_out_0_grant_bits_manager_xact_id,
  input   io_out_0_grant_bits_is_builtin_type,
  input  [3:0] io_out_0_grant_bits_g_type,
  input  [63:0] io_out_0_grant_bits_data,
  input   io_out_1_acquire_ready,
  output  io_out_1_acquire_valid,
  output [25:0] io_out_1_acquire_bits_addr_block,
  output [1:0] io_out_1_acquire_bits_client_xact_id,
  output [2:0] io_out_1_acquire_bits_addr_beat,
  output  io_out_1_acquire_bits_is_builtin_type,
  output [2:0] io_out_1_acquire_bits_a_type,
  output [11:0] io_out_1_acquire_bits_union,
  output [63:0] io_out_1_acquire_bits_data,
  output  io_out_1_grant_ready,
  input   io_out_1_grant_valid,
  input  [2:0] io_out_1_grant_bits_addr_beat,
  input  [1:0] io_out_1_grant_bits_client_xact_id,
  input   io_out_1_grant_bits_manager_xact_id,
  input   io_out_1_grant_bits_is_builtin_type,
  input  [3:0] io_out_1_grant_bits_g_type,
  input  [63:0] io_out_1_grant_bits_data,
  input   io_out_2_acquire_ready,
  output  io_out_2_acquire_valid,
  output [25:0] io_out_2_acquire_bits_addr_block,
  output [1:0] io_out_2_acquire_bits_client_xact_id,
  output [2:0] io_out_2_acquire_bits_addr_beat,
  output  io_out_2_acquire_bits_is_builtin_type,
  output [2:0] io_out_2_acquire_bits_a_type,
  output [11:0] io_out_2_acquire_bits_union,
  output [63:0] io_out_2_acquire_bits_data,
  output  io_out_2_grant_ready,
  input   io_out_2_grant_valid,
  input  [2:0] io_out_2_grant_bits_addr_beat,
  input  [1:0] io_out_2_grant_bits_client_xact_id,
  input   io_out_2_grant_bits_manager_xact_id,
  input   io_out_2_grant_bits_is_builtin_type,
  input  [3:0] io_out_2_grant_bits_g_type,
  input  [63:0] io_out_2_grant_bits_data,
  input   io_out_3_acquire_ready,
  output  io_out_3_acquire_valid,
  output [25:0] io_out_3_acquire_bits_addr_block,
  output [1:0] io_out_3_acquire_bits_client_xact_id,
  output [2:0] io_out_3_acquire_bits_addr_beat,
  output  io_out_3_acquire_bits_is_builtin_type,
  output [2:0] io_out_3_acquire_bits_a_type,
  output [11:0] io_out_3_acquire_bits_union,
  output [63:0] io_out_3_acquire_bits_data,
  output  io_out_3_grant_ready,
  input   io_out_3_grant_valid,
  input  [2:0] io_out_3_grant_bits_addr_beat,
  input  [1:0] io_out_3_grant_bits_client_xact_id,
  input   io_out_3_grant_bits_manager_xact_id,
  input   io_out_3_grant_bits_is_builtin_type,
  input  [3:0] io_out_3_grant_bits_g_type,
  input  [63:0] io_out_3_grant_bits_data,
  input   io_out_4_acquire_ready,
  output  io_out_4_acquire_valid,
  output [25:0] io_out_4_acquire_bits_addr_block,
  output [1:0] io_out_4_acquire_bits_client_xact_id,
  output [2:0] io_out_4_acquire_bits_addr_beat,
  output  io_out_4_acquire_bits_is_builtin_type,
  output [2:0] io_out_4_acquire_bits_a_type,
  output [11:0] io_out_4_acquire_bits_union,
  output [63:0] io_out_4_acquire_bits_data,
  output  io_out_4_grant_ready,
  input   io_out_4_grant_valid,
  input  [2:0] io_out_4_grant_bits_addr_beat,
  input  [1:0] io_out_4_grant_bits_client_xact_id,
  input   io_out_4_grant_bits_manager_xact_id,
  input   io_out_4_grant_bits_is_builtin_type,
  input  [3:0] io_out_4_grant_bits_g_type,
  input  [63:0] io_out_4_grant_bits_data,
  input   io_out_5_acquire_ready,
  output  io_out_5_acquire_valid,
  output [25:0] io_out_5_acquire_bits_addr_block,
  output [1:0] io_out_5_acquire_bits_client_xact_id,
  output [2:0] io_out_5_acquire_bits_addr_beat,
  output  io_out_5_acquire_bits_is_builtin_type,
  output [2:0] io_out_5_acquire_bits_a_type,
  output [11:0] io_out_5_acquire_bits_union,
  output [63:0] io_out_5_acquire_bits_data,
  output  io_out_5_grant_ready,
  input   io_out_5_grant_valid,
  input  [2:0] io_out_5_grant_bits_addr_beat,
  input  [1:0] io_out_5_grant_bits_client_xact_id,
  input   io_out_5_grant_bits_manager_xact_id,
  input   io_out_5_grant_bits_is_builtin_type,
  input  [3:0] io_out_5_grant_bits_g_type,
  input  [63:0] io_out_5_grant_bits_data
);
  wire  xbar_clk;
  wire  xbar_reset;
  wire  xbar_io_in_0_acquire_ready;
  wire  xbar_io_in_0_acquire_valid;
  wire [25:0] xbar_io_in_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_in_0_acquire_bits_addr_beat;
  wire  xbar_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_in_0_acquire_bits_a_type;
  wire [11:0] xbar_io_in_0_acquire_bits_union;
  wire [63:0] xbar_io_in_0_acquire_bits_data;
  wire  xbar_io_in_0_grant_ready;
  wire  xbar_io_in_0_grant_valid;
  wire [2:0] xbar_io_in_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_in_0_grant_bits_client_xact_id;
  wire  xbar_io_in_0_grant_bits_manager_xact_id;
  wire  xbar_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_in_0_grant_bits_g_type;
  wire [63:0] xbar_io_in_0_grant_bits_data;
  wire  xbar_io_out_0_acquire_ready;
  wire  xbar_io_out_0_acquire_valid;
  wire [25:0] xbar_io_out_0_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_0_acquire_bits_addr_beat;
  wire  xbar_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_0_acquire_bits_a_type;
  wire [11:0] xbar_io_out_0_acquire_bits_union;
  wire [63:0] xbar_io_out_0_acquire_bits_data;
  wire  xbar_io_out_0_grant_ready;
  wire  xbar_io_out_0_grant_valid;
  wire [2:0] xbar_io_out_0_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_0_grant_bits_client_xact_id;
  wire  xbar_io_out_0_grant_bits_manager_xact_id;
  wire  xbar_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_0_grant_bits_g_type;
  wire [63:0] xbar_io_out_0_grant_bits_data;
  wire  xbar_io_out_1_acquire_ready;
  wire  xbar_io_out_1_acquire_valid;
  wire [25:0] xbar_io_out_1_acquire_bits_addr_block;
  wire [1:0] xbar_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] xbar_io_out_1_acquire_bits_addr_beat;
  wire  xbar_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] xbar_io_out_1_acquire_bits_a_type;
  wire [11:0] xbar_io_out_1_acquire_bits_union;
  wire [63:0] xbar_io_out_1_acquire_bits_data;
  wire  xbar_io_out_1_grant_ready;
  wire  xbar_io_out_1_grant_valid;
  wire [2:0] xbar_io_out_1_grant_bits_addr_beat;
  wire [1:0] xbar_io_out_1_grant_bits_client_xact_id;
  wire  xbar_io_out_1_grant_bits_manager_xact_id;
  wire  xbar_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] xbar_io_out_1_grant_bits_g_type;
  wire [63:0] xbar_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_clk;
  wire  TileLinkRecursiveInterconnect_45_3478_reset;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_ready;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_data;
  ClientUncachedTileLinkIOCrossbar xbar (
    .clk(xbar_clk),
    .reset(xbar_reset),
    .io_in_0_acquire_ready(xbar_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(xbar_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(xbar_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(xbar_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(xbar_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(xbar_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(xbar_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(xbar_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(xbar_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(xbar_io_in_0_grant_ready),
    .io_in_0_grant_valid(xbar_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(xbar_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(xbar_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(xbar_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(xbar_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(xbar_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(xbar_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(xbar_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(xbar_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(xbar_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(xbar_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(xbar_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(xbar_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(xbar_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(xbar_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(xbar_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(xbar_io_out_0_grant_ready),
    .io_out_0_grant_valid(xbar_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(xbar_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(xbar_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(xbar_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(xbar_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(xbar_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(xbar_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(xbar_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(xbar_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(xbar_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(xbar_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(xbar_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(xbar_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(xbar_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(xbar_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(xbar_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(xbar_io_out_1_grant_ready),
    .io_out_1_grant_valid(xbar_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(xbar_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(xbar_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(xbar_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(xbar_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(xbar_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(xbar_io_out_1_grant_bits_data)
  );
  TileLinkRecursiveInterconnect_45 TileLinkRecursiveInterconnect_45_3478 (
    .clk(TileLinkRecursiveInterconnect_45_3478_clk),
    .reset(TileLinkRecursiveInterconnect_45_3478_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_ready),
    .io_out_4_grant_valid(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_data)
  );
  assign io_in_0_acquire_ready = xbar_io_in_0_acquire_ready;
  assign io_in_0_grant_valid = xbar_io_in_0_grant_valid;
  assign io_in_0_grant_bits_addr_beat = xbar_io_in_0_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = xbar_io_in_0_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = xbar_io_in_0_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = xbar_io_in_0_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = xbar_io_in_0_grant_bits_g_type;
  assign io_in_0_grant_bits_data = xbar_io_in_0_grant_bits_data;
  assign io_out_0_acquire_valid = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_valid;
  assign io_out_0_acquire_bits_addr_block = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_block;
  assign io_out_0_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_client_xact_id;
  assign io_out_0_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_addr_beat;
  assign io_out_0_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_is_builtin_type;
  assign io_out_0_acquire_bits_a_type = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_a_type;
  assign io_out_0_acquire_bits_union = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_union;
  assign io_out_0_acquire_bits_data = TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_bits_data;
  assign io_out_0_grant_ready = TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_ready;
  assign io_out_1_acquire_valid = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_valid;
  assign io_out_1_acquire_bits_addr_block = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_block;
  assign io_out_1_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_client_xact_id;
  assign io_out_1_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_addr_beat;
  assign io_out_1_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_1_acquire_bits_a_type = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_a_type;
  assign io_out_1_acquire_bits_union = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_union;
  assign io_out_1_acquire_bits_data = TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_bits_data;
  assign io_out_1_grant_ready = TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_ready;
  assign io_out_2_acquire_valid = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_valid;
  assign io_out_2_acquire_bits_addr_block = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_block;
  assign io_out_2_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_client_xact_id;
  assign io_out_2_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_addr_beat;
  assign io_out_2_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_is_builtin_type;
  assign io_out_2_acquire_bits_a_type = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_a_type;
  assign io_out_2_acquire_bits_union = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_union;
  assign io_out_2_acquire_bits_data = TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_bits_data;
  assign io_out_2_grant_ready = TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_ready;
  assign io_out_3_acquire_valid = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_valid;
  assign io_out_3_acquire_bits_addr_block = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_block;
  assign io_out_3_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_client_xact_id;
  assign io_out_3_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_addr_beat;
  assign io_out_3_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_is_builtin_type;
  assign io_out_3_acquire_bits_a_type = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_a_type;
  assign io_out_3_acquire_bits_union = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_union;
  assign io_out_3_acquire_bits_data = TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_bits_data;
  assign io_out_3_grant_ready = TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_ready;
  assign io_out_4_acquire_valid = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_valid;
  assign io_out_4_acquire_bits_addr_block = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_block;
  assign io_out_4_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_client_xact_id;
  assign io_out_4_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_addr_beat;
  assign io_out_4_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_is_builtin_type;
  assign io_out_4_acquire_bits_a_type = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_a_type;
  assign io_out_4_acquire_bits_union = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_union;
  assign io_out_4_acquire_bits_data = TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_bits_data;
  assign io_out_4_grant_ready = TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_ready;
  assign io_out_5_acquire_valid = xbar_io_out_1_acquire_valid;
  assign io_out_5_acquire_bits_addr_block = xbar_io_out_1_acquire_bits_addr_block;
  assign io_out_5_acquire_bits_client_xact_id = xbar_io_out_1_acquire_bits_client_xact_id;
  assign io_out_5_acquire_bits_addr_beat = xbar_io_out_1_acquire_bits_addr_beat;
  assign io_out_5_acquire_bits_is_builtin_type = xbar_io_out_1_acquire_bits_is_builtin_type;
  assign io_out_5_acquire_bits_a_type = xbar_io_out_1_acquire_bits_a_type;
  assign io_out_5_acquire_bits_union = xbar_io_out_1_acquire_bits_union;
  assign io_out_5_acquire_bits_data = xbar_io_out_1_acquire_bits_data;
  assign io_out_5_grant_ready = xbar_io_out_1_grant_ready;
  assign xbar_clk = clk;
  assign xbar_reset = reset;
  assign xbar_io_in_0_acquire_valid = io_in_0_acquire_valid;
  assign xbar_io_in_0_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign xbar_io_in_0_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign xbar_io_in_0_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign xbar_io_in_0_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign xbar_io_in_0_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign xbar_io_in_0_acquire_bits_union = io_in_0_acquire_bits_union;
  assign xbar_io_in_0_acquire_bits_data = io_in_0_acquire_bits_data;
  assign xbar_io_in_0_grant_ready = io_in_0_grant_ready;
  assign xbar_io_out_0_acquire_ready = TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_ready;
  assign xbar_io_out_0_grant_valid = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_valid;
  assign xbar_io_out_0_grant_bits_addr_beat = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_addr_beat;
  assign xbar_io_out_0_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_client_xact_id;
  assign xbar_io_out_0_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_manager_xact_id;
  assign xbar_io_out_0_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_is_builtin_type;
  assign xbar_io_out_0_grant_bits_g_type = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_g_type;
  assign xbar_io_out_0_grant_bits_data = TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_bits_data;
  assign xbar_io_out_1_acquire_ready = io_out_5_acquire_ready;
  assign xbar_io_out_1_grant_valid = io_out_5_grant_valid;
  assign xbar_io_out_1_grant_bits_addr_beat = io_out_5_grant_bits_addr_beat;
  assign xbar_io_out_1_grant_bits_client_xact_id = io_out_5_grant_bits_client_xact_id;
  assign xbar_io_out_1_grant_bits_manager_xact_id = io_out_5_grant_bits_manager_xact_id;
  assign xbar_io_out_1_grant_bits_is_builtin_type = io_out_5_grant_bits_is_builtin_type;
  assign xbar_io_out_1_grant_bits_g_type = io_out_5_grant_bits_g_type;
  assign xbar_io_out_1_grant_bits_data = io_out_5_grant_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_clk = clk;
  assign TileLinkRecursiveInterconnect_45_3478_reset = reset;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_valid = xbar_io_out_0_acquire_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_block = xbar_io_out_0_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_client_xact_id = xbar_io_out_0_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_addr_beat = xbar_io_out_0_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_is_builtin_type = xbar_io_out_0_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_a_type = xbar_io_out_0_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_union = xbar_io_out_0_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_acquire_bits_data = xbar_io_out_0_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_io_in_0_grant_ready = xbar_io_out_0_grant_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_acquire_ready = io_out_0_acquire_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_valid = io_out_0_grant_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_addr_beat = io_out_0_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_client_xact_id = io_out_0_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_manager_xact_id = io_out_0_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_is_builtin_type = io_out_0_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_g_type = io_out_0_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_0_grant_bits_data = io_out_0_grant_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_acquire_ready = io_out_1_acquire_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_valid = io_out_1_grant_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_addr_beat = io_out_1_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_client_xact_id = io_out_1_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_manager_xact_id = io_out_1_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_is_builtin_type = io_out_1_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_g_type = io_out_1_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_1_grant_bits_data = io_out_1_grant_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_acquire_ready = io_out_2_acquire_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_valid = io_out_2_grant_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_addr_beat = io_out_2_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_client_xact_id = io_out_2_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_manager_xact_id = io_out_2_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_is_builtin_type = io_out_2_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_g_type = io_out_2_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_2_grant_bits_data = io_out_2_grant_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_acquire_ready = io_out_3_acquire_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_valid = io_out_3_grant_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_addr_beat = io_out_3_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_client_xact_id = io_out_3_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_manager_xact_id = io_out_3_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_is_builtin_type = io_out_3_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_g_type = io_out_3_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_3_grant_bits_data = io_out_3_grant_bits_data;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_acquire_ready = io_out_4_acquire_ready;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_valid = io_out_4_grant_valid;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_addr_beat = io_out_4_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_client_xact_id = io_out_4_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_manager_xact_id = io_out_4_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_is_builtin_type = io_out_4_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_g_type = io_out_4_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_45_3478_io_out_4_grant_bits_data = io_out_4_grant_bits_data;
endmodule
module Queue_49(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [25:0] io_enq_bits_addr_block,
  input  [1:0] io_enq_bits_client_xact_id,
  input  [2:0] io_enq_bits_addr_beat,
  input   io_enq_bits_is_builtin_type,
  input  [2:0] io_enq_bits_a_type,
  input  [11:0] io_enq_bits_union,
  input  [63:0] io_enq_bits_data,
  input   io_deq_ready,
  output  io_deq_valid,
  output [25:0] io_deq_bits_addr_block,
  output [1:0] io_deq_bits_client_xact_id,
  output [2:0] io_deq_bits_addr_beat,
  output  io_deq_bits_is_builtin_type,
  output [2:0] io_deq_bits_a_type,
  output [11:0] io_deq_bits_union,
  output [63:0] io_deq_bits_data,
  output  io_count
);
  reg [25:0] ram_addr_block [0:0];
  reg [31:0] GEN_0;
  wire [25:0] ram_addr_block_T_254_data;
  wire  ram_addr_block_T_254_addr;
  wire  ram_addr_block_T_254_en;
  wire [25:0] ram_addr_block_T_224_data;
  wire  ram_addr_block_T_224_addr;
  wire  ram_addr_block_T_224_mask;
  wire  ram_addr_block_T_224_en;
  reg [1:0] ram_client_xact_id [0:0];
  reg [31:0] GEN_1;
  wire [1:0] ram_client_xact_id_T_254_data;
  wire  ram_client_xact_id_T_254_addr;
  wire  ram_client_xact_id_T_254_en;
  wire [1:0] ram_client_xact_id_T_224_data;
  wire  ram_client_xact_id_T_224_addr;
  wire  ram_client_xact_id_T_224_mask;
  wire  ram_client_xact_id_T_224_en;
  reg [2:0] ram_addr_beat [0:0];
  reg [31:0] GEN_2;
  wire [2:0] ram_addr_beat_T_254_data;
  wire  ram_addr_beat_T_254_addr;
  wire  ram_addr_beat_T_254_en;
  wire [2:0] ram_addr_beat_T_224_data;
  wire  ram_addr_beat_T_224_addr;
  wire  ram_addr_beat_T_224_mask;
  wire  ram_addr_beat_T_224_en;
  reg  ram_is_builtin_type [0:0];
  reg [31:0] GEN_3;
  wire  ram_is_builtin_type_T_254_data;
  wire  ram_is_builtin_type_T_254_addr;
  wire  ram_is_builtin_type_T_254_en;
  wire  ram_is_builtin_type_T_224_data;
  wire  ram_is_builtin_type_T_224_addr;
  wire  ram_is_builtin_type_T_224_mask;
  wire  ram_is_builtin_type_T_224_en;
  reg [2:0] ram_a_type [0:0];
  reg [31:0] GEN_4;
  wire [2:0] ram_a_type_T_254_data;
  wire  ram_a_type_T_254_addr;
  wire  ram_a_type_T_254_en;
  wire [2:0] ram_a_type_T_224_data;
  wire  ram_a_type_T_224_addr;
  wire  ram_a_type_T_224_mask;
  wire  ram_a_type_T_224_en;
  reg [11:0] ram_union [0:0];
  reg [31:0] GEN_5;
  wire [11:0] ram_union_T_254_data;
  wire  ram_union_T_254_addr;
  wire  ram_union_T_254_en;
  wire [11:0] ram_union_T_224_data;
  wire  ram_union_T_224_addr;
  wire  ram_union_T_224_mask;
  wire  ram_union_T_224_en;
  reg [63:0] ram_data [0:0];
  reg [63:0] GEN_6;
  wire [63:0] ram_data_T_254_data;
  wire  ram_data_T_254_addr;
  wire  ram_data_T_254_en;
  wire [63:0] ram_data_T_224_data;
  wire  ram_data_T_224_addr;
  wire  ram_data_T_224_mask;
  wire  ram_data_T_224_en;
  reg  maybe_full;
  reg [31:0] GEN_7;
  wire  T_221;
  wire  T_222;
  wire  do_enq;
  wire  T_223;
  wire  do_deq;
  wire  T_249;
  wire  GEN_17;
  wire  T_251;
  wire [1:0] T_277;
  wire  ptr_diff;
  wire [1:0] T_279;
  assign io_enq_ready = T_221;
  assign io_deq_valid = T_251;
  assign io_deq_bits_addr_block = ram_addr_block_T_254_data;
  assign io_deq_bits_client_xact_id = ram_client_xact_id_T_254_data;
  assign io_deq_bits_addr_beat = ram_addr_beat_T_254_data;
  assign io_deq_bits_is_builtin_type = ram_is_builtin_type_T_254_data;
  assign io_deq_bits_a_type = ram_a_type_T_254_data;
  assign io_deq_bits_union = ram_union_T_254_data;
  assign io_deq_bits_data = ram_data_T_254_data;
  assign io_count = T_279[0];
  assign ram_addr_block_T_254_addr = 1'h0;
  assign ram_addr_block_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_block_T_254_data = ram_addr_block[ram_addr_block_T_254_addr];
  `else
  assign ram_addr_block_T_254_data = ram_addr_block_T_254_addr >= 1'h1 ? $random : ram_addr_block[ram_addr_block_T_254_addr];
  `endif
  assign ram_addr_block_T_224_data = io_enq_bits_addr_block;
  assign ram_addr_block_T_224_addr = 1'h0;
  assign ram_addr_block_T_224_mask = do_enq;
  assign ram_addr_block_T_224_en = do_enq;
  assign ram_client_xact_id_T_254_addr = 1'h0;
  assign ram_client_xact_id_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_client_xact_id_T_254_data = ram_client_xact_id[ram_client_xact_id_T_254_addr];
  `else
  assign ram_client_xact_id_T_254_data = ram_client_xact_id_T_254_addr >= 1'h1 ? $random : ram_client_xact_id[ram_client_xact_id_T_254_addr];
  `endif
  assign ram_client_xact_id_T_224_data = io_enq_bits_client_xact_id;
  assign ram_client_xact_id_T_224_addr = 1'h0;
  assign ram_client_xact_id_T_224_mask = do_enq;
  assign ram_client_xact_id_T_224_en = do_enq;
  assign ram_addr_beat_T_254_addr = 1'h0;
  assign ram_addr_beat_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_beat_T_254_data = ram_addr_beat[ram_addr_beat_T_254_addr];
  `else
  assign ram_addr_beat_T_254_data = ram_addr_beat_T_254_addr >= 1'h1 ? $random : ram_addr_beat[ram_addr_beat_T_254_addr];
  `endif
  assign ram_addr_beat_T_224_data = io_enq_bits_addr_beat;
  assign ram_addr_beat_T_224_addr = 1'h0;
  assign ram_addr_beat_T_224_mask = do_enq;
  assign ram_addr_beat_T_224_en = do_enq;
  assign ram_is_builtin_type_T_254_addr = 1'h0;
  assign ram_is_builtin_type_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  `else
  assign ram_is_builtin_type_T_254_data = ram_is_builtin_type_T_254_addr >= 1'h1 ? $random : ram_is_builtin_type[ram_is_builtin_type_T_254_addr];
  `endif
  assign ram_is_builtin_type_T_224_data = io_enq_bits_is_builtin_type;
  assign ram_is_builtin_type_T_224_addr = 1'h0;
  assign ram_is_builtin_type_T_224_mask = do_enq;
  assign ram_is_builtin_type_T_224_en = do_enq;
  assign ram_a_type_T_254_addr = 1'h0;
  assign ram_a_type_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_a_type_T_254_data = ram_a_type[ram_a_type_T_254_addr];
  `else
  assign ram_a_type_T_254_data = ram_a_type_T_254_addr >= 1'h1 ? $random : ram_a_type[ram_a_type_T_254_addr];
  `endif
  assign ram_a_type_T_224_data = io_enq_bits_a_type;
  assign ram_a_type_T_224_addr = 1'h0;
  assign ram_a_type_T_224_mask = do_enq;
  assign ram_a_type_T_224_en = do_enq;
  assign ram_union_T_254_addr = 1'h0;
  assign ram_union_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_union_T_254_data = ram_union[ram_union_T_254_addr];
  `else
  assign ram_union_T_254_data = ram_union_T_254_addr >= 1'h1 ? $random : ram_union[ram_union_T_254_addr];
  `endif
  assign ram_union_T_224_data = io_enq_bits_union;
  assign ram_union_T_224_addr = 1'h0;
  assign ram_union_T_224_mask = do_enq;
  assign ram_union_T_224_en = do_enq;
  assign ram_data_T_254_addr = 1'h0;
  assign ram_data_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_254_data = ram_data[ram_data_T_254_addr];
  `else
  assign ram_data_T_254_data = ram_data_T_254_addr >= 1'h1 ? $random : ram_data[ram_data_T_254_addr];
  `endif
  assign ram_data_T_224_data = io_enq_bits_data;
  assign ram_data_T_224_addr = 1'h0;
  assign ram_data_T_224_mask = do_enq;
  assign ram_data_T_224_en = do_enq;
  assign T_221 = maybe_full == 1'h0;
  assign T_222 = io_enq_ready & io_enq_valid;
  assign do_enq = T_222;
  assign T_223 = io_deq_ready & io_deq_valid;
  assign do_deq = T_223;
  assign T_249 = do_enq != do_deq;
  assign GEN_17 = T_249 ? do_enq : maybe_full;
  assign T_251 = T_221 == 1'h0;
  assign T_277 = 1'h0 - 1'h0;
  assign ptr_diff = T_277[0:0];
  assign T_279 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_block[initvar] = GEN_0[25:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_client_xact_id[initvar] = GEN_1[1:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr_beat[initvar] = GEN_2[2:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_is_builtin_type[initvar] = GEN_3[0:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_a_type[initvar] = GEN_4[2:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_union[initvar] = GEN_5[11:0];
  GEN_6 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_6[63:0];
  GEN_7 = {1{$random}};
  maybe_full = GEN_7[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_block_T_224_en & ram_addr_block_T_224_mask) begin
      ram_addr_block[ram_addr_block_T_224_addr] <= ram_addr_block_T_224_data;
    end
    if(ram_client_xact_id_T_224_en & ram_client_xact_id_T_224_mask) begin
      ram_client_xact_id[ram_client_xact_id_T_224_addr] <= ram_client_xact_id_T_224_data;
    end
    if(ram_addr_beat_T_224_en & ram_addr_beat_T_224_mask) begin
      ram_addr_beat[ram_addr_beat_T_224_addr] <= ram_addr_beat_T_224_data;
    end
    if(ram_is_builtin_type_T_224_en & ram_is_builtin_type_T_224_mask) begin
      ram_is_builtin_type[ram_is_builtin_type_T_224_addr] <= ram_is_builtin_type_T_224_data;
    end
    if(ram_a_type_T_224_en & ram_a_type_T_224_mask) begin
      ram_a_type[ram_a_type_T_224_addr] <= ram_a_type_T_224_data;
    end
    if(ram_union_T_224_en & ram_union_T_224_mask) begin
      ram_union[ram_union_T_224_addr] <= ram_union_T_224_data;
    end
    if(ram_data_T_224_en & ram_data_T_224_mask) begin
      ram_data[ram_data_T_224_addr] <= ram_data_T_224_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_17;
    end
  end
endmodule
module RTC(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_irqs_0
);
  reg [63:0] regs_0;
  reg [63:0] GEN_6;
  reg [63:0] regs_1;
  reg [63:0] GEN_9;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire [2:0] T_461;
  wire [28:0] T_462;
  wire [31:0] full_addr;
  wire  addr;
  wire  T_464;
  wire  read;
  wire  T_466;
  wire  write;
  wire  T_468;
  wire  T_469;
  wire [7:0] GEN_14;
  wire [8:0] T_473;
  wire [7:0] T_474;
  wire [7:0] T_480_0;
  wire  T_483;
  wire  T_484;
  wire  T_488;
  wire [7:0] T_489;
  wire [7:0] T_491;
  wire [7:0] T_492;
  wire  T_493;
  wire  T_494;
  wire  T_495;
  wire  T_496;
  wire  T_497;
  wire  T_498;
  wire  T_499;
  wire  T_500;
  wire [7:0] GEN_15;
  wire [8:0] T_502;
  wire [7:0] T_503;
  wire [7:0] GEN_16;
  wire [8:0] T_505;
  wire [7:0] T_506;
  wire [7:0] GEN_17;
  wire [8:0] T_508;
  wire [7:0] T_509;
  wire [7:0] GEN_18;
  wire [8:0] T_511;
  wire [7:0] T_512;
  wire [7:0] GEN_19;
  wire [8:0] T_514;
  wire [7:0] T_515;
  wire [7:0] GEN_20;
  wire [8:0] T_517;
  wire [7:0] T_518;
  wire [7:0] GEN_21;
  wire [8:0] T_520;
  wire [7:0] T_521;
  wire [7:0] GEN_22;
  wire [8:0] T_523;
  wire [7:0] T_524;
  wire [7:0] T_530_0;
  wire [7:0] T_530_1;
  wire [7:0] T_530_2;
  wire [7:0] T_530_3;
  wire [7:0] T_530_4;
  wire [7:0] T_530_5;
  wire [7:0] T_530_6;
  wire [7:0] T_530_7;
  wire [15:0] T_532;
  wire [15:0] T_533;
  wire [31:0] T_534;
  wire [15:0] T_535;
  wire [15:0] T_536;
  wire [31:0] T_537;
  wire [63:0] wmask;
  wire  T_539;
  wire  T_540;
  wire  T_541;
  wire  T_542;
  wire  T_544;
  wire  T_561;
  wire [2:0] T_562;
  wire  T_563;
  wire [2:0] T_564;
  wire  T_565;
  wire [2:0] T_566;
  wire  T_567;
  wire [2:0] T_568;
  wire  T_569;
  wire [2:0] T_570;
  wire  T_571;
  wire [2:0] T_572;
  wire  T_573;
  wire [2:0] T_574;
  wire [2:0] T_599_addr_beat;
  wire [1:0] T_599_client_xact_id;
  wire  T_599_manager_xact_id;
  wire  T_599_is_builtin_type;
  wire [3:0] T_599_g_type;
  wire [63:0] T_599_data;
  wire [63:0] GEN_0;
  wire [63:0] GEN_3;
  wire  T_621;
  reg [6:0] T_623;
  reg [31:0] GEN_10;
  wire  T_625;
  wire [6:0] GEN_23;
  wire [7:0] T_627;
  wire [6:0] T_628;
  wire [6:0] GEN_4;
  wire [63:0] GEN_24;
  wire [64:0] T_631;
  wire [63:0] T_632;
  wire [63:0] GEN_5;
  wire  T_633;
  wire [63:0] T_634;
  wire [63:0] T_635;
  wire [63:0] GEN_1;
  wire [63:0] T_636;
  wire [63:0] T_637;
  wire [63:0] GEN_2;
  wire [63:0] GEN_7;
  wire [63:0] GEN_8;
  wire [63:0] GEN_11;
  wire [63:0] GEN_12;
  wire [63:0] GEN_13;
  Queue_49 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_599_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_599_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_599_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_599_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_599_g_type;
  assign io_tl_grant_bits_data = T_599_data;
  assign io_irqs_0 = T_621;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_461 = acq_io_deq_bits_union[11:9];
  assign T_462 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign full_addr = {T_462,T_461};
  assign addr = full_addr[3];
  assign T_464 = acq_io_deq_bits_a_type == 3'h0;
  assign read = acq_io_deq_bits_is_builtin_type & T_464;
  assign T_466 = acq_io_deq_bits_a_type == 3'h2;
  assign write = acq_io_deq_bits_is_builtin_type & T_466;
  assign T_468 = acq_io_deq_bits_a_type == 3'h4;
  assign T_469 = acq_io_deq_bits_is_builtin_type & T_468;
  assign GEN_14 = {{7'd0}, 1'h1};
  assign T_473 = 8'h0 - GEN_14;
  assign T_474 = T_473[7:0];
  assign T_480_0 = T_474;
  assign T_483 = acq_io_deq_bits_a_type == 3'h3;
  assign T_484 = acq_io_deq_bits_is_builtin_type & T_483;
  assign T_488 = T_484 | write;
  assign T_489 = acq_io_deq_bits_union[8:1];
  assign T_491 = T_488 ? T_489 : {{7'd0}, 1'h0};
  assign T_492 = T_469 ? T_480_0 : T_491;
  assign T_493 = T_492[0];
  assign T_494 = T_492[1];
  assign T_495 = T_492[2];
  assign T_496 = T_492[3];
  assign T_497 = T_492[4];
  assign T_498 = T_492[5];
  assign T_499 = T_492[6];
  assign T_500 = T_492[7];
  assign GEN_15 = {{7'd0}, T_493};
  assign T_502 = 8'h0 - GEN_15;
  assign T_503 = T_502[7:0];
  assign GEN_16 = {{7'd0}, T_494};
  assign T_505 = 8'h0 - GEN_16;
  assign T_506 = T_505[7:0];
  assign GEN_17 = {{7'd0}, T_495};
  assign T_508 = 8'h0 - GEN_17;
  assign T_509 = T_508[7:0];
  assign GEN_18 = {{7'd0}, T_496};
  assign T_511 = 8'h0 - GEN_18;
  assign T_512 = T_511[7:0];
  assign GEN_19 = {{7'd0}, T_497};
  assign T_514 = 8'h0 - GEN_19;
  assign T_515 = T_514[7:0];
  assign GEN_20 = {{7'd0}, T_498};
  assign T_517 = 8'h0 - GEN_20;
  assign T_518 = T_517[7:0];
  assign GEN_21 = {{7'd0}, T_499};
  assign T_520 = 8'h0 - GEN_21;
  assign T_521 = T_520[7:0];
  assign GEN_22 = {{7'd0}, T_500};
  assign T_523 = 8'h0 - GEN_22;
  assign T_524 = T_523[7:0];
  assign T_530_0 = T_503;
  assign T_530_1 = T_506;
  assign T_530_2 = T_509;
  assign T_530_3 = T_512;
  assign T_530_4 = T_515;
  assign T_530_5 = T_518;
  assign T_530_6 = T_521;
  assign T_530_7 = T_524;
  assign T_532 = {T_530_1,T_530_0};
  assign T_533 = {T_530_3,T_530_2};
  assign T_534 = {T_533,T_532};
  assign T_535 = {T_530_5,T_530_4};
  assign T_536 = {T_530_7,T_530_6};
  assign T_537 = {T_536,T_535};
  assign wmask = {T_537,T_534};
  assign T_539 = acq_io_deq_valid == 1'h0;
  assign T_540 = T_539 | read;
  assign T_541 = T_540 | write;
  assign T_542 = T_541 | reset;
  assign T_544 = T_542 == 1'h0;
  assign T_561 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_562 = T_561 ? 3'h1 : 3'h3;
  assign T_563 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_564 = T_563 ? 3'h1 : T_562;
  assign T_565 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_566 = T_565 ? 3'h4 : T_564;
  assign T_567 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_568 = T_567 ? 3'h3 : T_566;
  assign T_569 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_570 = T_569 ? 3'h3 : T_568;
  assign T_571 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_572 = T_571 ? 3'h5 : T_570;
  assign T_573 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_574 = T_573 ? 3'h4 : T_572;
  assign T_599_addr_beat = {{2'd0}, 1'h0};
  assign T_599_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_599_manager_xact_id = 1'h0;
  assign T_599_is_builtin_type = 1'h1;
  assign T_599_g_type = {{1'd0}, T_574};
  assign T_599_data = GEN_0;
  assign GEN_0 = GEN_3;
  assign GEN_3 = addr ? regs_1 : regs_0;
  assign T_621 = regs_0 >= regs_1;
  assign T_625 = T_623 == 7'h63;
  assign GEN_23 = {{6'd0}, 1'h1};
  assign T_627 = T_623 + GEN_23;
  assign T_628 = T_627[6:0];
  assign GEN_4 = T_625 ? {{6'd0}, 1'h0} : T_628;
  assign GEN_24 = {{63'd0}, 1'h1};
  assign T_631 = regs_0 + GEN_24;
  assign T_632 = T_631[63:0];
  assign GEN_5 = T_625 ? T_632 : regs_0;
  assign T_633 = acq_io_deq_valid & write;
  assign T_634 = acq_io_deq_bits_data & wmask;
  assign T_635 = ~ wmask;
  assign GEN_1 = GEN_3;
  assign T_636 = GEN_1 & T_635;
  assign T_637 = T_634 | T_636;
  assign GEN_2 = T_637;
  assign GEN_7 = 1'h0 == addr ? GEN_2 : GEN_5;
  assign GEN_8 = addr ? GEN_2 : regs_1;
  assign GEN_11 = T_633 ? GEN_7 : GEN_5;
  assign GEN_12 = T_633 ? GEN_8 : regs_1;
  assign GEN_13 = reset ? {{63'd0}, 1'h0} : GEN_11;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_6 = {2{$random}};
  regs_0 = GEN_6[63:0];
  GEN_9 = {2{$random}};
  regs_1 = GEN_9[63:0];
  GEN_10 = {1{$random}};
  T_623 = GEN_10[6:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      regs_0 <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      regs_1 <= GEN_12;
    end
    if(reset) begin
      T_623 <= 7'h0;
    end else begin
      T_623 <= GEN_4;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_544) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported RTC operation\n    at rtc.scala:32 assert(!acq.valid || read || write, \"unsupported RTC operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_544) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  output  io_harts_0,
  output  io_harts_1,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_477_0;
  wire  T_477_1;
  wire  T_477_2;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  T_489_0;
  wire  T_489_1;
  wire  threshold_0;
  wire  threshold_1;
  wire  T_502_0;
  wire  T_502_1;
  wire  T_502_2;
  reg  pending_0;
  reg [31:0] GEN_15;
  reg  pending_1;
  reg [31:0] GEN_18;
  reg  pending_2;
  reg [31:0] GEN_19;
  reg  enables_0_0;
  reg [31:0] GEN_29;
  reg  enables_0_1;
  reg [31:0] GEN_32;
  reg  enables_0_2;
  reg [31:0] GEN_33;
  reg  enables_1_0;
  reg [31:0] GEN_36;
  reg  enables_1_1;
  reg [31:0] GEN_37;
  reg  enables_1_2;
  reg [31:0] GEN_38;
  wire  T_545;
  wire  GEN_11;
  wire  T_549;
  wire  GEN_12;
  wire [1:0] maxDevs_0;
  wire [1:0] maxDevs_1;
  wire  T_559;
  wire [1:0] T_560;
  wire  T_561;
  wire [1:0] T_562;
  wire  T_567;
  wire [1:0] T_568;
  wire [1:0] T_570;
  wire  T_571;
  wire  T_572;
  wire  T_574;
  wire [1:0] T_575;
  wire [1:0] GEN_101;
  wire [2:0] T_577;
  wire [1:0] T_578;
  wire [1:0] T_579;
  reg [1:0] T_580;
  reg [31:0] GEN_41;
  reg [1:0] T_581;
  reg [31:0] GEN_43;
  wire [1:0] T_583;
  wire  T_584;
  wire  T_585;
  wire [1:0] T_586;
  wire  T_587;
  wire [1:0] T_588;
  wire  T_593;
  wire [1:0] T_594;
  wire  T_598;
  wire  T_600;
  wire [1:0] T_601;
  wire [1:0] T_605;
  reg [1:0] T_606;
  reg [31:0] GEN_44;
  reg [1:0] T_607;
  reg [31:0] GEN_47;
  wire [1:0] T_609;
  wire  T_610;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_634;
  wire  T_636;
  wire  T_637;
  wire  read;
  wire  T_640;
  wire  T_641;
  wire  write;
  wire  T_644;
  wire  T_645;
  wire  T_646;
  wire  T_647;
  wire  T_649;
  wire [2:0] T_650;
  wire [28:0] T_651;
  wire [31:0] T_652;
  wire [25:0] addr;
  wire [25:0] GEN_103;
  wire [26:0] T_654;
  wire [25:0] T_655;
  wire  claimant;
  wire  hart;
  wire [1:0] GEN_0;
  wire [1:0] GEN_13;
  wire [2:0] T_657;
  wire [1:0] myMaxDev;
  wire [63:0] rdata;
  wire  T_663;
  wire  T_664;
  wire [7:0] GEN_105;
  wire [8:0] T_668;
  wire [7:0] T_669;
  wire [7:0] T_675_0;
  wire  T_678;
  wire  T_679;
  wire  T_683;
  wire [7:0] T_684;
  wire [7:0] T_686;
  wire [7:0] T_687;
  wire  T_688;
  wire  T_689;
  wire  T_690;
  wire  T_691;
  wire  T_692;
  wire  T_693;
  wire  T_694;
  wire  T_695;
  wire [7:0] GEN_106;
  wire [8:0] T_697;
  wire [7:0] T_698;
  wire [7:0] GEN_107;
  wire [8:0] T_700;
  wire [7:0] T_701;
  wire [7:0] GEN_108;
  wire [8:0] T_703;
  wire [7:0] T_704;
  wire [7:0] GEN_109;
  wire [8:0] T_706;
  wire [7:0] T_707;
  wire [7:0] GEN_110;
  wire [8:0] T_709;
  wire [7:0] T_710;
  wire [7:0] GEN_111;
  wire [8:0] T_712;
  wire [7:0] T_713;
  wire [7:0] GEN_112;
  wire [8:0] T_715;
  wire [7:0] T_716;
  wire [7:0] GEN_113;
  wire [8:0] T_718;
  wire [7:0] T_719;
  wire [7:0] T_725_0;
  wire [7:0] T_725_1;
  wire [7:0] T_725_2;
  wire [7:0] T_725_3;
  wire [7:0] T_725_4;
  wire [7:0] T_725_5;
  wire [7:0] T_725_6;
  wire [7:0] T_725_7;
  wire [15:0] T_727;
  wire [15:0] T_728;
  wire [31:0] T_729;
  wire [15:0] T_730;
  wire [15:0] T_731;
  wire [31:0] T_732;
  wire [63:0] T_733;
  wire [63:0] T_734;
  wire [7:0] T_748_0;
  wire [7:0] T_760;
  wire  T_761;
  wire  T_762;
  wire  T_763;
  wire  T_764;
  wire  T_765;
  wire  T_766;
  wire  T_767;
  wire  T_768;
  wire [7:0] GEN_115;
  wire [8:0] T_770;
  wire [7:0] T_771;
  wire [7:0] GEN_116;
  wire [8:0] T_773;
  wire [7:0] T_774;
  wire [7:0] GEN_117;
  wire [8:0] T_776;
  wire [7:0] T_777;
  wire [7:0] GEN_118;
  wire [8:0] T_779;
  wire [7:0] T_780;
  wire [7:0] GEN_119;
  wire [8:0] T_782;
  wire [7:0] T_783;
  wire [7:0] GEN_120;
  wire [8:0] T_785;
  wire [7:0] T_786;
  wire [7:0] GEN_121;
  wire [8:0] T_788;
  wire [7:0] T_789;
  wire [7:0] GEN_122;
  wire [8:0] T_791;
  wire [7:0] T_792;
  wire [7:0] T_798_0;
  wire [7:0] T_798_1;
  wire [7:0] T_798_2;
  wire [7:0] T_798_3;
  wire [7:0] T_798_4;
  wire [7:0] T_798_5;
  wire [7:0] T_798_6;
  wire [7:0] T_798_7;
  wire [15:0] T_800;
  wire [15:0] T_801;
  wire [31:0] T_802;
  wire [15:0] T_803;
  wire [15:0] T_804;
  wire [31:0] T_805;
  wire [63:0] T_806;
  wire [63:0] T_807;
  wire [63:0] T_808;
  wire [63:0] masked_wdata;
  wire  T_810;
  wire [32:0] T_813;
  wire  GEN_1;
  wire  GEN_14;
  wire [33:0] T_814;
  wire [6:0] GEN_124;
  wire [7:0] T_816;
  wire [33:0] T_817;
  wire  T_818;
  wire  T_819;
  wire  GEN_2;
  wire [1:0] GEN_126;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_20;
  wire  GEN_21;
  wire [7:0] T_834_0;
  wire [7:0] T_846;
  wire  T_847;
  wire [31:0] T_848;
  wire [1:0] T_849;
  wire  GEN_3;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_22;
  wire  GEN_132;
  wire  GEN_23;
  wire  GEN_134;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire [2:0] T_851;
  wire [1:0] T_852;
  wire  GEN_4;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_39;
  wire  GEN_40;
  wire [63:0] GEN_42;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_50;
  wire  GEN_51;
  wire [25:0] GEN_141;
  wire  T_860;
  wire  T_862;
  wire  T_863;
  wire [26:0] T_865;
  wire [25:0] T_866;
  wire  T_867;
  wire  GEN_5;
  wire  GEN_52;
  wire  GEN_6;
  wire  GEN_53;
  wire [1:0] T_871;
  wire  GEN_7;
  wire  GEN_54;
  wire [2:0] T_872;
  wire  T_876;
  wire  GEN_8;
  wire  T_880;
  wire  GEN_9;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_63;
  wire  GEN_64;
  wire  T_884;
  wire  GEN_10;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_68;
  wire  GEN_69;
  wire [63:0] GEN_73;
  wire  GEN_83;
  wire [63:0] GEN_87;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_95;
  wire  GEN_96;
  wire [25:0] GEN_143;
  wire  T_886;
  wire  T_890;
  wire  T_891;
  wire  T_892;
  wire [1:0] T_894;
  wire [2:0] T_895;
  wire [2:0] T_898;
  wire [63:0] GEN_97;
  wire  T_905;
  wire  T_906;
  wire  T_907;
  wire  T_909;
  wire [31:0] T_911;
  wire [31:0] T_913;
  wire [63:0] T_914;
  wire [63:0] GEN_98;
  wire [31:0] T_918;
  wire [63:0] GEN_99;
  wire [63:0] GEN_100;
  wire  T_939;
  wire [2:0] T_940;
  wire  T_941;
  wire [2:0] T_942;
  wire  T_943;
  wire [2:0] T_944;
  wire  T_945;
  wire [2:0] T_946;
  wire  T_947;
  wire [2:0] T_948;
  wire  T_949;
  wire [2:0] T_950;
  wire  T_951;
  wire [2:0] T_952;
  wire [2:0] T_977_addr_beat;
  wire [1:0] T_977_client_xact_id;
  wire  T_977_manager_xact_id;
  wire  T_977_is_builtin_type;
  wire [3:0] T_977_g_type;
  wire [63:0] T_977_data;
  Queue_49 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_545;
  assign io_devices_0_complete = GEN_50;
  assign io_devices_1_ready = T_549;
  assign io_devices_1_complete = GEN_51;
  assign io_harts_0 = T_584;
  assign io_harts_1 = T_610;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_977_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_977_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_977_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_977_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_977_g_type;
  assign io_tl_grant_bits_data = T_977_data;
  assign T_477_0 = 1'h1;
  assign T_477_1 = 1'h1;
  assign T_477_2 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_477_1;
  assign priority_2 = T_477_2;
  assign T_489_0 = 1'h0;
  assign T_489_1 = 1'h0;
  assign threshold_0 = T_489_0;
  assign threshold_1 = T_489_1;
  assign T_502_0 = 1'h0;
  assign T_502_1 = 1'h0;
  assign T_502_2 = 1'h0;
  assign T_545 = pending_1 == 1'h0;
  assign GEN_11 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_549 = pending_2 == 1'h0;
  assign GEN_12 = io_devices_1_valid ? 1'h1 : pending_2;
  assign maxDevs_0 = T_580;
  assign maxDevs_1 = T_606;
  assign T_559 = pending_1 & enables_0_1;
  assign T_560 = {T_559,priority_1};
  assign T_561 = pending_2 & enables_0_2;
  assign T_562 = {T_561,priority_2};
  assign T_567 = 2'h2 >= T_560;
  assign T_568 = T_567 ? 2'h2 : T_560;
  assign T_570 = 1'h1 + 1'h0;
  assign T_571 = T_570[0:0];
  assign T_572 = T_567 ? 1'h0 : T_571;
  assign T_574 = T_568 >= T_562;
  assign T_575 = T_574 ? T_568 : T_562;
  assign GEN_101 = {{1'd0}, 1'h0};
  assign T_577 = 2'h2 + GEN_101;
  assign T_578 = T_577[1:0];
  assign T_579 = T_574 ? {{1'd0}, T_572} : T_578;
  assign T_583 = {1'h1,threshold_0};
  assign T_584 = T_581 > T_583;
  assign T_585 = pending_1 & enables_1_1;
  assign T_586 = {T_585,priority_1};
  assign T_587 = pending_2 & enables_1_2;
  assign T_588 = {T_587,priority_2};
  assign T_593 = 2'h2 >= T_586;
  assign T_594 = T_593 ? 2'h2 : T_586;
  assign T_598 = T_593 ? 1'h0 : T_571;
  assign T_600 = T_594 >= T_588;
  assign T_601 = T_600 ? T_594 : T_588;
  assign T_605 = T_600 ? {{1'd0}, T_598} : T_578;
  assign T_609 = {1'h1,threshold_1};
  assign T_610 = T_607 > T_609;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_634 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_636 = acq_io_deq_bits_a_type == 3'h0;
  assign T_637 = acq_io_deq_bits_is_builtin_type & T_636;
  assign read = T_634 & T_637;
  assign T_640 = acq_io_deq_bits_a_type == 3'h2;
  assign T_641 = acq_io_deq_bits_is_builtin_type & T_640;
  assign write = T_634 & T_641;
  assign T_644 = T_634 == 1'h0;
  assign T_645 = T_644 | read;
  assign T_646 = T_645 | write;
  assign T_647 = T_646 | reset;
  assign T_649 = T_647 == 1'h0;
  assign T_650 = acq_io_deq_bits_union[11:9];
  assign T_651 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_652 = {T_651,T_650};
  assign addr = T_652[25:0];
  assign GEN_103 = {{4'd0}, 22'h200000};
  assign T_654 = addr - GEN_103;
  assign T_655 = T_654[25:0];
  assign claimant = T_655[12];
  assign hart = GEN_83;
  assign GEN_0 = GEN_13;
  assign GEN_13 = claimant ? maxDevs_1 : maxDevs_0;
  assign T_657 = GEN_0 + GEN_101;
  assign myMaxDev = T_657[1:0];
  assign rdata = GEN_100;
  assign T_663 = acq_io_deq_bits_a_type == 3'h4;
  assign T_664 = acq_io_deq_bits_is_builtin_type & T_663;
  assign GEN_105 = {{7'd0}, 1'h1};
  assign T_668 = 8'h0 - GEN_105;
  assign T_669 = T_668[7:0];
  assign T_675_0 = T_669;
  assign T_678 = acq_io_deq_bits_a_type == 3'h3;
  assign T_679 = acq_io_deq_bits_is_builtin_type & T_678;
  assign T_683 = T_679 | T_641;
  assign T_684 = acq_io_deq_bits_union[8:1];
  assign T_686 = T_683 ? T_684 : {{7'd0}, 1'h0};
  assign T_687 = T_664 ? T_675_0 : T_686;
  assign T_688 = T_687[0];
  assign T_689 = T_687[1];
  assign T_690 = T_687[2];
  assign T_691 = T_687[3];
  assign T_692 = T_687[4];
  assign T_693 = T_687[5];
  assign T_694 = T_687[6];
  assign T_695 = T_687[7];
  assign GEN_106 = {{7'd0}, T_688};
  assign T_697 = 8'h0 - GEN_106;
  assign T_698 = T_697[7:0];
  assign GEN_107 = {{7'd0}, T_689};
  assign T_700 = 8'h0 - GEN_107;
  assign T_701 = T_700[7:0];
  assign GEN_108 = {{7'd0}, T_690};
  assign T_703 = 8'h0 - GEN_108;
  assign T_704 = T_703[7:0];
  assign GEN_109 = {{7'd0}, T_691};
  assign T_706 = 8'h0 - GEN_109;
  assign T_707 = T_706[7:0];
  assign GEN_110 = {{7'd0}, T_692};
  assign T_709 = 8'h0 - GEN_110;
  assign T_710 = T_709[7:0];
  assign GEN_111 = {{7'd0}, T_693};
  assign T_712 = 8'h0 - GEN_111;
  assign T_713 = T_712[7:0];
  assign GEN_112 = {{7'd0}, T_694};
  assign T_715 = 8'h0 - GEN_112;
  assign T_716 = T_715[7:0];
  assign GEN_113 = {{7'd0}, T_695};
  assign T_718 = 8'h0 - GEN_113;
  assign T_719 = T_718[7:0];
  assign T_725_0 = T_698;
  assign T_725_1 = T_701;
  assign T_725_2 = T_704;
  assign T_725_3 = T_707;
  assign T_725_4 = T_710;
  assign T_725_5 = T_713;
  assign T_725_6 = T_716;
  assign T_725_7 = T_719;
  assign T_727 = {T_725_1,T_725_0};
  assign T_728 = {T_725_3,T_725_2};
  assign T_729 = {T_728,T_727};
  assign T_730 = {T_725_5,T_725_4};
  assign T_731 = {T_725_7,T_725_6};
  assign T_732 = {T_731,T_730};
  assign T_733 = {T_732,T_729};
  assign T_734 = acq_io_deq_bits_data & T_733;
  assign T_748_0 = T_669;
  assign T_760 = T_664 ? T_748_0 : T_686;
  assign T_761 = T_760[0];
  assign T_762 = T_760[1];
  assign T_763 = T_760[2];
  assign T_764 = T_760[3];
  assign T_765 = T_760[4];
  assign T_766 = T_760[5];
  assign T_767 = T_760[6];
  assign T_768 = T_760[7];
  assign GEN_115 = {{7'd0}, T_761};
  assign T_770 = 8'h0 - GEN_115;
  assign T_771 = T_770[7:0];
  assign GEN_116 = {{7'd0}, T_762};
  assign T_773 = 8'h0 - GEN_116;
  assign T_774 = T_773[7:0];
  assign GEN_117 = {{7'd0}, T_763};
  assign T_776 = 8'h0 - GEN_117;
  assign T_777 = T_776[7:0];
  assign GEN_118 = {{7'd0}, T_764};
  assign T_779 = 8'h0 - GEN_118;
  assign T_780 = T_779[7:0];
  assign GEN_119 = {{7'd0}, T_765};
  assign T_782 = 8'h0 - GEN_119;
  assign T_783 = T_782[7:0];
  assign GEN_120 = {{7'd0}, T_766};
  assign T_785 = 8'h0 - GEN_120;
  assign T_786 = T_785[7:0];
  assign GEN_121 = {{7'd0}, T_767};
  assign T_788 = 8'h0 - GEN_121;
  assign T_789 = T_788[7:0];
  assign GEN_122 = {{7'd0}, T_768};
  assign T_791 = 8'h0 - GEN_122;
  assign T_792 = T_791[7:0];
  assign T_798_0 = T_771;
  assign T_798_1 = T_774;
  assign T_798_2 = T_777;
  assign T_798_3 = T_780;
  assign T_798_4 = T_783;
  assign T_798_5 = T_786;
  assign T_798_6 = T_789;
  assign T_798_7 = T_792;
  assign T_800 = {T_798_1,T_798_0};
  assign T_801 = {T_798_3,T_798_2};
  assign T_802 = {T_801,T_800};
  assign T_803 = {T_798_5,T_798_4};
  assign T_804 = {T_798_7,T_798_6};
  assign T_805 = {T_804,T_803};
  assign T_806 = {T_805,T_802};
  assign T_807 = ~ T_806;
  assign T_808 = rdata & T_807;
  assign masked_wdata = T_734 | T_808;
  assign T_810 = addr >= GEN_103;
  assign T_813 = {myMaxDev,31'h0};
  assign GEN_1 = GEN_14;
  assign GEN_14 = claimant ? threshold_1 : threshold_0;
  assign T_814 = {T_813,GEN_1};
  assign GEN_124 = {{6'd0}, 1'h0};
  assign T_816 = GEN_124 * 7'h40;
  assign T_817 = T_814 >> T_816;
  assign T_818 = addr[2];
  assign T_819 = read & T_818;
  assign GEN_2 = 1'h0;
  assign GEN_126 = {{1'd0}, 1'h1};
  assign GEN_16 = GEN_126 == myMaxDev ? GEN_2 : GEN_11;
  assign GEN_17 = 2'h2 == myMaxDev ? GEN_2 : GEN_12;
  assign GEN_20 = T_819 ? GEN_16 : GEN_11;
  assign GEN_21 = T_819 ? GEN_17 : GEN_12;
  assign T_834_0 = T_669;
  assign T_846 = T_664 ? T_834_0 : T_686;
  assign T_847 = T_846[4];
  assign T_848 = acq_io_deq_bits_data[63:32];
  assign T_849 = T_848[1:0];
  assign GEN_3 = GEN_26;
  assign GEN_129 = 1'h0 == hart;
  assign GEN_130 = GEN_126 == T_849;
  assign GEN_22 = GEN_129 & GEN_130 ? enables_0_1 : enables_0_0;
  assign GEN_132 = 2'h2 == T_849;
  assign GEN_23 = GEN_129 & GEN_132 ? enables_0_2 : GEN_22;
  assign GEN_134 = GEN_101 == T_849;
  assign GEN_24 = hart & GEN_134 ? enables_1_0 : GEN_23;
  assign GEN_25 = hart & GEN_130 ? enables_1_1 : GEN_24;
  assign GEN_26 = hart & GEN_132 ? enables_1_2 : GEN_25;
  assign T_851 = T_849 - GEN_126;
  assign T_852 = T_851[1:0];
  assign GEN_4 = 1'h1;
  assign GEN_27 = GEN_101 == T_852 ? GEN_4 : 1'h0;
  assign GEN_28 = GEN_126 == T_852 ? GEN_4 : 1'h0;
  assign GEN_30 = GEN_3 ? GEN_27 : 1'h0;
  assign GEN_31 = GEN_3 ? GEN_28 : 1'h0;
  assign GEN_34 = T_847 ? GEN_30 : 1'h0;
  assign GEN_35 = T_847 ? GEN_31 : 1'h0;
  assign GEN_39 = write ? GEN_34 : 1'h0;
  assign GEN_40 = write ? GEN_35 : 1'h0;
  assign GEN_42 = T_810 ? {{30'd0}, T_817} : 64'h0;
  assign GEN_45 = T_810 ? GEN_20 : GEN_11;
  assign GEN_46 = T_810 ? GEN_21 : GEN_12;
  assign GEN_50 = T_810 ? GEN_39 : 1'h0;
  assign GEN_51 = T_810 ? GEN_40 : 1'h0;
  assign GEN_141 = {{12'd0}, 14'h2000};
  assign T_860 = addr >= GEN_141;
  assign T_862 = T_810 == 1'h0;
  assign T_863 = T_862 & T_860;
  assign T_865 = addr - GEN_141;
  assign T_866 = T_865[25:0];
  assign T_867 = T_866[7];
  assign GEN_5 = GEN_52;
  assign GEN_52 = hart ? enables_1_2 : enables_0_2;
  assign GEN_6 = GEN_53;
  assign GEN_53 = hart ? enables_1_1 : enables_0_1;
  assign T_871 = {GEN_5,GEN_6};
  assign GEN_7 = GEN_54;
  assign GEN_54 = hart ? enables_1_0 : enables_0_0;
  assign T_872 = {T_871,GEN_7};
  assign T_876 = masked_wdata[0];
  assign GEN_8 = T_876;
  assign T_880 = masked_wdata[1];
  assign GEN_9 = T_880;
  assign GEN_60 = 1'h0 == T_867 ? GEN_9 : enables_0_1;
  assign GEN_61 = T_867 ? GEN_9 : enables_1_1;
  assign GEN_63 = write ? GEN_60 : enables_0_1;
  assign GEN_64 = write ? GEN_61 : enables_1_1;
  assign T_884 = masked_wdata[2];
  assign GEN_10 = T_884;
  assign GEN_65 = 1'h0 == T_867 ? GEN_10 : enables_0_2;
  assign GEN_66 = T_867 ? GEN_10 : enables_1_2;
  assign GEN_68 = write ? GEN_65 : enables_0_2;
  assign GEN_69 = write ? GEN_66 : enables_1_2;
  assign GEN_73 = 1'h1 ? {{61'd0}, T_872} : GEN_42;
  assign GEN_83 = T_863 ? T_867 : claimant;
  assign GEN_87 = T_863 ? GEN_73 : GEN_42;
  assign GEN_92 = T_863 ? GEN_63 : enables_0_1;
  assign GEN_93 = T_863 ? GEN_64 : enables_1_1;
  assign GEN_95 = T_863 ? GEN_68 : enables_0_2;
  assign GEN_96 = T_863 ? GEN_69 : enables_1_2;
  assign GEN_143 = {{13'd0}, 13'h1000};
  assign T_886 = addr >= GEN_143;
  assign T_890 = T_860 == 1'h0;
  assign T_891 = T_862 & T_890;
  assign T_892 = T_891 & T_886;
  assign T_894 = {pending_2,pending_1};
  assign T_895 = {T_894,pending_0};
  assign T_898 = T_895 >> T_816;
  assign GEN_97 = T_892 ? {{61'd0}, T_898} : GEN_87;
  assign T_905 = T_886 == 1'h0;
  assign T_906 = T_891 & T_905;
  assign T_907 = addr[3];
  assign T_909 = T_907 == 1'h0;
  assign T_911 = {31'h0,priority_0};
  assign T_913 = {31'h0,priority_1};
  assign T_914 = {T_913,T_911};
  assign GEN_98 = T_909 ? T_914 : GEN_97;
  assign T_918 = {31'h0,priority_2};
  assign GEN_99 = T_907 ? {{32'd0}, T_918} : GEN_98;
  assign GEN_100 = T_906 ? GEN_99 : GEN_97;
  assign T_939 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_940 = T_939 ? 3'h1 : 3'h3;
  assign T_941 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_942 = T_941 ? 3'h1 : T_940;
  assign T_943 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_944 = T_943 ? 3'h4 : T_942;
  assign T_945 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_946 = T_945 ? 3'h3 : T_944;
  assign T_947 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_948 = T_947 ? 3'h3 : T_946;
  assign T_949 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_950 = T_949 ? 3'h5 : T_948;
  assign T_951 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_952 = T_951 ? 3'h4 : T_950;
  assign T_977_addr_beat = {{2'd0}, 1'h0};
  assign T_977_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_977_manager_xact_id = 1'h0;
  assign T_977_is_builtin_type = 1'h1;
  assign T_977_g_type = {{1'd0}, T_952};
  assign T_977_data = rdata;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  pending_0 = GEN_15[0:0];
  GEN_18 = {1{$random}};
  pending_1 = GEN_18[0:0];
  GEN_19 = {1{$random}};
  pending_2 = GEN_19[0:0];
  GEN_29 = {1{$random}};
  enables_0_0 = GEN_29[0:0];
  GEN_32 = {1{$random}};
  enables_0_1 = GEN_32[0:0];
  GEN_33 = {1{$random}};
  enables_0_2 = GEN_33[0:0];
  GEN_36 = {1{$random}};
  enables_1_0 = GEN_36[0:0];
  GEN_37 = {1{$random}};
  enables_1_1 = GEN_37[0:0];
  GEN_38 = {1{$random}};
  enables_1_2 = GEN_38[0:0];
  GEN_41 = {1{$random}};
  T_580 = GEN_41[1:0];
  GEN_43 = {1{$random}};
  T_581 = GEN_43[1:0];
  GEN_44 = {1{$random}};
  T_606 = GEN_44[1:0];
  GEN_47 = {1{$random}};
  T_607 = GEN_47[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_502_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_502_1;
    end else begin
      pending_1 <= GEN_45;
    end
    if(reset) begin
      pending_2 <= T_502_2;
    end else begin
      pending_2 <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      enables_0_1 <= GEN_92;
    end
    if(1'h0) begin
    end else begin
      enables_0_2 <= GEN_95;
    end
    if(1'h0) begin
    end else begin
      enables_1_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      enables_1_1 <= GEN_93;
    end
    if(1'h0) begin
    end else begin
      enables_1_2 <= GEN_96;
    end
    if(1'h0) begin
    end else begin
      T_580 <= T_579;
    end
    if(1'h0) begin
    end else begin
      T_581 <= T_575;
    end
    if(1'h0) begin
    end else begin
      T_606 <= T_605;
    end
    if(1'h0) begin
    end else begin
      T_607 <= T_601;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_649) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at plic.scala:107 assert(!acq.fire() || read || write, \"unsupported PLIC operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_649) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module LevelGateway(
  input   clk,
  input   reset,
  input   io_interrupt,
  output  io_plic_valid,
  input   io_plic_ready,
  input   io_plic_complete
);
  reg  inFlight;
  reg [31:0] GEN_2;
  wire  T_6;
  wire  GEN_0;
  wire  GEN_1;
  wire  T_10;
  wire  T_11;
  assign io_plic_valid = T_11;
  assign T_6 = io_interrupt & io_plic_ready;
  assign GEN_0 = T_6 ? 1'h1 : inFlight;
  assign GEN_1 = io_plic_complete ? 1'h0 : GEN_0;
  assign T_10 = inFlight == 1'h0;
  assign T_11 = io_interrupt & T_10;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_2 = {1{$random}};
  inFlight = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      inFlight <= 1'h0;
    end else begin
      inFlight <= GEN_1;
    end
  end
endmodule
module DebugModule(
  input   clk,
  input   reset,
  output  io_db_req_ready,
  input   io_db_req_valid,
  input  [4:0] io_db_req_bits_addr,
  input  [1:0] io_db_req_bits_op,
  input  [33:0] io_db_req_bits_data,
  input   io_db_resp_ready,
  output  io_db_resp_valid,
  output [1:0] io_db_resp_bits_resp,
  output [33:0] io_db_resp_bits_data,
  output  io_debugInterrupts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_ndreset,
  output  io_fullreset
);
  wire  CONTROLReset_interrupt;
  wire  CONTROLReset_haltnot;
  wire [9:0] CONTROLReset_reserved0;
  wire [2:0] CONTROLReset_buserror;
  wire [2:0] CONTROLReset_serial;
  wire  CONTROLReset_autoincrement;
  wire [2:0] CONTROLReset_access;
  wire [9:0] CONTROLReset_hartid;
  wire  CONTROLReset_ndreset;
  wire  CONTROLReset_fullreset;
  wire  CONTROLWrEn;
  reg  CONTROLReg_interrupt;
  reg [31:0] GEN_26;
  reg  CONTROLReg_haltnot;
  reg [31:0] GEN_27;
  reg [9:0] CONTROLReg_reserved0;
  reg [31:0] GEN_28;
  reg [2:0] CONTROLReg_buserror;
  reg [31:0] GEN_29;
  reg [2:0] CONTROLReg_serial;
  reg [31:0] GEN_30;
  reg  CONTROLReg_autoincrement;
  reg [31:0] GEN_52;
  reg [2:0] CONTROLReg_access;
  reg [31:0] GEN_94;
  reg [9:0] CONTROLReg_hartid;
  reg [31:0] GEN_95;
  reg  CONTROLReg_ndreset;
  reg [31:0] GEN_97;
  reg  CONTROLReg_fullreset;
  reg [31:0] GEN_98;
  wire  CONTROLWrData_interrupt;
  wire  CONTROLWrData_haltnot;
  wire [9:0] CONTROLWrData_reserved0;
  wire [2:0] CONTROLWrData_buserror;
  wire [2:0] CONTROLWrData_serial;
  wire  CONTROLWrData_autoincrement;
  wire [2:0] CONTROLWrData_access;
  wire [9:0] CONTROLWrData_hartid;
  wire  CONTROLWrData_ndreset;
  wire  CONTROLWrData_fullreset;
  wire  CONTROLRdData_interrupt;
  wire  CONTROLRdData_haltnot;
  wire [9:0] CONTROLRdData_reserved0;
  wire [2:0] CONTROLRdData_buserror;
  wire [2:0] CONTROLRdData_serial;
  wire  CONTROLRdData_autoincrement;
  wire [2:0] CONTROLRdData_access;
  wire [9:0] CONTROLRdData_hartid;
  wire  CONTROLRdData_ndreset;
  wire  CONTROLRdData_fullreset;
  reg  ndresetCtrReg;
  reg [31:0] GEN_99;
  wire [1:0] DMINFORdData_reserved0;
  wire [6:0] DMINFORdData_abussize;
  wire [3:0] DMINFORdData_serialcount;
  wire  DMINFORdData_access128;
  wire  DMINFORdData_access64;
  wire  DMINFORdData_access32;
  wire  DMINFORdData_access16;
  wire  DMINFORdData_accesss8;
  wire [5:0] DMINFORdData_dramsize;
  wire  DMINFORdData_haltsum;
  wire [2:0] DMINFORdData_reserved1;
  wire  DMINFORdData_authenticated;
  wire  DMINFORdData_authbusy;
  wire [1:0] DMINFORdData_authtype;
  wire [1:0] DMINFORdData_version;
  wire  HALTSUMRdData_serialfull;
  wire  HALTSUMRdData_serialvalid;
  wire [31:0] HALTSUMRdData_acks;
  wire  RAMWrData_interrupt;
  wire  RAMWrData_haltnot;
  wire [31:0] RAMWrData_data;
  wire  RAMRdData_interrupt;
  wire  RAMRdData_haltnot;
  wire [31:0] RAMRdData_data;
  wire  SETHALTNOTWrEn;
  wire [9:0] SETHALTNOTWrData;
  wire  CLEARDEBINTWrEn;
  wire [9:0] CLEARDEBINTWrData;
  wire  T_655_0;
  reg  interruptRegs_0;
  reg [31:0] GEN_120;
  wire  T_666_0;
  reg  haltnotRegs_0;
  reg [31:0] GEN_121;
  wire [31:0] haltnotStatus_0;
  wire [31:0] rdHaltnotStatus;
  wire [31:0] GEN_118;
  wire  haltnotSummary;
  reg [63:0] ramMem [0:7];
  reg [63:0] GEN_122;
  wire [63:0] ramMem_T_853_data;
  wire [2:0] ramMem_T_853_addr;
  wire  ramMem_T_853_en;
  wire [63:0] ramMem_T_854_data;
  wire [2:0] ramMem_T_854_addr;
  wire  ramMem_T_854_mask;
  wire  ramMem_T_854_en;
  wire [2:0] ramAddr;
  wire [63:0] ramRdData;
  wire [63:0] ramWrData;
  wire [63:0] ramWrMask;
  wire  ramWrEn;
  wire [3:0] dbRamAddr;
  wire [31:0] dbRamRdData;
  wire [31:0] dbRamWrData;
  wire  dbRamWrEn;
  wire  dbRamRdEn;
  wire [2:0] sbRamAddr;
  wire [63:0] sbRamRdData;
  wire [63:0] sbRamWrData;
  wire  sbRamWrEn;
  wire  sbRamRdEn;
  wire [63:0] sbRomRdData;
  wire  dbRdEn;
  wire  dbWrEn;
  wire [33:0] dbRdData;
  reg  dbStateReg;
  reg [31:0] GEN_140;
  wire [1:0] dbResult_resp;
  wire [33:0] dbResult_data;
  wire [4:0] dbReq_addr;
  wire [1:0] dbReq_op;
  wire [33:0] dbReq_data;
  reg [1:0] dbRespReg_resp;
  reg [31:0] GEN_141;
  reg [33:0] dbRespReg_data;
  reg [63:0] GEN_142;
  wire  rdCondWrFailure;
  wire  dbWrNeeded;
  wire [11:0] sbAddr;
  wire [63:0] sbRdData;
  wire [63:0] sbWrData;
  wire [63:0] sbWrMask;
  wire  sbWrEn;
  wire  sbRdEn;
  wire  stallFromDb;
  wire  stallFromSb;
  wire [9:0] GEN_119;
  wire  T_720;
  wire  T_721;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_723;
  wire  T_724;
  wire  T_726;
  wire  T_727;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_731;
  wire  T_732;
  wire  T_733;
  wire  T_735;
  wire  GEN_15;
  wire  GEN_16;
  wire  T_738;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_741;
  wire  T_742;
  wire  T_745;
  wire  GEN_19;
  wire  GEN_20;
  wire  T_750;
  wire  T_751;
  wire  T_754;
  wire  GEN_21;
  wire  GEN_22;
  wire [3:0] T_782;
  wire [2:0] T_783;
  wire [31:0] T_801_0;
  wire [31:0] T_801_1;
  wire [31:0] dbRamWrMask_0;
  wire [31:0] dbRamWrMask_1;
  wire  T_806;
  wire [31:0] T_807;
  wire [31:0] T_808;
  wire [31:0] T_814_0;
  wire [31:0] T_814_1;
  wire [31:0] T_823_0;
  wire [31:0] T_823_1;
  wire [31:0] GEN_0;
  wire [31:0] GEN_23;
  wire [31:0] GEN_24;
  wire [31:0] GEN_1;
  wire [31:0] GEN_25;
  wire [63:0] T_831;
  wire [63:0] T_832;
  wire  T_833;
  wire  T_834;
  wire  T_835;
  wire  T_837;
  wire  T_838;
  wire  T_840;
  wire [63:0] dbRamWrDataVec;
  wire [63:0] T_841;
  wire [63:0] T_842;
  wire [63:0] T_843;
  wire [63:0] T_844;
  wire [63:0] T_845;
  wire [63:0] T_848;
  wire [63:0] T_849;
  wire  T_850;
  wire [2:0] T_851;
  wire [2:0] T_852;
  wire  T_855;
  wire  T_878_interrupt;
  wire  T_878_haltnot;
  wire [9:0] T_878_reserved0;
  wire [2:0] T_878_buserror;
  wire [2:0] T_878_serial;
  wire  T_878_autoincrement;
  wire [2:0] T_878_access;
  wire [9:0] T_878_hartid;
  wire  T_878_ndreset;
  wire  T_878_fullreset;
  wire  T_889;
  wire  T_890;
  wire [9:0] T_891;
  wire [2:0] T_892;
  wire  T_893;
  wire [2:0] T_894;
  wire [2:0] T_895;
  wire [9:0] T_896;
  wire  T_897;
  wire  T_898;
  wire  T_907_interrupt;
  wire  T_907_haltnot;
  wire [31:0] T_907_data;
  wire [31:0] T_911;
  wire  T_916;
  wire  T_918;
  wire  GEN_31;
  wire  T_920;
  wire  T_922;
  wire  T_923;
  wire  GEN_32;
  wire  T_927;
  wire  T_928;
  wire  GEN_33;
  wire  GEN_34;
  wire [9:0] GEN_35;
  wire [2:0] GEN_36;
  wire [2:0] GEN_37;
  wire  GEN_38;
  wire [2:0] GEN_39;
  wire [9:0] GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  T_931;
  wire  T_932;
  wire  T_933;
  wire  GEN_44;
  wire  T_936;
  wire  T_938;
  wire [1:0] T_941;
  wire  T_942;
  wire  T_943;
  wire  GEN_45;
  wire [9:0] GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  T_948;
  wire  GEN_49;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [4:0] GEN_123;
  wire  T_961;
  wire [31:0] GEN_50;
  wire [1:0] T_966;
  wire [33:0] T_967;
  wire [33:0] GEN_51;
  wire [1:0] T_973;
  wire [3:0] T_974;
  wire [13:0] T_975;
  wire [15:0] T_976;
  wire [5:0] T_977;
  wire [1:0] T_978;
  wire [11:0] T_979;
  wire [17:0] T_980;
  wire [33:0] T_981;
  wire [33:0] GEN_53;
  wire  T_983;
  wire  T_989;
  wire [2:0] T_990;
  wire [4:0] T_991;
  wire [3:0] T_992;
  wire [6:0] T_993;
  wire [10:0] T_994;
  wire [15:0] T_995;
  wire [1:0] T_996;
  wire [1:0] T_997;
  wire [3:0] T_998;
  wire [4:0] T_999;
  wire [8:0] T_1000;
  wire [13:0] T_1001;
  wire [17:0] T_1002;
  wire [33:0] T_1003;
  wire [33:0] GEN_54;
  wire  T_1005;
  wire  T_1012;
  wire  T_1013;
  wire  T_1014;
  wire [33:0] GEN_55;
  wire [2:0] T_1016;
  wire  T_1018;
  wire  T_1028;
  wire  T_1029;
  wire  T_1030;
  wire [33:0] GEN_56;
  wire  T_1043;
  wire  T_1044;
  wire [33:0] GEN_57;
  wire  T_1046;
  wire  T_1048;
  wire  T_1049;
  wire  T_1051;
  wire  T_1054;
  wire  T_1055;
  wire  T_1056;
  wire [1:0] T_1059;
  wire  T_1061;
  wire  T_1062;
  wire  T_1064;
  wire  T_1065;
  wire  T_1066;
  wire  T_1067;
  wire  T_1069;
  wire  T_1071;
  wire  GEN_58;
  wire [1:0] GEN_59;
  wire [33:0] GEN_60;
  wire  GEN_61;
  wire [1:0] GEN_62;
  wire [33:0] GEN_63;
  wire  T_1076;
  wire  T_1077;
  wire  GEN_64;
  wire [1:0] GEN_65;
  wire [33:0] GEN_66;
  wire  T_1081;
  wire  T_1082;
  wire  GEN_67;
  wire  GEN_68;
  wire [1:0] GEN_69;
  wire [33:0] GEN_70;
  wire [63:0] T_1113_0;
  wire [63:0] T_1113_1;
  wire [63:0] T_1113_2;
  wire [63:0] T_1113_3;
  wire [63:0] T_1113_4;
  wire [63:0] T_1113_5;
  wire [63:0] T_1113_6;
  wire [63:0] T_1113_7;
  wire [63:0] T_1113_8;
  wire [63:0] T_1113_9;
  wire [63:0] T_1113_10;
  wire [63:0] T_1113_11;
  wire [63:0] T_1113_12;
  wire [63:0] T_1113_13;
  wire [63:0] T_1113_14;
  wire [63:0] T_1113_15;
  wire [63:0] T_1113_16;
  wire [63:0] T_1113_17;
  wire [63:0] T_1113_18;
  wire [63:0] T_1113_19;
  wire [63:0] T_1113_20;
  wire [63:0] T_1113_21;
  wire [63:0] T_1113_22;
  wire [63:0] T_1113_23;
  wire [4:0] T_1116;
  wire [4:0] T_1117;
  wire [63:0] GEN_6;
  wire [4:0] GEN_124;
  wire [63:0] GEN_71;
  wire [4:0] GEN_125;
  wire [63:0] GEN_72;
  wire [4:0] GEN_126;
  wire [63:0] GEN_73;
  wire [4:0] GEN_127;
  wire [63:0] GEN_74;
  wire [4:0] GEN_128;
  wire [63:0] GEN_75;
  wire [4:0] GEN_129;
  wire [63:0] GEN_76;
  wire [4:0] GEN_130;
  wire [63:0] GEN_77;
  wire [4:0] GEN_131;
  wire [63:0] GEN_78;
  wire [4:0] GEN_132;
  wire [63:0] GEN_79;
  wire [4:0] GEN_133;
  wire [63:0] GEN_80;
  wire [4:0] GEN_134;
  wire [63:0] GEN_81;
  wire [4:0] GEN_135;
  wire [63:0] GEN_82;
  wire [4:0] GEN_136;
  wire [63:0] GEN_83;
  wire [4:0] GEN_137;
  wire [63:0] GEN_84;
  wire [4:0] GEN_138;
  wire [63:0] GEN_85;
  wire [63:0] GEN_86;
  wire [63:0] GEN_87;
  wire [63:0] GEN_88;
  wire [63:0] GEN_89;
  wire [63:0] GEN_90;
  wire [63:0] GEN_91;
  wire [63:0] GEN_92;
  wire [63:0] GEN_93;
  wire [31:0] T_1121;
  wire [31:0] T_1122;
  wire [31:0] T_1128_0;
  wire [31:0] T_1128_1;
  wire [31:0] T_1130;
  wire [31:0] T_1131;
  wire [31:0] T_1137_0;
  wire [31:0] T_1137_1;
  wire [31:0] GEN_7;
  wire [31:0] GEN_8;
  wire [3:0] T_1143;
  wire [3:0] GEN_139;
  wire  T_1145;
  wire  GEN_96;
  wire [8:0] T_1146;
  wire  T_1149;
  wire [31:0] GEN_9;
  wire  T_1153;
  wire  T_1154;
  wire  T_1155;
  wire  T_1159;
  wire [31:0] GEN_10;
  wire  T_1163;
  wire  T_1164;
  wire  T_1165;
  wire [63:0] GEN_100;
  wire  GEN_101;
  wire  T_1174;
  wire  T_1177;
  wire  T_1178;
  wire  T_1180;
  wire  T_1181;
  wire [63:0] GEN_102;
  wire  T_1185;
  wire  T_1186;
  wire [63:0] GEN_103;
  reg [25:0] sbAcqReg_addr_block;
  reg [31:0] GEN_153;
  reg [1:0] sbAcqReg_client_xact_id;
  reg [31:0] GEN_154;
  reg [2:0] sbAcqReg_addr_beat;
  reg [31:0] GEN_155;
  reg  sbAcqReg_is_builtin_type;
  reg [31:0] GEN_156;
  reg [2:0] sbAcqReg_a_type;
  reg [31:0] GEN_157;
  reg [11:0] sbAcqReg_union;
  reg [31:0] GEN_158;
  reg [63:0] sbAcqReg_data;
  reg [63:0] GEN_159;
  reg  sbAcqValidReg;
  reg [31:0] GEN_160;
  wire  T_1215;
  wire  sbReg_get;
  wire  T_1216;
  wire  sbReg_getblk;
  wire  T_1217;
  wire  sbReg_put;
  wire  T_1218;
  wire  sbReg_putblk;
  wire  sbMultibeat;
  wire [2:0] GEN_143;
  wire [3:0] T_1220;
  wire [2:0] sbBeatInc1;
  wire  sbLast;
  wire [2:0] T_1222;
  wire [28:0] T_1223;
  wire [31:0] T_1224;
  wire  T_1225;
  wire  T_1226;
  wire  T_1227;
  wire  T_1228;
  wire  T_1230;
  wire  T_1231;
  wire [7:0] GEN_144;
  wire [8:0] T_1235;
  wire [7:0] T_1236;
  wire [7:0] T_1242_0;
  wire  T_1250;
  wire [7:0] T_1251;
  wire [7:0] T_1253;
  wire [7:0] T_1254;
  wire  T_1255;
  wire  T_1256;
  wire  T_1257;
  wire  T_1258;
  wire  T_1259;
  wire  T_1260;
  wire  T_1261;
  wire  T_1262;
  wire [7:0] GEN_145;
  wire [8:0] T_1264;
  wire [7:0] T_1265;
  wire [7:0] GEN_146;
  wire [8:0] T_1267;
  wire [7:0] T_1268;
  wire [7:0] GEN_147;
  wire [8:0] T_1270;
  wire [7:0] T_1271;
  wire [7:0] GEN_148;
  wire [8:0] T_1273;
  wire [7:0] T_1274;
  wire [7:0] GEN_149;
  wire [8:0] T_1276;
  wire [7:0] T_1277;
  wire [7:0] GEN_150;
  wire [8:0] T_1279;
  wire [7:0] T_1280;
  wire [7:0] GEN_151;
  wire [8:0] T_1282;
  wire [7:0] T_1283;
  wire [7:0] GEN_152;
  wire [8:0] T_1285;
  wire [7:0] T_1286;
  wire [7:0] T_1292_0;
  wire [7:0] T_1292_1;
  wire [7:0] T_1292_2;
  wire [7:0] T_1292_3;
  wire [7:0] T_1292_4;
  wire [7:0] T_1292_5;
  wire [7:0] T_1292_6;
  wire [7:0] T_1292_7;
  wire [15:0] T_1294;
  wire [15:0] T_1295;
  wire [31:0] T_1296;
  wire [15:0] T_1297;
  wire [15:0] T_1298;
  wire [31:0] T_1299;
  wire [63:0] T_1300;
  wire  T_1301;
  wire [25:0] GEN_104;
  wire [1:0] GEN_105;
  wire [2:0] GEN_106;
  wire  GEN_107;
  wire [2:0] GEN_108;
  wire [11:0] GEN_109;
  wire [63:0] GEN_110;
  wire  GEN_111;
  wire  T_1303;
  wire  T_1305;
  wire  T_1306;
  wire  GEN_112;
  wire [2:0] GEN_113;
  wire  GEN_114;
  wire  T_1309;
  wire  GEN_115;
  wire [2:0] GEN_116;
  wire  GEN_117;
  wire  T_1327;
  wire [2:0] T_1328;
  wire  T_1329;
  wire [2:0] T_1330;
  wire  T_1331;
  wire [2:0] T_1332;
  wire  T_1333;
  wire [2:0] T_1334;
  wire  T_1335;
  wire [2:0] T_1336;
  wire  T_1337;
  wire [2:0] T_1338;
  wire  T_1339;
  wire [2:0] T_1340;
  wire [2:0] T_1364_addr_beat;
  wire [1:0] T_1364_client_xact_id;
  wire  T_1364_manager_xact_id;
  wire  T_1364_is_builtin_type;
  wire [3:0] T_1364_g_type;
  wire [63:0] T_1364_data;
  wire  T_1389;
  wire  T_1390;
  wire  T_1392;
  wire  T_1393;
  wire  T_1394;
  wire  sbStall;
  wire  T_1396;
  assign io_db_req_ready = T_1067;
  assign io_db_resp_valid = dbStateReg;
  assign io_db_resp_bits_resp = dbRespReg_resp;
  assign io_db_resp_bits_data = dbRespReg_data;
  assign io_debugInterrupts_0 = interruptRegs_0;
  assign io_tl_acquire_ready = T_1396;
  assign io_tl_grant_valid = sbAcqValidReg;
  assign io_tl_grant_bits_addr_beat = T_1364_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1364_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1364_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1364_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1364_g_type;
  assign io_tl_grant_bits_data = T_1364_data;
  assign io_ndreset = ndresetCtrReg;
  assign io_fullreset = CONTROLReg_fullreset;
  assign CONTROLReset_interrupt = 1'h0;
  assign CONTROLReset_haltnot = 1'h0;
  assign CONTROLReset_reserved0 = {{9'd0}, 1'h0};
  assign CONTROLReset_buserror = {{2'd0}, 1'h0};
  assign CONTROLReset_serial = {{2'd0}, 1'h0};
  assign CONTROLReset_autoincrement = 1'h0;
  assign CONTROLReset_access = {{1'd0}, 2'h2};
  assign CONTROLReset_hartid = {{9'd0}, 1'h0};
  assign CONTROLReset_ndreset = 1'h0;
  assign CONTROLReset_fullreset = 1'h0;
  assign CONTROLWrEn = GEN_32;
  assign CONTROLWrData_interrupt = T_878_interrupt;
  assign CONTROLWrData_haltnot = T_878_haltnot;
  assign CONTROLWrData_reserved0 = T_878_reserved0;
  assign CONTROLWrData_buserror = T_878_buserror;
  assign CONTROLWrData_serial = T_878_serial;
  assign CONTROLWrData_autoincrement = T_878_autoincrement;
  assign CONTROLWrData_access = T_878_access;
  assign CONTROLWrData_hartid = T_878_hartid;
  assign CONTROLWrData_ndreset = T_878_ndreset;
  assign CONTROLWrData_fullreset = T_878_fullreset;
  assign CONTROLRdData_interrupt = GEN_2;
  assign CONTROLRdData_haltnot = GEN_3;
  assign CONTROLRdData_reserved0 = CONTROLReg_reserved0;
  assign CONTROLRdData_buserror = CONTROLReg_buserror;
  assign CONTROLRdData_serial = CONTROLReg_serial;
  assign CONTROLRdData_autoincrement = CONTROLReg_autoincrement;
  assign CONTROLRdData_access = CONTROLReg_access;
  assign CONTROLRdData_hartid = CONTROLReg_hartid;
  assign CONTROLRdData_ndreset = ndresetCtrReg;
  assign CONTROLRdData_fullreset = CONTROLReg_fullreset;
  assign DMINFORdData_reserved0 = {{1'd0}, 1'h0};
  assign DMINFORdData_abussize = {{6'd0}, 1'h0};
  assign DMINFORdData_serialcount = {{3'd0}, 1'h0};
  assign DMINFORdData_access128 = 1'h0;
  assign DMINFORdData_access64 = 1'h0;
  assign DMINFORdData_access32 = 1'h0;
  assign DMINFORdData_access16 = 1'h0;
  assign DMINFORdData_accesss8 = 1'h0;
  assign DMINFORdData_dramsize = {{2'd0}, 4'hf};
  assign DMINFORdData_haltsum = 1'h0;
  assign DMINFORdData_reserved1 = {{2'd0}, 1'h0};
  assign DMINFORdData_authenticated = 1'h1;
  assign DMINFORdData_authbusy = 1'h0;
  assign DMINFORdData_authtype = {{1'd0}, 1'h0};
  assign DMINFORdData_version = {{1'd0}, 1'h1};
  assign HALTSUMRdData_serialfull = 1'h0;
  assign HALTSUMRdData_serialvalid = 1'h0;
  assign HALTSUMRdData_acks = {{31'd0}, haltnotSummary};
  assign RAMWrData_interrupt = T_907_interrupt;
  assign RAMWrData_haltnot = T_907_haltnot;
  assign RAMWrData_data = T_907_data;
  assign RAMRdData_interrupt = GEN_4;
  assign RAMRdData_haltnot = GEN_5;
  assign RAMRdData_data = dbRamRdData;
  assign SETHALTNOTWrEn = T_1155;
  assign SETHALTNOTWrData = GEN_7[9:0];
  assign CLEARDEBINTWrEn = T_1165;
  assign CLEARDEBINTWrData = GEN_8[9:0];
  assign T_655_0 = 1'h0;
  assign T_666_0 = 1'h0;
  assign haltnotStatus_0 = {{31'd0}, haltnotRegs_0};
  assign rdHaltnotStatus = GEN_50;
  assign GEN_118 = {{31'd0}, 1'h0};
  assign haltnotSummary = haltnotStatus_0 != GEN_118;
  assign ramMem_T_853_addr = ramAddr;
  assign ramMem_T_853_en = 1'h1;
  `ifdef SYNTHESIS
  assign ramMem_T_853_data = ramMem[ramMem_T_853_addr];
  `else
  assign ramMem_T_853_data = ramMem_T_853_addr >= 4'h8 ? $random : ramMem[ramMem_T_853_addr];
  `endif
  assign ramMem_T_854_data = ramWrData;
  assign ramMem_T_854_addr = ramAddr;
  assign ramMem_T_854_mask = ramWrEn;
  assign ramMem_T_854_en = ramWrEn;
  assign ramAddr = T_852;
  assign ramRdData = ramMem_T_853_data;
  assign ramWrData = T_849;
  assign ramWrMask = T_832;
  assign ramWrEn = T_855;
  assign dbRamAddr = T_782;
  assign dbRamRdData = GEN_1;
  assign dbRamWrData = dbReq_data[31:0];
  assign dbRamWrEn = GEN_31;
  assign dbRamRdEn = 1'h0;
  assign sbRamAddr = T_783;
  assign sbRamRdData = ramRdData;
  assign sbRamWrData = sbWrData;
  assign sbRamWrEn = GEN_96;
  assign sbRamRdEn = GEN_101;
  assign sbRomRdData = GEN_6;
  assign dbRdEn = T_1069;
  assign dbWrEn = T_1071;
  assign dbRdData = GEN_57;
  assign dbResult_resp = T_1059;
  assign dbResult_data = dbRdData;
  assign dbReq_addr = io_db_req_bits_addr;
  assign dbReq_op = io_db_req_bits_op;
  assign dbReq_data = io_db_req_bits_data;
  assign rdCondWrFailure = T_1049;
  assign dbWrNeeded = T_1056;
  assign sbAddr = T_1224[11:0];
  assign sbRdData = GEN_103;
  assign sbWrData = sbAcqReg_data;
  assign sbWrMask = T_1300;
  assign sbWrEn = T_1228;
  assign sbRdEn = T_1226;
  assign stallFromDb = 1'h0;
  assign stallFromSb = T_834;
  assign GEN_119 = {{9'd0}, 1'h0};
  assign T_720 = CONTROLWrData_hartid == GEN_119;
  assign T_721 = interruptRegs_0 | CONTROLWrData_interrupt;
  assign GEN_11 = T_720 ? T_721 : interruptRegs_0;
  assign GEN_12 = CONTROLWrEn ? GEN_11 : interruptRegs_0;
  assign T_723 = CONTROLWrEn == 1'h0;
  assign T_724 = T_723 & dbRamWrEn;
  assign T_726 = CONTROLReg_hartid == GEN_119;
  assign T_727 = interruptRegs_0 | RAMWrData_interrupt;
  assign GEN_13 = T_726 ? T_727 : GEN_12;
  assign GEN_14 = T_724 ? GEN_13 : GEN_12;
  assign T_731 = dbRamWrEn == 1'h0;
  assign T_732 = T_723 & T_731;
  assign T_733 = T_732 & CLEARDEBINTWrEn;
  assign T_735 = CLEARDEBINTWrData == 10'h0;
  assign GEN_15 = T_735 ? 1'h0 : GEN_14;
  assign GEN_16 = T_733 ? GEN_15 : GEN_14;
  assign T_738 = SETHALTNOTWrData == 10'h0;
  assign GEN_17 = T_738 ? 1'h1 : haltnotRegs_0;
  assign GEN_18 = SETHALTNOTWrEn ? GEN_17 : haltnotRegs_0;
  assign T_741 = SETHALTNOTWrEn == 1'h0;
  assign T_742 = T_741 & CONTROLWrEn;
  assign T_745 = haltnotRegs_0 & CONTROLWrData_haltnot;
  assign GEN_19 = T_720 ? T_745 : GEN_18;
  assign GEN_20 = T_742 ? GEN_19 : GEN_18;
  assign T_750 = T_741 & T_723;
  assign T_751 = T_750 & dbRamWrEn;
  assign T_754 = haltnotRegs_0 & RAMWrData_haltnot;
  assign GEN_21 = T_726 ? T_754 : GEN_20;
  assign GEN_22 = T_751 ? GEN_21 : GEN_20;
  assign T_782 = dbReq_addr[3:0];
  assign T_783 = sbAddr[5:3];
  assign T_801_0 = 32'hffffffff;
  assign T_801_1 = 32'hffffffff;
  assign dbRamWrMask_0 = GEN_23;
  assign dbRamWrMask_1 = GEN_24;
  assign T_806 = dbRamAddr[0];
  assign T_807 = ramRdData[31:0];
  assign T_808 = ramRdData[63:32];
  assign T_814_0 = T_807;
  assign T_814_1 = T_808;
  assign T_823_0 = 32'h0;
  assign T_823_1 = 32'h0;
  assign GEN_0 = 32'hffffffff;
  assign GEN_23 = 1'h0 == T_806 ? GEN_0 : T_823_0;
  assign GEN_24 = T_806 ? GEN_0 : T_823_1;
  assign GEN_1 = GEN_25;
  assign GEN_25 = T_806 ? T_814_1 : T_814_0;
  assign T_831 = {dbRamWrMask_1,dbRamWrMask_0};
  assign T_832 = sbRamWrEn ? sbWrMask : T_831;
  assign T_833 = dbRamWrEn | dbRamRdEn;
  assign T_834 = sbRamRdEn | sbRamWrEn;
  assign T_835 = T_833 & T_834;
  assign T_837 = T_835 == 1'h0;
  assign T_838 = T_837 | reset;
  assign T_840 = T_838 == 1'h0;
  assign dbRamWrDataVec = {dbRamWrData,dbRamWrData};
  assign T_841 = ramWrMask & sbRamWrData;
  assign T_842 = ~ ramWrMask;
  assign T_843 = T_842 & ramRdData;
  assign T_844 = T_841 | T_843;
  assign T_845 = ramWrMask & dbRamWrDataVec;
  assign T_848 = T_845 | T_843;
  assign T_849 = sbRamWrEn ? T_844 : T_848;
  assign T_850 = sbRamWrEn | sbRamRdEn;
  assign T_851 = dbRamAddr[3:1];
  assign T_852 = T_850 ? sbRamAddr : T_851;
  assign T_855 = sbRamWrEn | dbRamWrEn;
  assign T_878_interrupt = T_898;
  assign T_878_haltnot = T_897;
  assign T_878_reserved0 = T_896;
  assign T_878_buserror = T_895;
  assign T_878_serial = T_894;
  assign T_878_autoincrement = T_893;
  assign T_878_access = T_892;
  assign T_878_hartid = T_891;
  assign T_878_ndreset = T_890;
  assign T_878_fullreset = T_889;
  assign T_889 = dbReq_data[0];
  assign T_890 = dbReq_data[1];
  assign T_891 = dbReq_data[11:2];
  assign T_892 = dbReq_data[14:12];
  assign T_893 = dbReq_data[15];
  assign T_894 = dbReq_data[18:16];
  assign T_895 = dbReq_data[21:19];
  assign T_896 = dbReq_data[31:22];
  assign T_897 = dbReq_data[32];
  assign T_898 = dbReq_data[33];
  assign T_907_interrupt = T_898;
  assign T_907_haltnot = T_897;
  assign T_907_data = T_911;
  assign T_911 = dbReq_data[31:0];
  assign T_916 = dbReq_addr[4:4];
  assign T_918 = T_916 == 1'h0;
  assign GEN_31 = T_918 ? dbWrEn : 1'h0;
  assign T_920 = dbReq_addr == 5'h10;
  assign T_922 = T_918 == 1'h0;
  assign T_923 = T_922 & T_920;
  assign GEN_32 = T_923 ? dbWrEn : 1'h0;
  assign T_927 = T_920 == 1'h0;
  assign T_928 = T_922 & T_927;
  assign GEN_33 = reset ? CONTROLReset_interrupt : CONTROLReg_interrupt;
  assign GEN_34 = reset ? CONTROLReset_haltnot : CONTROLReg_haltnot;
  assign GEN_35 = reset ? CONTROLReset_reserved0 : CONTROLReg_reserved0;
  assign GEN_36 = reset ? CONTROLReset_buserror : CONTROLReg_buserror;
  assign GEN_37 = reset ? CONTROLReset_serial : CONTROLReg_serial;
  assign GEN_38 = reset ? CONTROLReset_autoincrement : CONTROLReg_autoincrement;
  assign GEN_39 = reset ? CONTROLReset_access : CONTROLReg_access;
  assign GEN_40 = reset ? CONTROLReset_hartid : CONTROLReg_hartid;
  assign GEN_41 = reset ? CONTROLReset_ndreset : CONTROLReg_ndreset;
  assign GEN_42 = reset ? CONTROLReset_fullreset : CONTROLReg_fullreset;
  assign GEN_43 = reset ? 1'h0 : ndresetCtrReg;
  assign T_931 = reset == 1'h0;
  assign T_932 = T_931 & CONTROLWrEn;
  assign T_933 = CONTROLReg_fullreset | CONTROLWrData_fullreset;
  assign GEN_44 = CONTROLWrData_ndreset ? 1'h1 : GEN_43;
  assign T_936 = CONTROLWrData_ndreset == 1'h0;
  assign T_938 = ndresetCtrReg == 1'h0;
  assign T_941 = ndresetCtrReg - 1'h1;
  assign T_942 = T_941[0:0];
  assign T_943 = T_938 ? 1'h0 : T_942;
  assign GEN_45 = T_936 ? T_943 : GEN_44;
  assign GEN_46 = T_932 ? CONTROLWrData_hartid : GEN_40;
  assign GEN_47 = T_932 ? T_933 : GEN_42;
  assign GEN_48 = T_932 ? GEN_45 : GEN_43;
  assign T_948 = T_931 & T_723;
  assign GEN_49 = T_948 ? T_943 : GEN_48;
  assign GEN_2 = interruptRegs_0;
  assign GEN_3 = haltnotRegs_0;
  assign GEN_4 = interruptRegs_0;
  assign GEN_5 = haltnotRegs_0;
  assign GEN_123 = {{4'd0}, 1'h0};
  assign T_961 = dbReq_addr == GEN_123;
  assign GEN_50 = T_961 ? haltnotStatus_0 : {{31'd0}, 1'h0};
  assign T_966 = {RAMRdData_interrupt,RAMRdData_haltnot};
  assign T_967 = {T_966,RAMRdData_data};
  assign GEN_51 = T_918 ? T_967 : {{33'd0}, 1'h0};
  assign T_973 = {CONTROLRdData_ndreset,CONTROLRdData_fullreset};
  assign T_974 = {CONTROLRdData_autoincrement,CONTROLRdData_access};
  assign T_975 = {T_974,CONTROLRdData_hartid};
  assign T_976 = {T_975,T_973};
  assign T_977 = {CONTROLRdData_buserror,CONTROLRdData_serial};
  assign T_978 = {CONTROLRdData_interrupt,CONTROLRdData_haltnot};
  assign T_979 = {T_978,CONTROLRdData_reserved0};
  assign T_980 = {T_979,T_977};
  assign T_981 = {T_980,T_976};
  assign GEN_53 = T_923 ? T_981 : GEN_51;
  assign T_983 = dbReq_addr == 5'h11;
  assign T_989 = T_928 & T_983;
  assign T_990 = {DMINFORdData_authbusy,DMINFORdData_authtype};
  assign T_991 = {T_990,DMINFORdData_version};
  assign T_992 = {DMINFORdData_reserved1,DMINFORdData_authenticated};
  assign T_993 = {DMINFORdData_dramsize,DMINFORdData_haltsum};
  assign T_994 = {T_993,T_992};
  assign T_995 = {T_994,T_991};
  assign T_996 = {DMINFORdData_access16,DMINFORdData_accesss8};
  assign T_997 = {DMINFORdData_access64,DMINFORdData_access32};
  assign T_998 = {T_997,T_996};
  assign T_999 = {DMINFORdData_serialcount,DMINFORdData_access128};
  assign T_1000 = {DMINFORdData_reserved0,DMINFORdData_abussize};
  assign T_1001 = {T_1000,T_999};
  assign T_1002 = {T_1001,T_998};
  assign T_1003 = {T_1002,T_995};
  assign GEN_54 = T_989 ? T_1003 : GEN_53;
  assign T_1005 = dbReq_addr == 5'h1b;
  assign T_1012 = T_983 == 1'h0;
  assign T_1013 = T_928 & T_1012;
  assign T_1014 = T_1013 & T_1005;
  assign GEN_55 = T_1014 ? {{33'd0}, 1'h0} : GEN_54;
  assign T_1016 = dbReq_addr[4:2];
  assign T_1018 = T_1016 == 3'h7;
  assign T_1028 = T_1005 == 1'h0;
  assign T_1029 = T_1013 & T_1028;
  assign T_1030 = T_1029 & T_1018;
  assign GEN_56 = T_1030 ? {{2'd0}, rdHaltnotStatus} : GEN_55;
  assign T_1043 = T_1018 == 1'h0;
  assign T_1044 = T_1029 & T_1043;
  assign GEN_57 = T_1044 ? {{33'd0}, 1'h0} : GEN_56;
  assign T_1046 = dbRdData[33];
  assign T_1048 = dbReq_op == 2'h3;
  assign T_1049 = T_1046 & T_1048;
  assign T_1051 = dbReq_op == 2'h2;
  assign T_1054 = ~ rdCondWrFailure;
  assign T_1055 = T_1048 & T_1054;
  assign T_1056 = T_1051 | T_1055;
  assign T_1059 = rdCondWrFailure ? 2'h1 : 2'h0;
  assign T_1061 = stallFromSb == 1'h0;
  assign T_1062 = dbStateReg == 1'h0;
  assign T_1064 = io_db_resp_ready & io_db_resp_valid;
  assign T_1065 = dbStateReg & T_1064;
  assign T_1066 = T_1062 | T_1065;
  assign T_1067 = T_1061 & T_1066;
  assign T_1069 = io_db_req_ready & io_db_req_valid;
  assign T_1071 = dbWrNeeded & T_1069;
  assign GEN_58 = T_1069 ? 1'h1 : dbStateReg;
  assign GEN_59 = T_1069 ? dbResult_resp : dbRespReg_resp;
  assign GEN_60 = T_1069 ? dbResult_data : dbRespReg_data;
  assign GEN_61 = T_1062 ? GEN_58 : dbStateReg;
  assign GEN_62 = T_1062 ? GEN_59 : dbRespReg_resp;
  assign GEN_63 = T_1062 ? GEN_60 : dbRespReg_data;
  assign T_1076 = T_1062 == 1'h0;
  assign T_1077 = T_1076 & dbStateReg;
  assign GEN_64 = T_1069 ? 1'h1 : GEN_61;
  assign GEN_65 = T_1069 ? dbResult_resp : GEN_62;
  assign GEN_66 = T_1069 ? dbResult_data : GEN_63;
  assign T_1081 = T_1069 == 1'h0;
  assign T_1082 = T_1081 & T_1064;
  assign GEN_67 = T_1082 ? 1'h0 : GEN_64;
  assign GEN_68 = T_1077 ? GEN_67 : GEN_61;
  assign GEN_69 = T_1077 ? GEN_65 : GEN_62;
  assign GEN_70 = T_1077 ? GEN_66 : GEN_63;
  assign T_1113_0 = 64'hc0006f0600006f;
  assign T_1113_1 = 64'h80006ffff00413;
  assign T_1113_2 = 64'hff0000f00000413;
  assign T_1113_3 = 64'h4c663f10024f3;
  assign T_1113_4 = 64'h180006f43c02483;
  assign T_1113_5 = 64'h4c66300149493;
  assign T_1113_6 = 64'h80006f43803483;
  assign T_1113_7 = 64'h42802e2300000013;
  assign T_1113_8 = 64'h10802023f1402473;
  assign T_1113_9 = 64'h8474137b002473;
  assign T_1113_10 = 64'h580006f00040463;
  assign T_1113_11 = 64'h7b2000737b202473;
  assign T_1113_12 = 64'h7b0024737b241073;
  assign T_1113_13 = 64'hf40404131c047413;
  assign T_1113_14 = 64'h100f02041863;
  assign T_1113_15 = 64'h44663f1002473;
  assign T_1113_16 = 64'h4000006742902e23;
  assign T_1113_17 = 64'h4466300141413;
  assign T_1113_18 = 64'h4000006742903c23;
  assign T_1113_19 = 64'h4000006700000013;
  assign T_1113_20 = 64'h10802623f1402473;
  assign T_1113_21 = 64'h7b0024737b046073;
  assign T_1113_22 = 64'hfe040ce302047413;
  assign T_1113_23 = 64'hfbdff06f;
  assign T_1116 = T_1117;
  assign T_1117 = sbAddr[7:3];
  assign GEN_6 = GEN_93;
  assign GEN_124 = {{4'd0}, 1'h1};
  assign GEN_71 = GEN_124 == T_1116 ? T_1113_1 : T_1113_0;
  assign GEN_125 = {{3'd0}, 2'h2};
  assign GEN_72 = GEN_125 == T_1116 ? T_1113_2 : GEN_71;
  assign GEN_126 = {{3'd0}, 2'h3};
  assign GEN_73 = GEN_126 == T_1116 ? T_1113_3 : GEN_72;
  assign GEN_127 = {{2'd0}, 3'h4};
  assign GEN_74 = GEN_127 == T_1116 ? T_1113_4 : GEN_73;
  assign GEN_128 = {{2'd0}, 3'h5};
  assign GEN_75 = GEN_128 == T_1116 ? T_1113_5 : GEN_74;
  assign GEN_129 = {{2'd0}, 3'h6};
  assign GEN_76 = GEN_129 == T_1116 ? T_1113_6 : GEN_75;
  assign GEN_130 = {{2'd0}, 3'h7};
  assign GEN_77 = GEN_130 == T_1116 ? T_1113_7 : GEN_76;
  assign GEN_131 = {{1'd0}, 4'h8};
  assign GEN_78 = GEN_131 == T_1116 ? T_1113_8 : GEN_77;
  assign GEN_132 = {{1'd0}, 4'h9};
  assign GEN_79 = GEN_132 == T_1116 ? T_1113_9 : GEN_78;
  assign GEN_133 = {{1'd0}, 4'ha};
  assign GEN_80 = GEN_133 == T_1116 ? T_1113_10 : GEN_79;
  assign GEN_134 = {{1'd0}, 4'hb};
  assign GEN_81 = GEN_134 == T_1116 ? T_1113_11 : GEN_80;
  assign GEN_135 = {{1'd0}, 4'hc};
  assign GEN_82 = GEN_135 == T_1116 ? T_1113_12 : GEN_81;
  assign GEN_136 = {{1'd0}, 4'hd};
  assign GEN_83 = GEN_136 == T_1116 ? T_1113_13 : GEN_82;
  assign GEN_137 = {{1'd0}, 4'he};
  assign GEN_84 = GEN_137 == T_1116 ? T_1113_14 : GEN_83;
  assign GEN_138 = {{1'd0}, 4'hf};
  assign GEN_85 = GEN_138 == T_1116 ? T_1113_15 : GEN_84;
  assign GEN_86 = 5'h10 == T_1116 ? T_1113_16 : GEN_85;
  assign GEN_87 = 5'h11 == T_1116 ? T_1113_17 : GEN_86;
  assign GEN_88 = 5'h12 == T_1116 ? T_1113_18 : GEN_87;
  assign GEN_89 = 5'h13 == T_1116 ? T_1113_19 : GEN_88;
  assign GEN_90 = 5'h14 == T_1116 ? T_1113_20 : GEN_89;
  assign GEN_91 = 5'h15 == T_1116 ? T_1113_21 : GEN_90;
  assign GEN_92 = 5'h16 == T_1116 ? T_1113_22 : GEN_91;
  assign GEN_93 = 5'h17 == T_1116 ? T_1113_23 : GEN_92;
  assign T_1121 = sbWrData[31:0];
  assign T_1122 = sbWrData[63:32];
  assign T_1128_0 = T_1121;
  assign T_1128_1 = T_1122;
  assign T_1130 = sbWrMask[31:0];
  assign T_1131 = sbWrMask[63:32];
  assign T_1137_0 = T_1130;
  assign T_1137_1 = T_1131;
  assign GEN_7 = T_1128_1;
  assign GEN_8 = T_1128_0;
  assign T_1143 = sbAddr[11:8];
  assign GEN_139 = {{1'd0}, 3'h4};
  assign T_1145 = T_1143 == GEN_139;
  assign GEN_96 = T_1145 ? sbWrEn : 1'h0;
  assign T_1146 = sbAddr[11:3];
  assign T_1149 = T_1146 == 9'h21;
  assign GEN_9 = T_1137_1;
  assign T_1153 = GEN_9 != GEN_118;
  assign T_1154 = T_1149 & T_1153;
  assign T_1155 = T_1154 & sbWrEn;
  assign T_1159 = T_1146 == 9'h20;
  assign GEN_10 = T_1137_0;
  assign T_1163 = GEN_10 != GEN_118;
  assign T_1164 = T_1159 & T_1163;
  assign T_1165 = T_1164 & sbWrEn;
  assign GEN_100 = T_1145 ? sbRamRdData : {{63'd0}, 1'h0};
  assign GEN_101 = T_1145 ? sbRdEn : 1'h0;
  assign T_1174 = T_1143 == 4'h8;
  assign T_1177 = T_1143 == 4'h9;
  assign T_1178 = T_1174 | T_1177;
  assign T_1180 = T_1145 == 1'h0;
  assign T_1181 = T_1180 & T_1178;
  assign GEN_102 = T_1181 ? sbRomRdData : GEN_100;
  assign T_1185 = T_1178 == 1'h0;
  assign T_1186 = T_1180 & T_1185;
  assign GEN_103 = T_1186 ? {{63'd0}, 1'h0} : GEN_102;
  assign T_1215 = sbAcqReg_a_type == 3'h0;
  assign sbReg_get = sbAcqReg_is_builtin_type & T_1215;
  assign T_1216 = sbAcqReg_a_type == 3'h1;
  assign sbReg_getblk = sbAcqReg_is_builtin_type & T_1216;
  assign T_1217 = sbAcqReg_a_type == 3'h2;
  assign sbReg_put = sbAcqReg_is_builtin_type & T_1217;
  assign T_1218 = sbAcqReg_a_type == 3'h3;
  assign sbReg_putblk = sbAcqReg_is_builtin_type & T_1218;
  assign sbMultibeat = sbReg_getblk & sbAcqValidReg;
  assign GEN_143 = {{2'd0}, 1'h1};
  assign T_1220 = sbAcqReg_addr_beat + GEN_143;
  assign sbBeatInc1 = T_1220[2:0];
  assign sbLast = sbAcqReg_addr_beat == 3'h7;
  assign T_1222 = sbAcqReg_union[11:9];
  assign T_1223 = {sbAcqReg_addr_block,sbAcqReg_addr_beat};
  assign T_1224 = {T_1223,T_1222};
  assign T_1225 = sbReg_get | sbReg_getblk;
  assign T_1226 = sbAcqValidReg & T_1225;
  assign T_1227 = sbReg_put | sbReg_putblk;
  assign T_1228 = sbAcqValidReg & T_1227;
  assign T_1230 = sbAcqReg_a_type == 3'h4;
  assign T_1231 = sbAcqReg_is_builtin_type & T_1230;
  assign GEN_144 = {{7'd0}, 1'h1};
  assign T_1235 = 8'h0 - GEN_144;
  assign T_1236 = T_1235[7:0];
  assign T_1242_0 = T_1236;
  assign T_1250 = sbReg_putblk | sbReg_put;
  assign T_1251 = sbAcqReg_union[8:1];
  assign T_1253 = T_1250 ? T_1251 : {{7'd0}, 1'h0};
  assign T_1254 = T_1231 ? T_1242_0 : T_1253;
  assign T_1255 = T_1254[0];
  assign T_1256 = T_1254[1];
  assign T_1257 = T_1254[2];
  assign T_1258 = T_1254[3];
  assign T_1259 = T_1254[4];
  assign T_1260 = T_1254[5];
  assign T_1261 = T_1254[6];
  assign T_1262 = T_1254[7];
  assign GEN_145 = {{7'd0}, T_1255};
  assign T_1264 = 8'h0 - GEN_145;
  assign T_1265 = T_1264[7:0];
  assign GEN_146 = {{7'd0}, T_1256};
  assign T_1267 = 8'h0 - GEN_146;
  assign T_1268 = T_1267[7:0];
  assign GEN_147 = {{7'd0}, T_1257};
  assign T_1270 = 8'h0 - GEN_147;
  assign T_1271 = T_1270[7:0];
  assign GEN_148 = {{7'd0}, T_1258};
  assign T_1273 = 8'h0 - GEN_148;
  assign T_1274 = T_1273[7:0];
  assign GEN_149 = {{7'd0}, T_1259};
  assign T_1276 = 8'h0 - GEN_149;
  assign T_1277 = T_1276[7:0];
  assign GEN_150 = {{7'd0}, T_1260};
  assign T_1279 = 8'h0 - GEN_150;
  assign T_1280 = T_1279[7:0];
  assign GEN_151 = {{7'd0}, T_1261};
  assign T_1282 = 8'h0 - GEN_151;
  assign T_1283 = T_1282[7:0];
  assign GEN_152 = {{7'd0}, T_1262};
  assign T_1285 = 8'h0 - GEN_152;
  assign T_1286 = T_1285[7:0];
  assign T_1292_0 = T_1265;
  assign T_1292_1 = T_1268;
  assign T_1292_2 = T_1271;
  assign T_1292_3 = T_1274;
  assign T_1292_4 = T_1277;
  assign T_1292_5 = T_1280;
  assign T_1292_6 = T_1283;
  assign T_1292_7 = T_1286;
  assign T_1294 = {T_1292_1,T_1292_0};
  assign T_1295 = {T_1292_3,T_1292_2};
  assign T_1296 = {T_1295,T_1294};
  assign T_1297 = {T_1292_5,T_1292_4};
  assign T_1298 = {T_1292_7,T_1292_6};
  assign T_1299 = {T_1298,T_1297};
  assign T_1300 = {T_1299,T_1296};
  assign T_1301 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign GEN_104 = T_1301 ? io_tl_acquire_bits_addr_block : sbAcqReg_addr_block;
  assign GEN_105 = T_1301 ? io_tl_acquire_bits_client_xact_id : sbAcqReg_client_xact_id;
  assign GEN_106 = T_1301 ? io_tl_acquire_bits_addr_beat : sbAcqReg_addr_beat;
  assign GEN_107 = T_1301 ? io_tl_acquire_bits_is_builtin_type : sbAcqReg_is_builtin_type;
  assign GEN_108 = T_1301 ? io_tl_acquire_bits_a_type : sbAcqReg_a_type;
  assign GEN_109 = T_1301 ? io_tl_acquire_bits_union : sbAcqReg_union;
  assign GEN_110 = T_1301 ? io_tl_acquire_bits_data : sbAcqReg_data;
  assign GEN_111 = T_1301 ? 1'h1 : sbAcqValidReg;
  assign T_1303 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_1305 = T_1301 == 1'h0;
  assign T_1306 = T_1305 & T_1303;
  assign GEN_112 = sbLast ? 1'h0 : GEN_111;
  assign GEN_113 = sbMultibeat ? sbBeatInc1 : GEN_106;
  assign GEN_114 = sbMultibeat ? GEN_112 : GEN_111;
  assign T_1309 = sbMultibeat == 1'h0;
  assign GEN_115 = T_1309 ? 1'h0 : GEN_114;
  assign GEN_116 = T_1306 ? GEN_113 : GEN_106;
  assign GEN_117 = T_1306 ? GEN_115 : GEN_111;
  assign T_1327 = 3'h6 == sbAcqReg_a_type;
  assign T_1328 = T_1327 ? 3'h1 : 3'h3;
  assign T_1329 = 3'h5 == sbAcqReg_a_type;
  assign T_1330 = T_1329 ? 3'h1 : T_1328;
  assign T_1331 = 3'h4 == sbAcqReg_a_type;
  assign T_1332 = T_1331 ? 3'h4 : T_1330;
  assign T_1333 = 3'h3 == sbAcqReg_a_type;
  assign T_1334 = T_1333 ? 3'h3 : T_1332;
  assign T_1335 = 3'h2 == sbAcqReg_a_type;
  assign T_1336 = T_1335 ? 3'h3 : T_1334;
  assign T_1337 = 3'h1 == sbAcqReg_a_type;
  assign T_1338 = T_1337 ? 3'h5 : T_1336;
  assign T_1339 = 3'h0 == sbAcqReg_a_type;
  assign T_1340 = T_1339 ? 3'h4 : T_1338;
  assign T_1364_addr_beat = sbAcqReg_addr_beat;
  assign T_1364_client_xact_id = sbAcqReg_client_xact_id;
  assign T_1364_manager_xact_id = 1'h0;
  assign T_1364_is_builtin_type = 1'h1;
  assign T_1364_g_type = {{1'd0}, T_1340};
  assign T_1364_data = sbRdData;
  assign T_1389 = sbLast == 1'h0;
  assign T_1390 = sbMultibeat & T_1389;
  assign T_1392 = io_tl_grant_ready == 1'h0;
  assign T_1393 = io_tl_grant_valid & T_1392;
  assign T_1394 = T_1390 | T_1393;
  assign sbStall = T_1394 | stallFromDb;
  assign T_1396 = sbStall == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_26 = {1{$random}};
  CONTROLReg_interrupt = GEN_26[0:0];
  GEN_27 = {1{$random}};
  CONTROLReg_haltnot = GEN_27[0:0];
  GEN_28 = {1{$random}};
  CONTROLReg_reserved0 = GEN_28[9:0];
  GEN_29 = {1{$random}};
  CONTROLReg_buserror = GEN_29[2:0];
  GEN_30 = {1{$random}};
  CONTROLReg_serial = GEN_30[2:0];
  GEN_52 = {1{$random}};
  CONTROLReg_autoincrement = GEN_52[0:0];
  GEN_94 = {1{$random}};
  CONTROLReg_access = GEN_94[2:0];
  GEN_95 = {1{$random}};
  CONTROLReg_hartid = GEN_95[9:0];
  GEN_97 = {1{$random}};
  CONTROLReg_ndreset = GEN_97[0:0];
  GEN_98 = {1{$random}};
  CONTROLReg_fullreset = GEN_98[0:0];
  GEN_99 = {1{$random}};
  ndresetCtrReg = GEN_99[0:0];
  GEN_120 = {1{$random}};
  interruptRegs_0 = GEN_120[0:0];
  GEN_121 = {1{$random}};
  haltnotRegs_0 = GEN_121[0:0];
  GEN_122 = {2{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    ramMem[initvar] = GEN_122[63:0];
  GEN_140 = {1{$random}};
  dbStateReg = GEN_140[0:0];
  GEN_141 = {1{$random}};
  dbRespReg_resp = GEN_141[1:0];
  GEN_142 = {2{$random}};
  dbRespReg_data = GEN_142[33:0];
  GEN_153 = {1{$random}};
  sbAcqReg_addr_block = GEN_153[25:0];
  GEN_154 = {1{$random}};
  sbAcqReg_client_xact_id = GEN_154[1:0];
  GEN_155 = {1{$random}};
  sbAcqReg_addr_beat = GEN_155[2:0];
  GEN_156 = {1{$random}};
  sbAcqReg_is_builtin_type = GEN_156[0:0];
  GEN_157 = {1{$random}};
  sbAcqReg_a_type = GEN_157[2:0];
  GEN_158 = {1{$random}};
  sbAcqReg_union = GEN_158[11:0];
  GEN_159 = {2{$random}};
  sbAcqReg_data = GEN_159[63:0];
  GEN_160 = {1{$random}};
  sbAcqValidReg = GEN_160[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      CONTROLReg_interrupt <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_haltnot <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_reserved0 <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_buserror <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_serial <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_autoincrement <= GEN_38;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_access <= GEN_39;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_hartid <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_ndreset <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      CONTROLReg_fullreset <= GEN_47;
    end
    if(1'h0) begin
    end else begin
      ndresetCtrReg <= GEN_49;
    end
    if(reset) begin
      interruptRegs_0 <= T_655_0;
    end else begin
      interruptRegs_0 <= GEN_16;
    end
    if(reset) begin
      haltnotRegs_0 <= T_666_0;
    end else begin
      haltnotRegs_0 <= GEN_22;
    end
    if(ramMem_T_854_en & ramMem_T_854_mask) begin
      ramMem[ramMem_T_854_addr] <= ramMem_T_854_data;
    end
    if(reset) begin
      dbStateReg <= 1'h0;
    end else begin
      dbStateReg <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      dbRespReg_resp <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      dbRespReg_data <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_addr_block <= GEN_104;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_client_xact_id <= GEN_105;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_addr_beat <= GEN_116;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_is_builtin_type <= GEN_107;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_a_type <= GEN_108;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_union <= GEN_109;
    end
    if(1'h0) begin
    end else begin
      sbAcqReg_data <= GEN_110;
    end
    if(reset) begin
      sbAcqValidReg <= 1'h0;
    end else begin
      sbAcqValidReg <= GEN_117;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_840) begin
          $fwrite(32'h80000002,"Assertion failed: Stall logic should have prevented concurrent SB/DB RAM Access\n    at debug.scala:623 assert (!((dbRamWrEn | dbRamRdEn) & (sbRamRdEn | sbRamWrEn)), \"Stall logic should have prevented concurrent SB/DB RAM Access\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_840) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module PRCI(
  input   clk,
  input   reset,
  input   io_interrupts_0_mtip,
  input   io_interrupts_0_meip,
  input   io_interrupts_0_seip,
  input   io_interrupts_0_debug,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  output  io_tiles_0_reset,
  output  io_tiles_0_id,
  output  io_tiles_0_interrupts_mtip,
  output  io_tiles_0_interrupts_meip,
  output  io_tiles_0_interrupts_seip,
  output  io_tiles_0_interrupts_debug,
  output  io_tiles_0_interrupts_msip
);
  wire  T_529_0;
  reg  ipi_0;
  reg [31:0] GEN_2;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_562;
  wire  write;
  wire [31:0] rdata;
  wire  T_565;
  wire  T_566;
  wire [7:0] GEN_5;
  wire [8:0] T_570;
  wire [7:0] T_571;
  wire [7:0] T_577_0;
  wire  T_580;
  wire  T_581;
  wire  T_585;
  wire [7:0] T_586;
  wire [7:0] T_588;
  wire [7:0] T_589;
  wire  T_590;
  wire  T_591;
  wire  T_592;
  wire  T_593;
  wire  T_594;
  wire  T_595;
  wire  T_596;
  wire  T_597;
  wire [7:0] GEN_6;
  wire [8:0] T_599;
  wire [7:0] T_600;
  wire [7:0] GEN_7;
  wire [8:0] T_602;
  wire [7:0] T_603;
  wire [7:0] GEN_8;
  wire [8:0] T_605;
  wire [7:0] T_606;
  wire [7:0] GEN_9;
  wire [8:0] T_608;
  wire [7:0] T_609;
  wire [7:0] GEN_10;
  wire [8:0] T_611;
  wire [7:0] T_612;
  wire [7:0] GEN_11;
  wire [8:0] T_614;
  wire [7:0] T_615;
  wire [7:0] GEN_12;
  wire [8:0] T_617;
  wire [7:0] T_618;
  wire [7:0] GEN_13;
  wire [8:0] T_620;
  wire [7:0] T_621;
  wire [7:0] T_627_0;
  wire [7:0] T_627_1;
  wire [7:0] T_627_2;
  wire [7:0] T_627_3;
  wire [7:0] T_627_4;
  wire [7:0] T_627_5;
  wire [7:0] T_627_6;
  wire [7:0] T_627_7;
  wire [15:0] T_629;
  wire [15:0] T_630;
  wire [31:0] T_631;
  wire [15:0] T_632;
  wire [15:0] T_633;
  wire [31:0] T_634;
  wire [63:0] T_635;
  wire [63:0] T_636;
  wire [7:0] T_650_0;
  wire [7:0] T_662;
  wire  T_663;
  wire  T_664;
  wire  T_665;
  wire  T_666;
  wire  T_667;
  wire  T_668;
  wire  T_669;
  wire  T_670;
  wire [7:0] GEN_15;
  wire [8:0] T_672;
  wire [7:0] T_673;
  wire [7:0] GEN_16;
  wire [8:0] T_675;
  wire [7:0] T_676;
  wire [7:0] GEN_17;
  wire [8:0] T_678;
  wire [7:0] T_679;
  wire [7:0] GEN_18;
  wire [8:0] T_681;
  wire [7:0] T_682;
  wire [7:0] GEN_19;
  wire [8:0] T_684;
  wire [7:0] T_685;
  wire [7:0] GEN_20;
  wire [8:0] T_687;
  wire [7:0] T_688;
  wire [7:0] GEN_21;
  wire [8:0] T_690;
  wire [7:0] T_691;
  wire [7:0] GEN_22;
  wire [8:0] T_693;
  wire [7:0] T_694;
  wire [7:0] T_700_0;
  wire [7:0] T_700_1;
  wire [7:0] T_700_2;
  wire [7:0] T_700_3;
  wire [7:0] T_700_4;
  wire [7:0] T_700_5;
  wire [7:0] T_700_6;
  wire [7:0] T_700_7;
  wire [15:0] T_702;
  wire [15:0] T_703;
  wire [31:0] T_704;
  wire [15:0] T_705;
  wire [15:0] T_706;
  wire [31:0] T_707;
  wire [63:0] T_708;
  wire [63:0] T_709;
  wire [63:0] GEN_23;
  wire [63:0] T_710;
  wire [63:0] masked_wdata;
  wire  T_727;
  wire [2:0] T_728;
  wire  T_729;
  wire [2:0] T_730;
  wire  T_731;
  wire [2:0] T_732;
  wire  T_733;
  wire [2:0] T_734;
  wire  T_735;
  wire [2:0] T_736;
  wire  T_737;
  wire [2:0] T_738;
  wire  T_739;
  wire [2:0] T_740;
  wire [2:0] T_765_addr_beat;
  wire [1:0] T_765_client_xact_id;
  wire  T_765_manager_xact_id;
  wire  T_765_is_builtin_type;
  wire [3:0] T_765_g_type;
  wire [63:0] T_765_data;
  wire [31:0] T_791;
  wire  T_792;
  wire  GEN_0;
  wire [31:0] GEN_3;
  wire  GEN_4;
  reg  GEN_1;
  reg [31:0] GEN_14;
  Queue_49 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_765_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_765_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_765_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_765_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_765_g_type;
  assign io_tl_grant_bits_data = T_765_data;
  assign io_tiles_0_reset = GEN_1;
  assign io_tiles_0_id = 1'h0;
  assign io_tiles_0_interrupts_mtip = io_interrupts_0_mtip;
  assign io_tiles_0_interrupts_meip = io_interrupts_0_meip;
  assign io_tiles_0_interrupts_seip = io_interrupts_0_seip;
  assign io_tiles_0_interrupts_debug = io_interrupts_0_debug;
  assign io_tiles_0_interrupts_msip = ipi_0;
  assign T_529_0 = 1'h0;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_562 = acq_io_deq_bits_a_type == 3'h2;
  assign write = acq_io_deq_bits_is_builtin_type & T_562;
  assign rdata = GEN_3;
  assign T_565 = acq_io_deq_bits_a_type == 3'h4;
  assign T_566 = acq_io_deq_bits_is_builtin_type & T_565;
  assign GEN_5 = {{7'd0}, 1'h1};
  assign T_570 = 8'h0 - GEN_5;
  assign T_571 = T_570[7:0];
  assign T_577_0 = T_571;
  assign T_580 = acq_io_deq_bits_a_type == 3'h3;
  assign T_581 = acq_io_deq_bits_is_builtin_type & T_580;
  assign T_585 = T_581 | write;
  assign T_586 = acq_io_deq_bits_union[8:1];
  assign T_588 = T_585 ? T_586 : {{7'd0}, 1'h0};
  assign T_589 = T_566 ? T_577_0 : T_588;
  assign T_590 = T_589[0];
  assign T_591 = T_589[1];
  assign T_592 = T_589[2];
  assign T_593 = T_589[3];
  assign T_594 = T_589[4];
  assign T_595 = T_589[5];
  assign T_596 = T_589[6];
  assign T_597 = T_589[7];
  assign GEN_6 = {{7'd0}, T_590};
  assign T_599 = 8'h0 - GEN_6;
  assign T_600 = T_599[7:0];
  assign GEN_7 = {{7'd0}, T_591};
  assign T_602 = 8'h0 - GEN_7;
  assign T_603 = T_602[7:0];
  assign GEN_8 = {{7'd0}, T_592};
  assign T_605 = 8'h0 - GEN_8;
  assign T_606 = T_605[7:0];
  assign GEN_9 = {{7'd0}, T_593};
  assign T_608 = 8'h0 - GEN_9;
  assign T_609 = T_608[7:0];
  assign GEN_10 = {{7'd0}, T_594};
  assign T_611 = 8'h0 - GEN_10;
  assign T_612 = T_611[7:0];
  assign GEN_11 = {{7'd0}, T_595};
  assign T_614 = 8'h0 - GEN_11;
  assign T_615 = T_614[7:0];
  assign GEN_12 = {{7'd0}, T_596};
  assign T_617 = 8'h0 - GEN_12;
  assign T_618 = T_617[7:0];
  assign GEN_13 = {{7'd0}, T_597};
  assign T_620 = 8'h0 - GEN_13;
  assign T_621 = T_620[7:0];
  assign T_627_0 = T_600;
  assign T_627_1 = T_603;
  assign T_627_2 = T_606;
  assign T_627_3 = T_609;
  assign T_627_4 = T_612;
  assign T_627_5 = T_615;
  assign T_627_6 = T_618;
  assign T_627_7 = T_621;
  assign T_629 = {T_627_1,T_627_0};
  assign T_630 = {T_627_3,T_627_2};
  assign T_631 = {T_630,T_629};
  assign T_632 = {T_627_5,T_627_4};
  assign T_633 = {T_627_7,T_627_6};
  assign T_634 = {T_633,T_632};
  assign T_635 = {T_634,T_631};
  assign T_636 = acq_io_deq_bits_data & T_635;
  assign T_650_0 = T_571;
  assign T_662 = T_566 ? T_650_0 : T_588;
  assign T_663 = T_662[0];
  assign T_664 = T_662[1];
  assign T_665 = T_662[2];
  assign T_666 = T_662[3];
  assign T_667 = T_662[4];
  assign T_668 = T_662[5];
  assign T_669 = T_662[6];
  assign T_670 = T_662[7];
  assign GEN_15 = {{7'd0}, T_663};
  assign T_672 = 8'h0 - GEN_15;
  assign T_673 = T_672[7:0];
  assign GEN_16 = {{7'd0}, T_664};
  assign T_675 = 8'h0 - GEN_16;
  assign T_676 = T_675[7:0];
  assign GEN_17 = {{7'd0}, T_665};
  assign T_678 = 8'h0 - GEN_17;
  assign T_679 = T_678[7:0];
  assign GEN_18 = {{7'd0}, T_666};
  assign T_681 = 8'h0 - GEN_18;
  assign T_682 = T_681[7:0];
  assign GEN_19 = {{7'd0}, T_667};
  assign T_684 = 8'h0 - GEN_19;
  assign T_685 = T_684[7:0];
  assign GEN_20 = {{7'd0}, T_668};
  assign T_687 = 8'h0 - GEN_20;
  assign T_688 = T_687[7:0];
  assign GEN_21 = {{7'd0}, T_669};
  assign T_690 = 8'h0 - GEN_21;
  assign T_691 = T_690[7:0];
  assign GEN_22 = {{7'd0}, T_670};
  assign T_693 = 8'h0 - GEN_22;
  assign T_694 = T_693[7:0];
  assign T_700_0 = T_673;
  assign T_700_1 = T_676;
  assign T_700_2 = T_679;
  assign T_700_3 = T_682;
  assign T_700_4 = T_685;
  assign T_700_5 = T_688;
  assign T_700_6 = T_691;
  assign T_700_7 = T_694;
  assign T_702 = {T_700_1,T_700_0};
  assign T_703 = {T_700_3,T_700_2};
  assign T_704 = {T_703,T_702};
  assign T_705 = {T_700_5,T_700_4};
  assign T_706 = {T_700_7,T_700_6};
  assign T_707 = {T_706,T_705};
  assign T_708 = {T_707,T_704};
  assign T_709 = ~ T_708;
  assign GEN_23 = {{32'd0}, rdata};
  assign T_710 = GEN_23 & T_709;
  assign masked_wdata = T_636 | T_710;
  assign T_727 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_728 = T_727 ? 3'h1 : 3'h3;
  assign T_729 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_730 = T_729 ? 3'h1 : T_728;
  assign T_731 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_732 = T_731 ? 3'h4 : T_730;
  assign T_733 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_734 = T_733 ? 3'h3 : T_732;
  assign T_735 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_736 = T_735 ? 3'h3 : T_734;
  assign T_737 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_738 = T_737 ? 3'h5 : T_736;
  assign T_739 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_740 = T_739 ? 3'h4 : T_738;
  assign T_765_addr_beat = {{2'd0}, 1'h0};
  assign T_765_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_765_manager_xact_id = 1'h0;
  assign T_765_is_builtin_type = 1'h1;
  assign T_765_g_type = {{1'd0}, T_740};
  assign T_765_data = {{32'd0}, rdata};
  assign T_791 = {31'h0,ipi_0};
  assign T_792 = masked_wdata[0];
  assign GEN_0 = write ? T_792 : ipi_0;
  assign GEN_3 = write ? T_791 : {{31'd0}, 1'h0};
  assign GEN_4 = write ? GEN_0 : ipi_0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_2 = {1{$random}};
  ipi_0 = GEN_2[0:0];
  GEN_14 = {1{$random}};
  GEN_1 = GEN_14[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      ipi_0 <= T_529_0;
    end else begin
      ipi_0 <= GEN_4;
    end
  end
endmodule
module ROMSlave(
  input   clk,
  input   reset,
  output  io_acquire_ready,
  input   io_acquire_valid,
  input  [25:0] io_acquire_bits_addr_block,
  input  [1:0] io_acquire_bits_client_xact_id,
  input  [2:0] io_acquire_bits_addr_beat,
  input   io_acquire_bits_is_builtin_type,
  input  [2:0] io_acquire_bits_a_type,
  input  [11:0] io_acquire_bits_union,
  input  [63:0] io_acquire_bits_data,
  input   io_grant_ready,
  output  io_grant_valid,
  output [2:0] io_grant_bits_addr_beat,
  output [1:0] io_grant_bits_client_xact_id,
  output  io_grant_bits_manager_xact_id,
  output  io_grant_bits_is_builtin_type,
  output [3:0] io_grant_bits_g_type,
  output [63:0] io_grant_bits_data
);
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_446;
  wire  single_beat;
  wire  T_448;
  wire  multi_beat;
  wire  T_450;
  wire  T_451;
  wire  T_452;
  wire  T_453;
  wire  T_455;
  reg [2:0] addr_beat;
  reg [31:0] GEN_136;
  wire  T_457;
  wire [2:0] GEN_72;
  wire [3:0] T_459;
  wire [2:0] T_460;
  wire [2:0] GEN_1;
  wire  T_461;
  wire [2:0] GEN_2;
  wire [63:0] rom_0;
  wire [63:0] rom_1;
  wire [63:0] rom_2;
  wire [63:0] rom_3;
  wire [63:0] rom_4;
  wire [63:0] rom_5;
  wire [63:0] rom_6;
  wire [63:0] rom_7;
  wire [63:0] rom_8;
  wire [63:0] rom_9;
  wire [63:0] rom_10;
  wire [63:0] rom_11;
  wire [63:0] rom_12;
  wire [63:0] rom_13;
  wire [63:0] rom_14;
  wire [63:0] rom_15;
  wire [63:0] rom_16;
  wire [63:0] rom_17;
  wire [63:0] rom_18;
  wire [63:0] rom_19;
  wire [63:0] rom_20;
  wire [63:0] rom_21;
  wire [63:0] rom_22;
  wire [63:0] rom_23;
  wire [63:0] rom_24;
  wire [63:0] rom_25;
  wire [63:0] rom_26;
  wire [63:0] rom_27;
  wire [63:0] rom_28;
  wire [63:0] rom_29;
  wire [63:0] rom_30;
  wire [63:0] rom_31;
  wire [63:0] rom_32;
  wire [63:0] rom_33;
  wire [63:0] rom_34;
  wire [63:0] rom_35;
  wire [63:0] rom_36;
  wire [63:0] rom_37;
  wire [63:0] rom_38;
  wire [63:0] rom_39;
  wire [63:0] rom_40;
  wire [63:0] rom_41;
  wire [63:0] rom_42;
  wire [63:0] rom_43;
  wire [63:0] rom_44;
  wire [63:0] rom_45;
  wire [63:0] rom_46;
  wire [63:0] rom_47;
  wire [63:0] rom_48;
  wire [63:0] rom_49;
  wire [63:0] rom_50;
  wire [63:0] rom_51;
  wire [63:0] rom_52;
  wire [63:0] rom_53;
  wire [63:0] rom_54;
  wire [63:0] rom_55;
  wire [63:0] rom_56;
  wire [63:0] rom_57;
  wire [63:0] rom_58;
  wire [63:0] rom_59;
  wire [63:0] rom_60;
  wire [63:0] rom_61;
  wire [63:0] rom_62;
  wire [63:0] rom_63;
  wire [63:0] rom_64;
  wire [63:0] rom_65;
  wire [63:0] rom_66;
  wire [63:0] rom_67;
  wire [63:0] rom_68;
  wire [63:0] rom_69;
  wire [28:0] raddr;
  wire [6:0] T_538;
  wire  T_540;
  wire  T_542;
  wire  last;
  wire  T_543;
  wire  T_560;
  wire [2:0] T_561;
  wire  T_562;
  wire [2:0] T_563;
  wire  T_564;
  wire [2:0] T_565;
  wire  T_566;
  wire [2:0] T_567;
  wire  T_568;
  wire [2:0] T_569;
  wire  T_570;
  wire [2:0] T_571;
  wire  T_572;
  wire [2:0] T_573;
  wire [2:0] T_597_addr_beat;
  wire [1:0] T_597_client_xact_id;
  wire  T_597_manager_xact_id;
  wire  T_597_is_builtin_type;
  wire [3:0] T_597_g_type;
  wire [63:0] T_597_data;
  wire [63:0] GEN_0;
  wire [6:0] GEN_73;
  wire [63:0] GEN_3;
  wire [6:0] GEN_74;
  wire [63:0] GEN_4;
  wire [6:0] GEN_75;
  wire [63:0] GEN_5;
  wire [6:0] GEN_76;
  wire [63:0] GEN_6;
  wire [6:0] GEN_77;
  wire [63:0] GEN_7;
  wire [6:0] GEN_78;
  wire [63:0] GEN_8;
  wire [6:0] GEN_79;
  wire [63:0] GEN_9;
  wire [6:0] GEN_80;
  wire [63:0] GEN_10;
  wire [6:0] GEN_81;
  wire [63:0] GEN_11;
  wire [6:0] GEN_82;
  wire [63:0] GEN_12;
  wire [6:0] GEN_83;
  wire [63:0] GEN_13;
  wire [6:0] GEN_84;
  wire [63:0] GEN_14;
  wire [6:0] GEN_85;
  wire [63:0] GEN_15;
  wire [6:0] GEN_86;
  wire [63:0] GEN_16;
  wire [6:0] GEN_87;
  wire [63:0] GEN_17;
  wire [6:0] GEN_88;
  wire [63:0] GEN_18;
  wire [6:0] GEN_89;
  wire [63:0] GEN_19;
  wire [6:0] GEN_90;
  wire [63:0] GEN_20;
  wire [6:0] GEN_91;
  wire [63:0] GEN_21;
  wire [6:0] GEN_92;
  wire [63:0] GEN_22;
  wire [6:0] GEN_93;
  wire [63:0] GEN_23;
  wire [6:0] GEN_94;
  wire [63:0] GEN_24;
  wire [6:0] GEN_95;
  wire [63:0] GEN_25;
  wire [6:0] GEN_96;
  wire [63:0] GEN_26;
  wire [6:0] GEN_97;
  wire [63:0] GEN_27;
  wire [6:0] GEN_98;
  wire [63:0] GEN_28;
  wire [6:0] GEN_99;
  wire [63:0] GEN_29;
  wire [6:0] GEN_100;
  wire [63:0] GEN_30;
  wire [6:0] GEN_101;
  wire [63:0] GEN_31;
  wire [6:0] GEN_102;
  wire [63:0] GEN_32;
  wire [6:0] GEN_103;
  wire [63:0] GEN_33;
  wire [6:0] GEN_104;
  wire [63:0] GEN_34;
  wire [6:0] GEN_105;
  wire [63:0] GEN_35;
  wire [6:0] GEN_106;
  wire [63:0] GEN_36;
  wire [6:0] GEN_107;
  wire [63:0] GEN_37;
  wire [6:0] GEN_108;
  wire [63:0] GEN_38;
  wire [6:0] GEN_109;
  wire [63:0] GEN_39;
  wire [6:0] GEN_110;
  wire [63:0] GEN_40;
  wire [6:0] GEN_111;
  wire [63:0] GEN_41;
  wire [6:0] GEN_112;
  wire [63:0] GEN_42;
  wire [6:0] GEN_113;
  wire [63:0] GEN_43;
  wire [6:0] GEN_114;
  wire [63:0] GEN_44;
  wire [6:0] GEN_115;
  wire [63:0] GEN_45;
  wire [6:0] GEN_116;
  wire [63:0] GEN_46;
  wire [6:0] GEN_117;
  wire [63:0] GEN_47;
  wire [6:0] GEN_118;
  wire [63:0] GEN_48;
  wire [6:0] GEN_119;
  wire [63:0] GEN_49;
  wire [6:0] GEN_120;
  wire [63:0] GEN_50;
  wire [6:0] GEN_121;
  wire [63:0] GEN_51;
  wire [6:0] GEN_122;
  wire [63:0] GEN_52;
  wire [6:0] GEN_123;
  wire [63:0] GEN_53;
  wire [6:0] GEN_124;
  wire [63:0] GEN_54;
  wire [6:0] GEN_125;
  wire [63:0] GEN_55;
  wire [6:0] GEN_126;
  wire [63:0] GEN_56;
  wire [6:0] GEN_127;
  wire [63:0] GEN_57;
  wire [6:0] GEN_128;
  wire [63:0] GEN_58;
  wire [6:0] GEN_129;
  wire [63:0] GEN_59;
  wire [6:0] GEN_130;
  wire [63:0] GEN_60;
  wire [6:0] GEN_131;
  wire [63:0] GEN_61;
  wire [6:0] GEN_132;
  wire [63:0] GEN_62;
  wire [6:0] GEN_133;
  wire [63:0] GEN_63;
  wire [6:0] GEN_134;
  wire [63:0] GEN_64;
  wire [6:0] GEN_135;
  wire [63:0] GEN_65;
  wire [63:0] GEN_66;
  wire [63:0] GEN_67;
  wire [63:0] GEN_68;
  wire [63:0] GEN_69;
  wire [63:0] GEN_70;
  wire [63:0] GEN_71;
  Queue_49 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_acquire_ready = acq_io_enq_ready;
  assign io_grant_valid = acq_io_deq_valid;
  assign io_grant_bits_addr_beat = T_597_addr_beat;
  assign io_grant_bits_client_xact_id = T_597_client_xact_id;
  assign io_grant_bits_manager_xact_id = T_597_manager_xact_id;
  assign io_grant_bits_is_builtin_type = T_597_is_builtin_type;
  assign io_grant_bits_g_type = T_597_g_type;
  assign io_grant_bits_data = T_597_data;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_acquire_bits_union;
  assign acq_io_enq_bits_data = io_acquire_bits_data;
  assign acq_io_deq_ready = T_543;
  assign T_446 = acq_io_deq_bits_a_type == 3'h0;
  assign single_beat = acq_io_deq_bits_is_builtin_type & T_446;
  assign T_448 = acq_io_deq_bits_a_type == 3'h1;
  assign multi_beat = acq_io_deq_bits_is_builtin_type & T_448;
  assign T_450 = acq_io_deq_valid == 1'h0;
  assign T_451 = T_450 | single_beat;
  assign T_452 = T_451 | multi_beat;
  assign T_453 = T_452 | reset;
  assign T_455 = T_453 == 1'h0;
  assign T_457 = io_grant_ready & io_grant_valid;
  assign GEN_72 = {{2'd0}, 1'h1};
  assign T_459 = addr_beat + GEN_72;
  assign T_460 = T_459[2:0];
  assign GEN_1 = T_457 ? T_460 : addr_beat;
  assign T_461 = io_acquire_ready & io_acquire_valid;
  assign GEN_2 = T_461 ? io_acquire_bits_addr_beat : GEN_1;
  assign rom_0 = 64'h280677ffff297;
  assign rom_1 = 64'h102000000000;
  assign rom_2 = 64'h0;
  assign rom_3 = 64'h0;
  assign rom_4 = 64'h6d726f6674616c70;
  assign rom_5 = 64'h6e657620200a7b20;
  assign rom_6 = 64'h3b62637520726f64;
  assign rom_7 = 64'h206863726120200a;
  assign rom_8 = 64'ha3b74656b636f72;
  assign rom_9 = 64'h2063696c700a3b7d;
  assign rom_10 = 64'h6f69727020200a7b;
  assign rom_11 = 64'h3478302079746972;
  assign rom_12 = 64'h3b30303030303030;
  assign rom_13 = 64'h69646e657020200a;
  assign rom_14 = 64'h303034783020676e;
  assign rom_15 = 64'h200a3b3030303130;
  assign rom_16 = 64'h3220737665646e20;
  assign rom_17 = 64'h6374720a3b7d0a3b;
  assign rom_18 = 64'h64646120200a7b20;
  assign rom_19 = 64'h3030303278302072;
  assign rom_20 = 64'h6d61720a3b7d0a3b;
  assign rom_21 = 64'h7b203020200a7b20;
  assign rom_22 = 64'h646461202020200a;
  assign rom_23 = 64'h3030303878302072;
  assign rom_24 = 64'h20200a3b30303030;
  assign rom_25 = 64'h3020657a69732020;
  assign rom_26 = 64'h3030303030303878;
  assign rom_27 = 64'ha3b7d20200a3b30;
  assign rom_28 = 64'h2065726f630a3b7d;
  assign rom_29 = 64'ha7b203020200a7b;
  assign rom_30 = 64'ha7b203020202020;
  assign rom_31 = 64'h7369202020202020;
  assign rom_32 = 64'h6d69343676722061;
  assign rom_33 = 64'h2020200a3b646661;
  assign rom_34 = 64'h63656d6974202020;
  assign rom_35 = 64'h303032783020706d;
  assign rom_36 = 64'h20202020200a3b38;
  assign rom_37 = 64'h3478302069706920;
  assign rom_38 = 64'h3b30303030303034;
  assign rom_39 = 64'h702020202020200a;
  assign rom_40 = 64'h20200a7b2063696c;
  assign rom_41 = 64'h206d202020202020;
  assign rom_42 = 64'h2020202020200a7b;
  assign rom_43 = 64'h7830206569202020;
  assign rom_44 = 64'h3030303230303034;
  assign rom_45 = 64'h2020202020200a3b;
  assign rom_46 = 64'h7365726874202020;
  assign rom_47 = 64'h3032303478302068;
  assign rom_48 = 64'h20200a3b30303030;
  assign rom_49 = 64'h6320202020202020;
  assign rom_50 = 64'h347830206d69616c;
  assign rom_51 = 64'h3b34303030303230;
  assign rom_52 = 64'h202020202020200a;
  assign rom_53 = 64'h202020200a3b7d20;
  assign rom_54 = 64'ha7b207320202020;
  assign rom_55 = 64'h2020202020202020;
  assign rom_56 = 64'h3034783020656920;
  assign rom_57 = 64'ha3b303830323030;
  assign rom_58 = 64'h2020202020202020;
  assign rom_59 = 64'h2068736572687420;
  assign rom_60 = 64'h3031303230347830;
  assign rom_61 = 64'h202020200a3b3030;
  assign rom_62 = 64'h616c632020202020;
  assign rom_63 = 64'h3230347830206d69;
  assign rom_64 = 64'h200a3b3430303130;
  assign rom_65 = 64'h7d20202020202020;
  assign rom_66 = 64'h2020202020200a3b;
  assign rom_67 = 64'h7d202020200a3b7d;
  assign rom_68 = 64'h7d0a3b7d20200a3b;
  assign rom_69 = 64'ha3b;
  assign raddr = {acq_io_deq_bits_addr_block,addr_beat};
  assign T_538 = raddr[6:0];
  assign T_540 = multi_beat == 1'h0;
  assign T_542 = addr_beat == 3'h7;
  assign last = T_540 | T_542;
  assign T_543 = io_grant_ready & last;
  assign T_560 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_561 = T_560 ? 3'h1 : 3'h3;
  assign T_562 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_563 = T_562 ? 3'h1 : T_561;
  assign T_564 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_565 = T_564 ? 3'h4 : T_563;
  assign T_566 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_567 = T_566 ? 3'h3 : T_565;
  assign T_568 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_569 = T_568 ? 3'h3 : T_567;
  assign T_570 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_571 = T_570 ? 3'h5 : T_569;
  assign T_572 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_573 = T_572 ? 3'h4 : T_571;
  assign T_597_addr_beat = addr_beat;
  assign T_597_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_597_manager_xact_id = 1'h0;
  assign T_597_is_builtin_type = 1'h1;
  assign T_597_g_type = {{1'd0}, T_573};
  assign T_597_data = GEN_0;
  assign GEN_0 = GEN_71;
  assign GEN_73 = {{6'd0}, 1'h1};
  assign GEN_3 = GEN_73 == T_538 ? rom_1 : rom_0;
  assign GEN_74 = {{5'd0}, 2'h2};
  assign GEN_4 = GEN_74 == T_538 ? rom_2 : GEN_3;
  assign GEN_75 = {{5'd0}, 2'h3};
  assign GEN_5 = GEN_75 == T_538 ? rom_3 : GEN_4;
  assign GEN_76 = {{4'd0}, 3'h4};
  assign GEN_6 = GEN_76 == T_538 ? rom_4 : GEN_5;
  assign GEN_77 = {{4'd0}, 3'h5};
  assign GEN_7 = GEN_77 == T_538 ? rom_5 : GEN_6;
  assign GEN_78 = {{4'd0}, 3'h6};
  assign GEN_8 = GEN_78 == T_538 ? rom_6 : GEN_7;
  assign GEN_79 = {{4'd0}, 3'h7};
  assign GEN_9 = GEN_79 == T_538 ? rom_7 : GEN_8;
  assign GEN_80 = {{3'd0}, 4'h8};
  assign GEN_10 = GEN_80 == T_538 ? rom_8 : GEN_9;
  assign GEN_81 = {{3'd0}, 4'h9};
  assign GEN_11 = GEN_81 == T_538 ? rom_9 : GEN_10;
  assign GEN_82 = {{3'd0}, 4'ha};
  assign GEN_12 = GEN_82 == T_538 ? rom_10 : GEN_11;
  assign GEN_83 = {{3'd0}, 4'hb};
  assign GEN_13 = GEN_83 == T_538 ? rom_11 : GEN_12;
  assign GEN_84 = {{3'd0}, 4'hc};
  assign GEN_14 = GEN_84 == T_538 ? rom_12 : GEN_13;
  assign GEN_85 = {{3'd0}, 4'hd};
  assign GEN_15 = GEN_85 == T_538 ? rom_13 : GEN_14;
  assign GEN_86 = {{3'd0}, 4'he};
  assign GEN_16 = GEN_86 == T_538 ? rom_14 : GEN_15;
  assign GEN_87 = {{3'd0}, 4'hf};
  assign GEN_17 = GEN_87 == T_538 ? rom_15 : GEN_16;
  assign GEN_88 = {{2'd0}, 5'h10};
  assign GEN_18 = GEN_88 == T_538 ? rom_16 : GEN_17;
  assign GEN_89 = {{2'd0}, 5'h11};
  assign GEN_19 = GEN_89 == T_538 ? rom_17 : GEN_18;
  assign GEN_90 = {{2'd0}, 5'h12};
  assign GEN_20 = GEN_90 == T_538 ? rom_18 : GEN_19;
  assign GEN_91 = {{2'd0}, 5'h13};
  assign GEN_21 = GEN_91 == T_538 ? rom_19 : GEN_20;
  assign GEN_92 = {{2'd0}, 5'h14};
  assign GEN_22 = GEN_92 == T_538 ? rom_20 : GEN_21;
  assign GEN_93 = {{2'd0}, 5'h15};
  assign GEN_23 = GEN_93 == T_538 ? rom_21 : GEN_22;
  assign GEN_94 = {{2'd0}, 5'h16};
  assign GEN_24 = GEN_94 == T_538 ? rom_22 : GEN_23;
  assign GEN_95 = {{2'd0}, 5'h17};
  assign GEN_25 = GEN_95 == T_538 ? rom_23 : GEN_24;
  assign GEN_96 = {{2'd0}, 5'h18};
  assign GEN_26 = GEN_96 == T_538 ? rom_24 : GEN_25;
  assign GEN_97 = {{2'd0}, 5'h19};
  assign GEN_27 = GEN_97 == T_538 ? rom_25 : GEN_26;
  assign GEN_98 = {{2'd0}, 5'h1a};
  assign GEN_28 = GEN_98 == T_538 ? rom_26 : GEN_27;
  assign GEN_99 = {{2'd0}, 5'h1b};
  assign GEN_29 = GEN_99 == T_538 ? rom_27 : GEN_28;
  assign GEN_100 = {{2'd0}, 5'h1c};
  assign GEN_30 = GEN_100 == T_538 ? rom_28 : GEN_29;
  assign GEN_101 = {{2'd0}, 5'h1d};
  assign GEN_31 = GEN_101 == T_538 ? rom_29 : GEN_30;
  assign GEN_102 = {{2'd0}, 5'h1e};
  assign GEN_32 = GEN_102 == T_538 ? rom_30 : GEN_31;
  assign GEN_103 = {{2'd0}, 5'h1f};
  assign GEN_33 = GEN_103 == T_538 ? rom_31 : GEN_32;
  assign GEN_104 = {{1'd0}, 6'h20};
  assign GEN_34 = GEN_104 == T_538 ? rom_32 : GEN_33;
  assign GEN_105 = {{1'd0}, 6'h21};
  assign GEN_35 = GEN_105 == T_538 ? rom_33 : GEN_34;
  assign GEN_106 = {{1'd0}, 6'h22};
  assign GEN_36 = GEN_106 == T_538 ? rom_34 : GEN_35;
  assign GEN_107 = {{1'd0}, 6'h23};
  assign GEN_37 = GEN_107 == T_538 ? rom_35 : GEN_36;
  assign GEN_108 = {{1'd0}, 6'h24};
  assign GEN_38 = GEN_108 == T_538 ? rom_36 : GEN_37;
  assign GEN_109 = {{1'd0}, 6'h25};
  assign GEN_39 = GEN_109 == T_538 ? rom_37 : GEN_38;
  assign GEN_110 = {{1'd0}, 6'h26};
  assign GEN_40 = GEN_110 == T_538 ? rom_38 : GEN_39;
  assign GEN_111 = {{1'd0}, 6'h27};
  assign GEN_41 = GEN_111 == T_538 ? rom_39 : GEN_40;
  assign GEN_112 = {{1'd0}, 6'h28};
  assign GEN_42 = GEN_112 == T_538 ? rom_40 : GEN_41;
  assign GEN_113 = {{1'd0}, 6'h29};
  assign GEN_43 = GEN_113 == T_538 ? rom_41 : GEN_42;
  assign GEN_114 = {{1'd0}, 6'h2a};
  assign GEN_44 = GEN_114 == T_538 ? rom_42 : GEN_43;
  assign GEN_115 = {{1'd0}, 6'h2b};
  assign GEN_45 = GEN_115 == T_538 ? rom_43 : GEN_44;
  assign GEN_116 = {{1'd0}, 6'h2c};
  assign GEN_46 = GEN_116 == T_538 ? rom_44 : GEN_45;
  assign GEN_117 = {{1'd0}, 6'h2d};
  assign GEN_47 = GEN_117 == T_538 ? rom_45 : GEN_46;
  assign GEN_118 = {{1'd0}, 6'h2e};
  assign GEN_48 = GEN_118 == T_538 ? rom_46 : GEN_47;
  assign GEN_119 = {{1'd0}, 6'h2f};
  assign GEN_49 = GEN_119 == T_538 ? rom_47 : GEN_48;
  assign GEN_120 = {{1'd0}, 6'h30};
  assign GEN_50 = GEN_120 == T_538 ? rom_48 : GEN_49;
  assign GEN_121 = {{1'd0}, 6'h31};
  assign GEN_51 = GEN_121 == T_538 ? rom_49 : GEN_50;
  assign GEN_122 = {{1'd0}, 6'h32};
  assign GEN_52 = GEN_122 == T_538 ? rom_50 : GEN_51;
  assign GEN_123 = {{1'd0}, 6'h33};
  assign GEN_53 = GEN_123 == T_538 ? rom_51 : GEN_52;
  assign GEN_124 = {{1'd0}, 6'h34};
  assign GEN_54 = GEN_124 == T_538 ? rom_52 : GEN_53;
  assign GEN_125 = {{1'd0}, 6'h35};
  assign GEN_55 = GEN_125 == T_538 ? rom_53 : GEN_54;
  assign GEN_126 = {{1'd0}, 6'h36};
  assign GEN_56 = GEN_126 == T_538 ? rom_54 : GEN_55;
  assign GEN_127 = {{1'd0}, 6'h37};
  assign GEN_57 = GEN_127 == T_538 ? rom_55 : GEN_56;
  assign GEN_128 = {{1'd0}, 6'h38};
  assign GEN_58 = GEN_128 == T_538 ? rom_56 : GEN_57;
  assign GEN_129 = {{1'd0}, 6'h39};
  assign GEN_59 = GEN_129 == T_538 ? rom_57 : GEN_58;
  assign GEN_130 = {{1'd0}, 6'h3a};
  assign GEN_60 = GEN_130 == T_538 ? rom_58 : GEN_59;
  assign GEN_131 = {{1'd0}, 6'h3b};
  assign GEN_61 = GEN_131 == T_538 ? rom_59 : GEN_60;
  assign GEN_132 = {{1'd0}, 6'h3c};
  assign GEN_62 = GEN_132 == T_538 ? rom_60 : GEN_61;
  assign GEN_133 = {{1'd0}, 6'h3d};
  assign GEN_63 = GEN_133 == T_538 ? rom_61 : GEN_62;
  assign GEN_134 = {{1'd0}, 6'h3e};
  assign GEN_64 = GEN_134 == T_538 ? rom_62 : GEN_63;
  assign GEN_135 = {{1'd0}, 6'h3f};
  assign GEN_65 = GEN_135 == T_538 ? rom_63 : GEN_64;
  assign GEN_66 = 7'h40 == T_538 ? rom_64 : GEN_65;
  assign GEN_67 = 7'h41 == T_538 ? rom_65 : GEN_66;
  assign GEN_68 = 7'h42 == T_538 ? rom_66 : GEN_67;
  assign GEN_69 = 7'h43 == T_538 ? rom_67 : GEN_68;
  assign GEN_70 = 7'h44 == T_538 ? rom_68 : GEN_69;
  assign GEN_71 = 7'h45 == T_538 ? rom_69 : GEN_70;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_136 = {1{$random}};
  addr_beat = GEN_136[2:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      addr_beat <= GEN_2;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported ROMSlave operation\n    at rom.scala:15 assert(!acq.valid || single_beat || multi_beat, \"unsupported ROMSlave operation\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_455) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_55(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [4:0] io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output [4:0] io_deq_bits,
  output  io_count
);
  reg [4:0] ram [0:0];
  reg [31:0] GEN_0;
  wire [4:0] ram_T_34_data;
  wire  ram_T_34_addr;
  wire  ram_T_34_en;
  wire [4:0] ram_T_26_data;
  wire  ram_T_26_addr;
  wire  ram_T_26_mask;
  wire  ram_T_26_en;
  reg  maybe_full;
  reg [31:0] GEN_1;
  wire  T_23;
  wire  T_24;
  wire  do_enq;
  wire  T_25;
  wire  do_deq;
  wire  T_29;
  wire  GEN_5;
  wire  T_31;
  wire [1:0] T_35;
  wire  ptr_diff;
  wire [1:0] T_37;
  assign io_enq_ready = T_23;
  assign io_deq_valid = T_31;
  assign io_deq_bits = ram_T_34_data;
  assign io_count = T_37[0];
  assign ram_T_34_addr = 1'h0;
  assign ram_T_34_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_T_34_data = ram[ram_T_34_addr];
  `else
  assign ram_T_34_data = ram_T_34_addr >= 1'h1 ? $random : ram[ram_T_34_addr];
  `endif
  assign ram_T_26_data = io_enq_bits;
  assign ram_T_26_addr = 1'h0;
  assign ram_T_26_mask = do_enq;
  assign ram_T_26_en = do_enq;
  assign T_23 = maybe_full == 1'h0;
  assign T_24 = io_enq_ready & io_enq_valid;
  assign do_enq = T_24;
  assign T_25 = io_deq_ready & io_deq_valid;
  assign do_deq = T_25;
  assign T_29 = do_enq != do_deq;
  assign GEN_5 = T_29 ? do_enq : maybe_full;
  assign T_31 = T_23 == 1'h0;
  assign T_35 = 1'h0 - 1'h0;
  assign ptr_diff = T_35[0:0];
  assign T_37 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = GEN_0[4:0];
  GEN_1 = {1{$random}};
  maybe_full = GEN_1[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_T_26_en & ram_T_26_mask) begin
      ram[ram_T_26_addr] <= ram_T_26_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_5;
    end
  end
endmodule
module NastiErrorSlave(
  input   clk,
  input   reset,
  output  io_aw_ready,
  input   io_aw_valid,
  input  [31:0] io_aw_bits_addr,
  input  [7:0] io_aw_bits_len,
  input  [2:0] io_aw_bits_size,
  input  [1:0] io_aw_bits_burst,
  input   io_aw_bits_lock,
  input  [3:0] io_aw_bits_cache,
  input  [2:0] io_aw_bits_prot,
  input  [3:0] io_aw_bits_qos,
  input  [3:0] io_aw_bits_region,
  input  [4:0] io_aw_bits_id,
  input   io_aw_bits_user,
  output  io_w_ready,
  input   io_w_valid,
  input  [63:0] io_w_bits_data,
  input   io_w_bits_last,
  input  [4:0] io_w_bits_id,
  input  [7:0] io_w_bits_strb,
  input   io_w_bits_user,
  input   io_b_ready,
  output  io_b_valid,
  output [1:0] io_b_bits_resp,
  output [4:0] io_b_bits_id,
  output  io_b_bits_user,
  output  io_ar_ready,
  input   io_ar_valid,
  input  [31:0] io_ar_bits_addr,
  input  [7:0] io_ar_bits_len,
  input  [2:0] io_ar_bits_size,
  input  [1:0] io_ar_bits_burst,
  input   io_ar_bits_lock,
  input  [3:0] io_ar_bits_cache,
  input  [2:0] io_ar_bits_prot,
  input  [3:0] io_ar_bits_qos,
  input  [3:0] io_ar_bits_region,
  input  [4:0] io_ar_bits_id,
  input   io_ar_bits_user,
  input   io_r_ready,
  output  io_r_valid,
  output [1:0] io_r_bits_resp,
  output [63:0] io_r_bits_data,
  output  io_r_bits_last,
  output [4:0] io_r_bits_id,
  output  io_r_bits_user
);
  wire  T_323;
  wire  T_325;
  wire  T_326;
  wire  r_queue_clk;
  wire  r_queue_reset;
  wire  r_queue_io_enq_ready;
  wire  r_queue_io_enq_valid;
  wire [31:0] r_queue_io_enq_bits_addr;
  wire [7:0] r_queue_io_enq_bits_len;
  wire [2:0] r_queue_io_enq_bits_size;
  wire [1:0] r_queue_io_enq_bits_burst;
  wire  r_queue_io_enq_bits_lock;
  wire [3:0] r_queue_io_enq_bits_cache;
  wire [2:0] r_queue_io_enq_bits_prot;
  wire [3:0] r_queue_io_enq_bits_qos;
  wire [3:0] r_queue_io_enq_bits_region;
  wire [4:0] r_queue_io_enq_bits_id;
  wire  r_queue_io_enq_bits_user;
  wire  r_queue_io_deq_ready;
  wire  r_queue_io_deq_valid;
  wire [31:0] r_queue_io_deq_bits_addr;
  wire [7:0] r_queue_io_deq_bits_len;
  wire [2:0] r_queue_io_deq_bits_size;
  wire [1:0] r_queue_io_deq_bits_burst;
  wire  r_queue_io_deq_bits_lock;
  wire [3:0] r_queue_io_deq_bits_cache;
  wire [2:0] r_queue_io_deq_bits_prot;
  wire [3:0] r_queue_io_deq_bits_qos;
  wire [3:0] r_queue_io_deq_bits_region;
  wire [4:0] r_queue_io_deq_bits_id;
  wire  r_queue_io_deq_bits_user;
  wire  r_queue_io_count;
  reg  responding;
  reg [31:0] GEN_12;
  reg [7:0] beats_left;
  reg [31:0] GEN_13;
  wire  T_344;
  wire  T_345;
  wire  GEN_0;
  wire [7:0] GEN_1;
  wire  T_347;
  wire [7:0] GEN_8;
  wire  T_350;
  wire  T_351;
  wire  T_352;
  wire  GEN_2;
  wire  T_358;
  wire [7:0] GEN_10;
  wire [8:0] T_360;
  wire [7:0] T_361;
  wire [7:0] GEN_3;
  wire  GEN_4;
  wire [7:0] GEN_5;
  reg  draining;
  reg [31:0] GEN_14;
  wire  GEN_6;
  wire  T_365;
  wire  T_366;
  wire  GEN_7;
  wire  b_queue_clk;
  wire  b_queue_reset;
  wire  b_queue_io_enq_ready;
  wire  b_queue_io_enq_valid;
  wire [4:0] b_queue_io_enq_bits;
  wire  b_queue_io_deq_ready;
  wire  b_queue_io_deq_valid;
  wire [4:0] b_queue_io_deq_bits;
  wire  b_queue_io_count;
  wire  T_370;
  wire  T_371;
  wire  T_374;
  wire  T_377;
  wire  T_381;
  reg  GEN_9;
  reg [31:0] GEN_15;
  reg  GEN_11;
  reg [31:0] GEN_16;
  Queue_39 r_queue (
    .clk(r_queue_clk),
    .reset(r_queue_reset),
    .io_enq_ready(r_queue_io_enq_ready),
    .io_enq_valid(r_queue_io_enq_valid),
    .io_enq_bits_addr(r_queue_io_enq_bits_addr),
    .io_enq_bits_len(r_queue_io_enq_bits_len),
    .io_enq_bits_size(r_queue_io_enq_bits_size),
    .io_enq_bits_burst(r_queue_io_enq_bits_burst),
    .io_enq_bits_lock(r_queue_io_enq_bits_lock),
    .io_enq_bits_cache(r_queue_io_enq_bits_cache),
    .io_enq_bits_prot(r_queue_io_enq_bits_prot),
    .io_enq_bits_qos(r_queue_io_enq_bits_qos),
    .io_enq_bits_region(r_queue_io_enq_bits_region),
    .io_enq_bits_id(r_queue_io_enq_bits_id),
    .io_enq_bits_user(r_queue_io_enq_bits_user),
    .io_deq_ready(r_queue_io_deq_ready),
    .io_deq_valid(r_queue_io_deq_valid),
    .io_deq_bits_addr(r_queue_io_deq_bits_addr),
    .io_deq_bits_len(r_queue_io_deq_bits_len),
    .io_deq_bits_size(r_queue_io_deq_bits_size),
    .io_deq_bits_burst(r_queue_io_deq_bits_burst),
    .io_deq_bits_lock(r_queue_io_deq_bits_lock),
    .io_deq_bits_cache(r_queue_io_deq_bits_cache),
    .io_deq_bits_prot(r_queue_io_deq_bits_prot),
    .io_deq_bits_qos(r_queue_io_deq_bits_qos),
    .io_deq_bits_region(r_queue_io_deq_bits_region),
    .io_deq_bits_id(r_queue_io_deq_bits_id),
    .io_deq_bits_user(r_queue_io_deq_bits_user),
    .io_count(r_queue_io_count)
  );
  Queue_55 b_queue (
    .clk(b_queue_clk),
    .reset(b_queue_reset),
    .io_enq_ready(b_queue_io_enq_ready),
    .io_enq_valid(b_queue_io_enq_valid),
    .io_enq_bits(b_queue_io_enq_bits),
    .io_deq_ready(b_queue_io_deq_ready),
    .io_deq_valid(b_queue_io_deq_valid),
    .io_deq_bits(b_queue_io_deq_bits),
    .io_count(b_queue_io_count)
  );
  assign io_aw_ready = T_374;
  assign io_w_ready = draining;
  assign io_b_valid = T_377;
  assign io_b_bits_resp = 2'h3;
  assign io_b_bits_id = b_queue_io_deq_bits;
  assign io_b_bits_user = GEN_9;
  assign io_ar_ready = r_queue_io_enq_ready;
  assign io_r_valid = T_347;
  assign io_r_bits_resp = 2'h3;
  assign io_r_bits_data = {{63'd0}, 1'h0};
  assign io_r_bits_last = T_350;
  assign io_r_bits_id = r_queue_io_deq_bits_id;
  assign io_r_bits_user = GEN_11;
  assign T_323 = io_ar_ready & io_ar_valid;
  assign T_325 = reset == 1'h0;
  assign T_326 = io_aw_ready & io_aw_valid;
  assign r_queue_clk = clk;
  assign r_queue_reset = reset;
  assign r_queue_io_enq_valid = io_ar_valid;
  assign r_queue_io_enq_bits_addr = io_ar_bits_addr;
  assign r_queue_io_enq_bits_len = io_ar_bits_len;
  assign r_queue_io_enq_bits_size = io_ar_bits_size;
  assign r_queue_io_enq_bits_burst = io_ar_bits_burst;
  assign r_queue_io_enq_bits_lock = io_ar_bits_lock;
  assign r_queue_io_enq_bits_cache = io_ar_bits_cache;
  assign r_queue_io_enq_bits_prot = io_ar_bits_prot;
  assign r_queue_io_enq_bits_qos = io_ar_bits_qos;
  assign r_queue_io_enq_bits_region = io_ar_bits_region;
  assign r_queue_io_enq_bits_id = io_ar_bits_id;
  assign r_queue_io_enq_bits_user = io_ar_bits_user;
  assign r_queue_io_deq_ready = T_352;
  assign T_344 = responding == 1'h0;
  assign T_345 = T_344 & r_queue_io_deq_valid;
  assign GEN_0 = T_345 ? 1'h1 : responding;
  assign GEN_1 = T_345 ? r_queue_io_deq_bits_len : beats_left;
  assign T_347 = r_queue_io_deq_valid & responding;
  assign GEN_8 = {{7'd0}, 1'h0};
  assign T_350 = beats_left == GEN_8;
  assign T_351 = io_r_ready & io_r_valid;
  assign T_352 = T_351 & io_r_bits_last;
  assign GEN_2 = T_350 ? 1'h0 : GEN_0;
  assign T_358 = T_350 == 1'h0;
  assign GEN_10 = {{7'd0}, 1'h1};
  assign T_360 = beats_left - GEN_10;
  assign T_361 = T_360[7:0];
  assign GEN_3 = T_358 ? T_361 : GEN_1;
  assign GEN_4 = T_351 ? GEN_2 : GEN_0;
  assign GEN_5 = T_351 ? GEN_3 : GEN_1;
  assign GEN_6 = T_326 ? 1'h1 : draining;
  assign T_365 = io_w_ready & io_w_valid;
  assign T_366 = T_365 & io_w_bits_last;
  assign GEN_7 = T_366 ? 1'h0 : GEN_6;
  assign b_queue_clk = clk;
  assign b_queue_reset = reset;
  assign b_queue_io_enq_valid = T_371;
  assign b_queue_io_enq_bits = io_aw_bits_id;
  assign b_queue_io_deq_ready = T_381;
  assign T_370 = draining == 1'h0;
  assign T_371 = io_aw_valid & T_370;
  assign T_374 = b_queue_io_enq_ready & T_370;
  assign T_377 = b_queue_io_deq_valid & T_370;
  assign T_381 = io_b_ready & T_370;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_12 = {1{$random}};
  responding = GEN_12[0:0];
  GEN_13 = {1{$random}};
  beats_left = GEN_13[7:0];
  GEN_14 = {1{$random}};
  draining = GEN_14[0:0];
  GEN_15 = {1{$random}};
  GEN_9 = GEN_15[0:0];
  GEN_16 = {1{$random}};
  GEN_11 = GEN_16[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      responding <= 1'h0;
    end else begin
      responding <= GEN_4;
    end
    if(reset) begin
      beats_left <= 8'h0;
    end else begin
      beats_left <= GEN_5;
    end
    if(reset) begin
      draining <= 1'h0;
    end else begin
      draining <= GEN_7;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_323 & T_325) begin
          $fwrite(32'h80000002,"Invalid read address %h\n",io_ar_bits_addr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_326 & T_325) begin
          $fwrite(32'h80000002,"Invalid write address %h\n",io_aw_bits_addr);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module ReorderQueue_57(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_data_addr_beat,
  input   io_enq_bits_data_subblock,
  input  [4:0] io_enq_bits_tag,
  input   io_deq_valid,
  input  [4:0] io_deq_tag,
  output [2:0] io_deq_data_addr_beat,
  output  io_deq_data_subblock,
  output  io_deq_matches
);
  reg [2:0] roq_data_addr_beat [0:3];
  reg [31:0] GEN_11;
  wire [2:0] roq_data_addr_beat_T_254_data;
  wire [1:0] roq_data_addr_beat_T_254_addr;
  wire  roq_data_addr_beat_T_254_en;
  wire [2:0] roq_data_addr_beat_T_276_data;
  wire [1:0] roq_data_addr_beat_T_276_addr;
  wire  roq_data_addr_beat_T_276_mask;
  wire  roq_data_addr_beat_T_276_en;
  reg  roq_data_subblock [0:3];
  reg [31:0] GEN_12;
  wire  roq_data_subblock_T_254_data;
  wire [1:0] roq_data_subblock_T_254_addr;
  wire  roq_data_subblock_T_254_en;
  wire  roq_data_subblock_T_276_data;
  wire [1:0] roq_data_subblock_T_276_addr;
  wire  roq_data_subblock_T_276_mask;
  wire  roq_data_subblock_T_276_en;
  reg [4:0] roq_tags_0;
  reg [31:0] GEN_13;
  reg [4:0] roq_tags_1;
  reg [31:0] GEN_14;
  reg [4:0] roq_tags_2;
  reg [31:0] GEN_15;
  reg [4:0] roq_tags_3;
  reg [31:0] GEN_16;
  wire  T_218_0;
  wire  T_218_1;
  wire  T_218_2;
  wire  T_218_3;
  reg  roq_free_0;
  reg [31:0] GEN_17;
  reg  roq_free_1;
  reg [31:0] GEN_18;
  reg  roq_free_2;
  reg [31:0] GEN_23;
  reg  roq_free_3;
  reg [31:0] GEN_32;
  wire [1:0] T_227;
  wire [1:0] T_228;
  wire [1:0] roq_enq_addr;
  wire  T_229;
  wire  T_231;
  wire  T_232;
  wire  T_233;
  wire  T_235;
  wire  T_236;
  wire  T_237;
  wire  T_239;
  wire  T_240;
  wire  T_241;
  wire  T_243;
  wire  T_244;
  wire [1:0] T_249;
  wire [1:0] T_250;
  wire [1:0] roq_deq_addr;
  wire  T_251;
  wire  T_252;
  wire  T_253;
  wire  T_272;
  wire  T_273;
  wire  T_274;
  wire  T_275;
  wire [4:0] GEN_0;
  wire [1:0] GEN_37;
  wire [4:0] GEN_3;
  wire [1:0] GEN_38;
  wire [4:0] GEN_4;
  wire [4:0] GEN_5;
  wire [4:0] GEN_6;
  wire  GEN_1;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [4:0] GEN_19;
  wire [4:0] GEN_20;
  wire [4:0] GEN_21;
  wire [4:0] GEN_22;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_2;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  assign io_enq_ready = T_253;
  assign io_deq_data_addr_beat = roq_data_addr_beat_T_254_data;
  assign io_deq_data_subblock = roq_data_subblock_T_254_data;
  assign io_deq_matches = T_274;
  assign roq_data_addr_beat_T_254_addr = roq_deq_addr;
  assign roq_data_addr_beat_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_addr_beat_T_254_data = roq_data_addr_beat[roq_data_addr_beat_T_254_addr];
  `else
  assign roq_data_addr_beat_T_254_data = roq_data_addr_beat_T_254_addr >= 3'h4 ? $random : roq_data_addr_beat[roq_data_addr_beat_T_254_addr];
  `endif
  assign roq_data_addr_beat_T_276_data = io_enq_bits_data_addr_beat;
  assign roq_data_addr_beat_T_276_addr = roq_enq_addr;
  assign roq_data_addr_beat_T_276_mask = T_275;
  assign roq_data_addr_beat_T_276_en = T_275;
  assign roq_data_subblock_T_254_addr = roq_deq_addr;
  assign roq_data_subblock_T_254_en = 1'h1;
  `ifdef SYNTHESIS
  assign roq_data_subblock_T_254_data = roq_data_subblock[roq_data_subblock_T_254_addr];
  `else
  assign roq_data_subblock_T_254_data = roq_data_subblock_T_254_addr >= 3'h4 ? $random : roq_data_subblock[roq_data_subblock_T_254_addr];
  `endif
  assign roq_data_subblock_T_276_data = io_enq_bits_data_subblock;
  assign roq_data_subblock_T_276_addr = roq_enq_addr;
  assign roq_data_subblock_T_276_mask = T_275;
  assign roq_data_subblock_T_276_en = T_275;
  assign T_218_0 = 1'h1;
  assign T_218_1 = 1'h1;
  assign T_218_2 = 1'h1;
  assign T_218_3 = 1'h1;
  assign T_227 = roq_free_2 ? 2'h2 : 2'h3;
  assign T_228 = roq_free_1 ? {{1'd0}, 1'h1} : T_227;
  assign roq_enq_addr = roq_free_0 ? {{1'd0}, 1'h0} : T_228;
  assign T_229 = roq_tags_0 == io_deq_tag;
  assign T_231 = roq_free_0 == 1'h0;
  assign T_232 = T_229 & T_231;
  assign T_233 = roq_tags_1 == io_deq_tag;
  assign T_235 = roq_free_1 == 1'h0;
  assign T_236 = T_233 & T_235;
  assign T_237 = roq_tags_2 == io_deq_tag;
  assign T_239 = roq_free_2 == 1'h0;
  assign T_240 = T_237 & T_239;
  assign T_241 = roq_tags_3 == io_deq_tag;
  assign T_243 = roq_free_3 == 1'h0;
  assign T_244 = T_241 & T_243;
  assign T_249 = T_240 ? 2'h2 : 2'h3;
  assign T_250 = T_236 ? {{1'd0}, 1'h1} : T_249;
  assign roq_deq_addr = T_232 ? {{1'd0}, 1'h0} : T_250;
  assign T_251 = roq_free_0 | roq_free_1;
  assign T_252 = T_251 | roq_free_2;
  assign T_253 = T_252 | roq_free_3;
  assign T_272 = T_232 | T_236;
  assign T_273 = T_272 | T_240;
  assign T_274 = T_273 | T_244;
  assign T_275 = io_enq_valid & io_enq_ready;
  assign GEN_0 = io_enq_bits_tag;
  assign GEN_37 = {{1'd0}, 1'h0};
  assign GEN_3 = GEN_37 == roq_enq_addr ? GEN_0 : roq_tags_0;
  assign GEN_38 = {{1'd0}, 1'h1};
  assign GEN_4 = GEN_38 == roq_enq_addr ? GEN_0 : roq_tags_1;
  assign GEN_5 = 2'h2 == roq_enq_addr ? GEN_0 : roq_tags_2;
  assign GEN_6 = 2'h3 == roq_enq_addr ? GEN_0 : roq_tags_3;
  assign GEN_1 = 1'h0;
  assign GEN_7 = GEN_37 == roq_enq_addr ? GEN_1 : roq_free_0;
  assign GEN_8 = GEN_38 == roq_enq_addr ? GEN_1 : roq_free_1;
  assign GEN_9 = 2'h2 == roq_enq_addr ? GEN_1 : roq_free_2;
  assign GEN_10 = 2'h3 == roq_enq_addr ? GEN_1 : roq_free_3;
  assign GEN_19 = T_275 ? GEN_3 : roq_tags_0;
  assign GEN_20 = T_275 ? GEN_4 : roq_tags_1;
  assign GEN_21 = T_275 ? GEN_5 : roq_tags_2;
  assign GEN_22 = T_275 ? GEN_6 : roq_tags_3;
  assign GEN_24 = T_275 ? GEN_7 : roq_free_0;
  assign GEN_25 = T_275 ? GEN_8 : roq_free_1;
  assign GEN_26 = T_275 ? GEN_9 : roq_free_2;
  assign GEN_27 = T_275 ? GEN_10 : roq_free_3;
  assign GEN_2 = 1'h1;
  assign GEN_28 = GEN_37 == roq_deq_addr ? GEN_2 : GEN_24;
  assign GEN_29 = GEN_38 == roq_deq_addr ? GEN_2 : GEN_25;
  assign GEN_30 = 2'h2 == roq_deq_addr ? GEN_2 : GEN_26;
  assign GEN_31 = 2'h3 == roq_deq_addr ? GEN_2 : GEN_27;
  assign GEN_33 = io_deq_valid ? GEN_28 : GEN_24;
  assign GEN_34 = io_deq_valid ? GEN_29 : GEN_25;
  assign GEN_35 = io_deq_valid ? GEN_30 : GEN_26;
  assign GEN_36 = io_deq_valid ? GEN_31 : GEN_27;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_11 = {1{$random}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    roq_data_addr_beat[initvar] = GEN_11[2:0];
  GEN_12 = {1{$random}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    roq_data_subblock[initvar] = GEN_12[0:0];
  GEN_13 = {1{$random}};
  roq_tags_0 = GEN_13[4:0];
  GEN_14 = {1{$random}};
  roq_tags_1 = GEN_14[4:0];
  GEN_15 = {1{$random}};
  roq_tags_2 = GEN_15[4:0];
  GEN_16 = {1{$random}};
  roq_tags_3 = GEN_16[4:0];
  GEN_17 = {1{$random}};
  roq_free_0 = GEN_17[0:0];
  GEN_18 = {1{$random}};
  roq_free_1 = GEN_18[0:0];
  GEN_23 = {1{$random}};
  roq_free_2 = GEN_23[0:0];
  GEN_32 = {1{$random}};
  roq_free_3 = GEN_32[0:0];
  end
`endif
  always @(posedge clk) begin
    if(roq_data_addr_beat_T_276_en & roq_data_addr_beat_T_276_mask) begin
      roq_data_addr_beat[roq_data_addr_beat_T_276_addr] <= roq_data_addr_beat_T_276_data;
    end
    if(roq_data_subblock_T_276_en & roq_data_subblock_T_276_mask) begin
      roq_data_subblock[roq_data_subblock_T_276_addr] <= roq_data_subblock_T_276_data;
    end
    if(1'h0) begin
    end else begin
      roq_tags_0 <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      roq_tags_1 <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      roq_tags_2 <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      roq_tags_3 <= GEN_22;
    end
    if(reset) begin
      roq_free_0 <= T_218_0;
    end else begin
      roq_free_0 <= GEN_33;
    end
    if(reset) begin
      roq_free_1 <= T_218_1;
    end else begin
      roq_free_1 <= GEN_34;
    end
    if(reset) begin
      roq_free_2 <= T_218_2;
    end else begin
      roq_free_2 <= GEN_35;
    end
    if(reset) begin
      roq_free_3 <= T_218_3;
    end else begin
      roq_free_3 <= GEN_36;
    end
  end
endmodule
module NastiIOTileLinkIOIdMapper_58(
  input   clk,
  input   reset,
  input   io_req_valid,
  output  io_req_ready,
  input  [1:0] io_req_tl_id,
  output [4:0] io_req_nasti_id,
  input   io_resp_valid,
  output  io_resp_matches,
  input  [4:0] io_resp_nasti_id,
  output [1:0] io_resp_tl_id
);
  assign io_req_ready = 1'h1;
  assign io_req_nasti_id = {{3'd0}, io_req_tl_id};
  assign io_resp_matches = 1'h1;
  assign io_resp_tl_id = io_resp_nasti_id[1:0];
endmodule
module Arbiter_60(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_is_builtin_type,
  input  [3:0] io_in_0_bits_g_type,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_client_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_is_builtin_type,
  input  [3:0] io_in_1_bits_g_type,
  input  [63:0] io_in_1_bits_data,
  input   io_in_1_bits_client_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_client_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [1:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire [63:0] GEN_6;
  wire  GEN_7;
  wire  T_542;
  wire  T_544;
  wire  T_546;
  wire  T_547;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_544;
  assign io_out_valid = T_547;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_manager_xact_id = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_g_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_client_id = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_manager_xact_id : io_in_1_bits_manager_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_is_builtin_type : io_in_1_bits_is_builtin_type;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_g_type : io_in_1_bits_g_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_client_id : io_in_1_bits_client_id;
  assign T_542 = io_in_0_valid == 1'h0;
  assign T_544 = T_542 & io_out_ready;
  assign T_546 = T_542 == 1'h0;
  assign T_547 = T_546 | io_in_1_valid;
endmodule
module NastiIOTileLinkIOConverter_56(
  input   clk,
  input   reset,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data,
  input   io_nasti_aw_ready,
  output  io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  output [7:0] io_nasti_aw_bits_len,
  output [2:0] io_nasti_aw_bits_size,
  output [1:0] io_nasti_aw_bits_burst,
  output  io_nasti_aw_bits_lock,
  output [3:0] io_nasti_aw_bits_cache,
  output [2:0] io_nasti_aw_bits_prot,
  output [3:0] io_nasti_aw_bits_qos,
  output [3:0] io_nasti_aw_bits_region,
  output [4:0] io_nasti_aw_bits_id,
  output  io_nasti_aw_bits_user,
  input   io_nasti_w_ready,
  output  io_nasti_w_valid,
  output [63:0] io_nasti_w_bits_data,
  output  io_nasti_w_bits_last,
  output [4:0] io_nasti_w_bits_id,
  output [7:0] io_nasti_w_bits_strb,
  output  io_nasti_w_bits_user,
  output  io_nasti_b_ready,
  input   io_nasti_b_valid,
  input  [1:0] io_nasti_b_bits_resp,
  input  [4:0] io_nasti_b_bits_id,
  input   io_nasti_b_bits_user,
  input   io_nasti_ar_ready,
  output  io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output [7:0] io_nasti_ar_bits_len,
  output [2:0] io_nasti_ar_bits_size,
  output [1:0] io_nasti_ar_bits_burst,
  output  io_nasti_ar_bits_lock,
  output [3:0] io_nasti_ar_bits_cache,
  output [2:0] io_nasti_ar_bits_prot,
  output [3:0] io_nasti_ar_bits_qos,
  output [3:0] io_nasti_ar_bits_region,
  output [4:0] io_nasti_ar_bits_id,
  output  io_nasti_ar_bits_user,
  output  io_nasti_r_ready,
  input   io_nasti_r_valid,
  input  [1:0] io_nasti_r_bits_resp,
  input  [63:0] io_nasti_r_bits_data,
  input   io_nasti_r_bits_last,
  input  [4:0] io_nasti_r_bits_id,
  input   io_nasti_r_bits_user
);
  wire [2:0] T_593_0;
  wire [2:0] T_593_1;
  wire [2:0] T_593_2;
  wire  T_595;
  wire  T_596;
  wire  T_597;
  wire  T_600;
  wire  T_601;
  wire  has_data;
  wire [2:0] T_610_0;
  wire [2:0] T_610_1;
  wire [2:0] T_610_2;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire  T_617;
  wire  T_618;
  wire  is_subblock;
  wire [2:0] T_627_0;
  wire  T_629;
  wire  is_multibeat;
  wire  T_632;
  wire  T_633;
  reg [2:0] tl_cnt_out;
  reg [31:0] GEN_15;
  wire  T_636;
  wire [2:0] GEN_6;
  wire [3:0] T_638;
  wire [2:0] T_639;
  wire [2:0] GEN_0;
  wire  tl_wrap_out;
  wire  T_641;
  wire  get_valid;
  wire  put_valid;
  wire  roq_clk;
  wire  roq_reset;
  wire  roq_io_enq_ready;
  wire  roq_io_enq_valid;
  wire [2:0] roq_io_enq_bits_data_addr_beat;
  wire  roq_io_enq_bits_data_subblock;
  wire [4:0] roq_io_enq_bits_tag;
  wire  roq_io_deq_valid;
  wire [4:0] roq_io_deq_tag;
  wire [2:0] roq_io_deq_data_addr_beat;
  wire  roq_io_deq_data_subblock;
  wire  roq_io_deq_matches;
  wire  get_id_mapper_clk;
  wire  get_id_mapper_reset;
  wire  get_id_mapper_io_req_valid;
  wire  get_id_mapper_io_req_ready;
  wire [1:0] get_id_mapper_io_req_tl_id;
  wire [4:0] get_id_mapper_io_req_nasti_id;
  wire  get_id_mapper_io_resp_valid;
  wire  get_id_mapper_io_resp_matches;
  wire [4:0] get_id_mapper_io_resp_nasti_id;
  wire [1:0] get_id_mapper_io_resp_tl_id;
  wire  put_id_mapper_clk;
  wire  put_id_mapper_reset;
  wire  put_id_mapper_io_req_valid;
  wire  put_id_mapper_io_req_ready;
  wire [1:0] put_id_mapper_io_req_tl_id;
  wire [4:0] put_id_mapper_io_req_nasti_id;
  wire  put_id_mapper_io_resp_valid;
  wire  put_id_mapper_io_resp_matches;
  wire [4:0] put_id_mapper_io_resp_nasti_id;
  wire [1:0] put_id_mapper_io_resp_tl_id;
  wire [2:0] GEN_7;
  wire  T_661;
  wire  put_id_mask;
  wire  T_663;
  wire  put_id_ready;
  reg  w_inflight;
  reg [31:0] GEN_16;
  wire  aw_ready;
  wire  T_665;
  wire  T_667;
  wire  T_668;
  reg [2:0] nasti_cnt_out;
  reg [31:0] GEN_17;
  wire  T_671;
  wire [3:0] T_673;
  wire [2:0] T_674;
  wire [2:0] GEN_1;
  wire  nasti_wrap_out;
  wire  T_675;
  wire  T_676;
  wire  T_678;
  wire  T_679;
  wire  T_680;
  wire  T_681;
  wire  T_683;
  wire  T_684;
  wire  T_685;
  wire  T_686;
  wire  T_687;
  wire  T_689;
  wire [2:0] T_690;
  wire [28:0] T_691;
  wire [31:0] T_692;
  wire [2:0] T_693;
  wire  T_703;
  wire [2:0] T_704;
  wire  T_705;
  wire [2:0] T_706;
  wire  T_707;
  wire [2:0] T_708;
  wire  T_709;
  wire [2:0] T_710;
  wire  T_711;
  wire [2:0] T_712;
  wire  T_713;
  wire [2:0] T_714;
  wire  T_715;
  wire [2:0] T_716;
  wire  T_717;
  wire [2:0] T_718;
  wire [2:0] T_720;
  wire [2:0] T_723;
  wire [31:0] T_736_addr;
  wire [7:0] T_736_len;
  wire [2:0] T_736_size;
  wire [1:0] T_736_burst;
  wire  T_736_lock;
  wire [3:0] T_736_cache;
  wire [2:0] T_736_prot;
  wire [3:0] T_736_qos;
  wire [3:0] T_736_region;
  wire [4:0] T_736_id;
  wire  T_736_user;
  wire  T_755;
  wire  T_756;
  wire  T_757;
  wire  T_758;
  wire [2:0] T_765;
  wire [31:0] T_778_addr;
  wire [7:0] T_778_len;
  wire [2:0] T_778_size;
  wire [1:0] T_778_burst;
  wire  T_778_lock;
  wire [3:0] T_778_cache;
  wire [2:0] T_778_prot;
  wire [3:0] T_778_qos;
  wire [3:0] T_778_region;
  wire [4:0] T_778_id;
  wire  T_778_user;
  wire  T_797;
  wire  T_799;
  wire  T_800;
  wire [7:0] GEN_9;
  wire [8:0] T_804;
  wire [7:0] T_805;
  wire [7:0] T_811_0;
  wire  T_814;
  wire  T_815;
  wire  T_817;
  wire  T_818;
  wire  T_819;
  wire [7:0] T_820;
  wire [7:0] T_822;
  wire [7:0] T_823;
  wire  T_825;
  wire  T_826;
  wire [63:0] T_833_data;
  wire  T_833_last;
  wire [4:0] T_833_id;
  wire [7:0] T_833_strb;
  wire  T_833_user;
  wire  T_844;
  wire  T_845;
  wire  T_846;
  wire  T_847;
  wire  T_848;
  wire  T_852;
  wire  T_853;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  T_856;
  wire [2:0] T_864_0;
  wire [3:0] GEN_10;
  wire  T_866;
  wire  T_874_0;
  wire [3:0] GEN_11;
  wire  T_876;
  wire  T_879;
  wire  T_881;
  reg [2:0] tl_cnt_in;
  reg [31:0] GEN_18;
  wire [3:0] T_886;
  wire [2:0] T_887;
  wire [2:0] GEN_5;
  wire  gnt_arb_clk;
  wire  gnt_arb_reset;
  wire  gnt_arb_io_in_0_ready;
  wire  gnt_arb_io_in_0_valid;
  wire [2:0] gnt_arb_io_in_0_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_0_bits_client_xact_id;
  wire  gnt_arb_io_in_0_bits_manager_xact_id;
  wire  gnt_arb_io_in_0_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_0_bits_g_type;
  wire [63:0] gnt_arb_io_in_0_bits_data;
  wire  gnt_arb_io_in_0_bits_client_id;
  wire  gnt_arb_io_in_1_ready;
  wire  gnt_arb_io_in_1_valid;
  wire [2:0] gnt_arb_io_in_1_bits_addr_beat;
  wire [1:0] gnt_arb_io_in_1_bits_client_xact_id;
  wire  gnt_arb_io_in_1_bits_manager_xact_id;
  wire  gnt_arb_io_in_1_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_in_1_bits_g_type;
  wire [63:0] gnt_arb_io_in_1_bits_data;
  wire  gnt_arb_io_in_1_bits_client_id;
  wire  gnt_arb_io_out_ready;
  wire  gnt_arb_io_out_valid;
  wire [2:0] gnt_arb_io_out_bits_addr_beat;
  wire [1:0] gnt_arb_io_out_bits_client_xact_id;
  wire  gnt_arb_io_out_bits_manager_xact_id;
  wire  gnt_arb_io_out_bits_is_builtin_type;
  wire [3:0] gnt_arb_io_out_bits_g_type;
  wire [63:0] gnt_arb_io_out_bits_data;
  wire  gnt_arb_io_out_bits_client_id;
  wire  gnt_arb_io_chosen;
  wire [2:0] T_914;
  wire [2:0] T_916;
  wire [2:0] T_939_addr_beat;
  wire [1:0] T_939_client_xact_id;
  wire  T_939_manager_xact_id;
  wire  T_939_is_builtin_type;
  wire [3:0] T_939_g_type;
  wire [63:0] T_939_data;
  wire  T_962;
  wire  T_963;
  wire  T_964;
  wire  T_966;
  wire  T_969;
  wire  T_970;
  wire  T_972;
  wire [2:0] T_1000_addr_beat;
  wire [1:0] T_1000_client_xact_id;
  wire  T_1000_manager_xact_id;
  wire  T_1000_is_builtin_type;
  wire [3:0] T_1000_g_type;
  wire [63:0] T_1000_data;
  wire  T_1023;
  wire  T_1024;
  wire  T_1025;
  wire  T_1027;
  wire  T_1029;
  wire [1:0] GEN_13;
  wire  T_1031;
  wire  T_1032;
  wire  T_1033;
  wire  T_1035;
  wire  T_1037;
  wire  T_1039;
  wire  T_1040;
  wire  T_1041;
  wire  T_1043;
  reg [4:0] GEN_8;
  reg [31:0] GEN_19;
  reg  GEN_12;
  reg [31:0] GEN_20;
  reg  GEN_14;
  reg [31:0] GEN_21;
  ReorderQueue_57 roq (
    .clk(roq_clk),
    .reset(roq_reset),
    .io_enq_ready(roq_io_enq_ready),
    .io_enq_valid(roq_io_enq_valid),
    .io_enq_bits_data_addr_beat(roq_io_enq_bits_data_addr_beat),
    .io_enq_bits_data_subblock(roq_io_enq_bits_data_subblock),
    .io_enq_bits_tag(roq_io_enq_bits_tag),
    .io_deq_valid(roq_io_deq_valid),
    .io_deq_tag(roq_io_deq_tag),
    .io_deq_data_addr_beat(roq_io_deq_data_addr_beat),
    .io_deq_data_subblock(roq_io_deq_data_subblock),
    .io_deq_matches(roq_io_deq_matches)
  );
  NastiIOTileLinkIOIdMapper_58 get_id_mapper (
    .clk(get_id_mapper_clk),
    .reset(get_id_mapper_reset),
    .io_req_valid(get_id_mapper_io_req_valid),
    .io_req_ready(get_id_mapper_io_req_ready),
    .io_req_tl_id(get_id_mapper_io_req_tl_id),
    .io_req_nasti_id(get_id_mapper_io_req_nasti_id),
    .io_resp_valid(get_id_mapper_io_resp_valid),
    .io_resp_matches(get_id_mapper_io_resp_matches),
    .io_resp_nasti_id(get_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(get_id_mapper_io_resp_tl_id)
  );
  NastiIOTileLinkIOIdMapper_58 put_id_mapper (
    .clk(put_id_mapper_clk),
    .reset(put_id_mapper_reset),
    .io_req_valid(put_id_mapper_io_req_valid),
    .io_req_ready(put_id_mapper_io_req_ready),
    .io_req_tl_id(put_id_mapper_io_req_tl_id),
    .io_req_nasti_id(put_id_mapper_io_req_nasti_id),
    .io_resp_valid(put_id_mapper_io_resp_valid),
    .io_resp_matches(put_id_mapper_io_resp_matches),
    .io_resp_nasti_id(put_id_mapper_io_resp_nasti_id),
    .io_resp_tl_id(put_id_mapper_io_resp_tl_id)
  );
  Arbiter_60 gnt_arb (
    .clk(gnt_arb_clk),
    .reset(gnt_arb_reset),
    .io_in_0_ready(gnt_arb_io_in_0_ready),
    .io_in_0_valid(gnt_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(gnt_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_client_xact_id(gnt_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_manager_xact_id(gnt_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_is_builtin_type(gnt_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_g_type(gnt_arb_io_in_0_bits_g_type),
    .io_in_0_bits_data(gnt_arb_io_in_0_bits_data),
    .io_in_0_bits_client_id(gnt_arb_io_in_0_bits_client_id),
    .io_in_1_ready(gnt_arb_io_in_1_ready),
    .io_in_1_valid(gnt_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(gnt_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_client_xact_id(gnt_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_manager_xact_id(gnt_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_is_builtin_type(gnt_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_g_type(gnt_arb_io_in_1_bits_g_type),
    .io_in_1_bits_data(gnt_arb_io_in_1_bits_data),
    .io_in_1_bits_client_id(gnt_arb_io_in_1_bits_client_id),
    .io_out_ready(gnt_arb_io_out_ready),
    .io_out_valid(gnt_arb_io_out_valid),
    .io_out_bits_addr_beat(gnt_arb_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(gnt_arb_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(gnt_arb_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(gnt_arb_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(gnt_arb_io_out_bits_g_type),
    .io_out_bits_data(gnt_arb_io_out_bits_data),
    .io_out_bits_client_id(gnt_arb_io_out_bits_client_id),
    .io_chosen(gnt_arb_io_chosen)
  );
  assign io_tl_acquire_ready = T_848;
  assign io_tl_grant_valid = gnt_arb_io_out_valid;
  assign io_tl_grant_bits_addr_beat = gnt_arb_io_out_bits_addr_beat;
  assign io_tl_grant_bits_client_xact_id = gnt_arb_io_out_bits_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = gnt_arb_io_out_bits_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = gnt_arb_io_out_bits_is_builtin_type;
  assign io_tl_grant_bits_g_type = gnt_arb_io_out_bits_g_type;
  assign io_tl_grant_bits_data = gnt_arb_io_out_bits_data;
  assign io_nasti_aw_valid = T_758;
  assign io_nasti_aw_bits_addr = T_778_addr;
  assign io_nasti_aw_bits_len = T_778_len;
  assign io_nasti_aw_bits_size = T_778_size;
  assign io_nasti_aw_bits_burst = T_778_burst;
  assign io_nasti_aw_bits_lock = T_778_lock;
  assign io_nasti_aw_bits_cache = T_778_cache;
  assign io_nasti_aw_bits_prot = T_778_prot;
  assign io_nasti_aw_bits_qos = T_778_qos;
  assign io_nasti_aw_bits_region = T_778_region;
  assign io_nasti_aw_bits_id = T_778_id;
  assign io_nasti_aw_bits_user = T_778_user;
  assign io_nasti_w_valid = T_797;
  assign io_nasti_w_bits_data = T_833_data;
  assign io_nasti_w_bits_last = T_833_last;
  assign io_nasti_w_bits_id = T_833_id;
  assign io_nasti_w_bits_strb = T_833_strb;
  assign io_nasti_w_bits_user = T_833_user;
  assign io_nasti_b_ready = gnt_arb_io_in_1_ready;
  assign io_nasti_ar_valid = T_689;
  assign io_nasti_ar_bits_addr = T_736_addr;
  assign io_nasti_ar_bits_len = T_736_len;
  assign io_nasti_ar_bits_size = T_736_size;
  assign io_nasti_ar_bits_burst = T_736_burst;
  assign io_nasti_ar_bits_lock = T_736_lock;
  assign io_nasti_ar_bits_cache = T_736_cache;
  assign io_nasti_ar_bits_prot = T_736_prot;
  assign io_nasti_ar_bits_qos = T_736_qos;
  assign io_nasti_ar_bits_region = T_736_region;
  assign io_nasti_ar_bits_id = T_736_id;
  assign io_nasti_ar_bits_user = T_736_user;
  assign io_nasti_r_ready = gnt_arb_io_in_0_ready;
  assign T_593_0 = 3'h2;
  assign T_593_1 = 3'h3;
  assign T_593_2 = 3'h4;
  assign T_595 = T_593_0 == io_tl_acquire_bits_a_type;
  assign T_596 = T_593_1 == io_tl_acquire_bits_a_type;
  assign T_597 = T_593_2 == io_tl_acquire_bits_a_type;
  assign T_600 = T_595 | T_596;
  assign T_601 = T_600 | T_597;
  assign has_data = io_tl_acquire_bits_is_builtin_type & T_601;
  assign T_610_0 = 3'h2;
  assign T_610_1 = 3'h0;
  assign T_610_2 = 3'h4;
  assign T_612 = T_610_0 == io_tl_acquire_bits_a_type;
  assign T_613 = T_610_1 == io_tl_acquire_bits_a_type;
  assign T_614 = T_610_2 == io_tl_acquire_bits_a_type;
  assign T_617 = T_612 | T_613;
  assign T_618 = T_617 | T_614;
  assign is_subblock = io_tl_acquire_bits_is_builtin_type & T_618;
  assign T_627_0 = 3'h3;
  assign T_629 = T_627_0 == io_tl_acquire_bits_a_type;
  assign is_multibeat = io_tl_acquire_bits_is_builtin_type & T_629;
  assign T_632 = io_tl_acquire_ready & io_tl_acquire_valid;
  assign T_633 = T_632 & is_multibeat;
  assign T_636 = tl_cnt_out == 3'h7;
  assign GEN_6 = {{2'd0}, 1'h1};
  assign T_638 = tl_cnt_out + GEN_6;
  assign T_639 = T_638[2:0];
  assign GEN_0 = T_633 ? T_639 : tl_cnt_out;
  assign tl_wrap_out = T_633 & T_636;
  assign T_641 = has_data == 1'h0;
  assign get_valid = io_tl_acquire_valid & T_641;
  assign put_valid = io_tl_acquire_valid & has_data;
  assign roq_clk = clk;
  assign roq_reset = reset;
  assign roq_io_enq_valid = T_676;
  assign roq_io_enq_bits_data_addr_beat = io_tl_acquire_bits_addr_beat;
  assign roq_io_enq_bits_data_subblock = is_subblock;
  assign roq_io_enq_bits_tag = io_nasti_ar_bits_id;
  assign roq_io_deq_valid = T_679;
  assign roq_io_deq_tag = io_nasti_r_bits_id;
  assign get_id_mapper_clk = clk;
  assign get_id_mapper_reset = reset;
  assign get_id_mapper_io_req_valid = T_681;
  assign get_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign get_id_mapper_io_resp_valid = T_683;
  assign get_id_mapper_io_resp_nasti_id = io_nasti_r_bits_id;
  assign put_id_mapper_clk = clk;
  assign put_id_mapper_reset = reset;
  assign put_id_mapper_io_req_valid = T_686;
  assign put_id_mapper_io_req_tl_id = io_tl_acquire_bits_client_xact_id;
  assign put_id_mapper_io_resp_valid = T_687;
  assign put_id_mapper_io_resp_nasti_id = io_nasti_b_bits_id;
  assign GEN_7 = {{2'd0}, 1'h0};
  assign T_661 = io_tl_acquire_bits_addr_beat == GEN_7;
  assign put_id_mask = is_subblock | T_661;
  assign T_663 = put_id_mask == 1'h0;
  assign put_id_ready = put_id_mapper_io_req_ready | T_663;
  assign aw_ready = w_inflight | io_nasti_aw_ready;
  assign T_665 = io_nasti_r_ready & io_nasti_r_valid;
  assign T_667 = roq_io_deq_data_subblock == 1'h0;
  assign T_668 = T_665 & T_667;
  assign T_671 = nasti_cnt_out == 3'h7;
  assign T_673 = nasti_cnt_out + GEN_6;
  assign T_674 = T_673[2:0];
  assign GEN_1 = T_668 ? T_674 : nasti_cnt_out;
  assign nasti_wrap_out = T_668 & T_671;
  assign T_675 = get_valid & io_nasti_ar_ready;
  assign T_676 = T_675 & get_id_mapper_io_req_ready;
  assign T_678 = nasti_wrap_out | roq_io_deq_data_subblock;
  assign T_679 = T_665 & T_678;
  assign T_680 = get_valid & roq_io_enq_ready;
  assign T_681 = T_680 & io_nasti_ar_ready;
  assign T_683 = T_665 & io_nasti_r_bits_last;
  assign T_684 = put_valid & aw_ready;
  assign T_685 = T_684 & io_nasti_w_ready;
  assign T_686 = T_685 & put_id_mask;
  assign T_687 = io_nasti_b_ready & io_nasti_b_valid;
  assign T_689 = T_680 & get_id_mapper_io_req_ready;
  assign T_690 = io_tl_acquire_bits_union[11:9];
  assign T_691 = {io_tl_acquire_bits_addr_block,io_tl_acquire_bits_addr_beat};
  assign T_692 = {T_691,T_690};
  assign T_693 = io_tl_acquire_bits_union[8:6];
  assign T_703 = 3'h7 == T_693;
  assign T_704 = T_703 ? {{1'd0}, 2'h3} : 3'h7;
  assign T_705 = 3'h3 == T_693;
  assign T_706 = T_705 ? {{1'd0}, 2'h3} : T_704;
  assign T_707 = 3'h6 == T_693;
  assign T_708 = T_707 ? {{1'd0}, 2'h2} : T_706;
  assign T_709 = 3'h2 == T_693;
  assign T_710 = T_709 ? {{1'd0}, 2'h2} : T_708;
  assign T_711 = 3'h5 == T_693;
  assign T_712 = T_711 ? {{2'd0}, 1'h1} : T_710;
  assign T_713 = 3'h1 == T_693;
  assign T_714 = T_713 ? {{2'd0}, 1'h1} : T_712;
  assign T_715 = 3'h4 == T_693;
  assign T_716 = T_715 ? {{2'd0}, 1'h0} : T_714;
  assign T_717 = 3'h0 == T_693;
  assign T_718 = T_717 ? {{2'd0}, 1'h0} : T_716;
  assign T_720 = is_subblock ? T_718 : {{1'd0}, 2'h3};
  assign T_723 = is_subblock ? {{2'd0}, 1'h0} : 3'h7;
  assign T_736_addr = T_692;
  assign T_736_len = {{5'd0}, T_723};
  assign T_736_size = T_720;
  assign T_736_burst = 2'h1;
  assign T_736_lock = 1'h0;
  assign T_736_cache = {{3'd0}, 1'h0};
  assign T_736_prot = {{2'd0}, 1'h0};
  assign T_736_qos = {{3'd0}, 1'h0};
  assign T_736_region = {{3'd0}, 1'h0};
  assign T_736_id = get_id_mapper_io_req_nasti_id;
  assign T_736_user = 1'h0;
  assign T_755 = w_inflight == 1'h0;
  assign T_756 = put_valid & io_nasti_w_ready;
  assign T_757 = T_756 & put_id_ready;
  assign T_758 = T_757 & T_755;
  assign T_765 = is_multibeat ? 3'h7 : {{2'd0}, 1'h0};
  assign T_778_addr = T_692;
  assign T_778_len = {{5'd0}, T_765};
  assign T_778_size = {{1'd0}, 2'h3};
  assign T_778_burst = 2'h1;
  assign T_778_lock = 1'h0;
  assign T_778_cache = 4'h0;
  assign T_778_prot = 3'h0;
  assign T_778_qos = 4'h0;
  assign T_778_region = 4'h0;
  assign T_778_id = put_id_mapper_io_req_nasti_id;
  assign T_778_user = 1'h0;
  assign T_797 = T_684 & put_id_ready;
  assign T_799 = io_tl_acquire_bits_a_type == 3'h4;
  assign T_800 = io_tl_acquire_bits_is_builtin_type & T_799;
  assign GEN_9 = {{7'd0}, 1'h1};
  assign T_804 = 8'h0 - GEN_9;
  assign T_805 = T_804[7:0];
  assign T_811_0 = T_805;
  assign T_814 = io_tl_acquire_bits_a_type == 3'h3;
  assign T_815 = io_tl_acquire_bits_is_builtin_type & T_814;
  assign T_817 = io_tl_acquire_bits_a_type == 3'h2;
  assign T_818 = io_tl_acquire_bits_is_builtin_type & T_817;
  assign T_819 = T_815 | T_818;
  assign T_820 = io_tl_acquire_bits_union[8:1];
  assign T_822 = T_819 ? T_820 : {{7'd0}, 1'h0};
  assign T_823 = T_800 ? T_811_0 : T_822;
  assign T_825 = T_632 & is_subblock;
  assign T_826 = tl_wrap_out | T_825;
  assign T_833_data = io_tl_acquire_bits_data;
  assign T_833_last = T_826;
  assign T_833_id = GEN_8;
  assign T_833_strb = T_823;
  assign T_833_user = 1'h0;
  assign T_844 = aw_ready & io_nasti_w_ready;
  assign T_845 = T_844 & put_id_ready;
  assign T_846 = roq_io_enq_ready & io_nasti_ar_ready;
  assign T_847 = T_846 & get_id_mapper_io_req_ready;
  assign T_848 = has_data ? T_845 : T_847;
  assign T_852 = T_755 & T_632;
  assign T_853 = T_852 & is_multibeat;
  assign GEN_2 = T_853 ? 1'h1 : w_inflight;
  assign GEN_3 = tl_wrap_out ? 1'h0 : GEN_2;
  assign GEN_4 = w_inflight ? GEN_3 : GEN_2;
  assign T_856 = io_tl_grant_ready & io_tl_grant_valid;
  assign T_864_0 = 3'h5;
  assign GEN_10 = {{1'd0}, T_864_0};
  assign T_866 = GEN_10 == io_tl_grant_bits_g_type;
  assign T_874_0 = 1'h0;
  assign GEN_11 = {{3'd0}, T_874_0};
  assign T_876 = GEN_11 == io_tl_grant_bits_g_type;
  assign T_879 = io_tl_grant_bits_is_builtin_type ? T_866 : T_876;
  assign T_881 = T_856 & T_879;
  assign T_886 = tl_cnt_in + GEN_6;
  assign T_887 = T_886[2:0];
  assign GEN_5 = T_881 ? T_887 : tl_cnt_in;
  assign gnt_arb_clk = clk;
  assign gnt_arb_reset = reset;
  assign gnt_arb_io_in_0_valid = io_nasti_r_valid;
  assign gnt_arb_io_in_0_bits_addr_beat = T_939_addr_beat;
  assign gnt_arb_io_in_0_bits_client_xact_id = T_939_client_xact_id;
  assign gnt_arb_io_in_0_bits_manager_xact_id = T_939_manager_xact_id;
  assign gnt_arb_io_in_0_bits_is_builtin_type = T_939_is_builtin_type;
  assign gnt_arb_io_in_0_bits_g_type = T_939_g_type;
  assign gnt_arb_io_in_0_bits_data = T_939_data;
  assign gnt_arb_io_in_0_bits_client_id = GEN_12;
  assign gnt_arb_io_in_1_valid = io_nasti_b_valid;
  assign gnt_arb_io_in_1_bits_addr_beat = T_1000_addr_beat;
  assign gnt_arb_io_in_1_bits_client_xact_id = T_1000_client_xact_id;
  assign gnt_arb_io_in_1_bits_manager_xact_id = T_1000_manager_xact_id;
  assign gnt_arb_io_in_1_bits_is_builtin_type = T_1000_is_builtin_type;
  assign gnt_arb_io_in_1_bits_g_type = T_1000_g_type;
  assign gnt_arb_io_in_1_bits_data = T_1000_data;
  assign gnt_arb_io_in_1_bits_client_id = GEN_14;
  assign gnt_arb_io_out_ready = io_tl_grant_ready;
  assign T_914 = roq_io_deq_data_subblock ? 3'h4 : 3'h5;
  assign T_916 = roq_io_deq_data_subblock ? roq_io_deq_data_addr_beat : tl_cnt_in;
  assign T_939_addr_beat = T_916;
  assign T_939_client_xact_id = get_id_mapper_io_resp_tl_id;
  assign T_939_manager_xact_id = 1'h0;
  assign T_939_is_builtin_type = 1'h1;
  assign T_939_g_type = {{1'd0}, T_914};
  assign T_939_data = io_nasti_r_bits_data;
  assign T_962 = gnt_arb_io_in_0_valid == 1'h0;
  assign T_963 = T_962 | roq_io_deq_matches;
  assign T_964 = T_963 | reset;
  assign T_966 = T_964 == 1'h0;
  assign T_969 = T_962 | get_id_mapper_io_resp_matches;
  assign T_970 = T_969 | reset;
  assign T_972 = T_970 == 1'h0;
  assign T_1000_addr_beat = {{2'd0}, 1'h0};
  assign T_1000_client_xact_id = put_id_mapper_io_resp_tl_id;
  assign T_1000_manager_xact_id = 1'h0;
  assign T_1000_is_builtin_type = 1'h1;
  assign T_1000_g_type = {{1'd0}, 3'h3};
  assign T_1000_data = {{63'd0}, 1'h0};
  assign T_1023 = gnt_arb_io_in_1_valid == 1'h0;
  assign T_1024 = T_1023 | put_id_mapper_io_resp_matches;
  assign T_1025 = T_1024 | reset;
  assign T_1027 = T_1025 == 1'h0;
  assign T_1029 = io_nasti_r_valid == 1'h0;
  assign GEN_13 = {{1'd0}, 1'h0};
  assign T_1031 = io_nasti_r_bits_resp == GEN_13;
  assign T_1032 = T_1029 | T_1031;
  assign T_1033 = T_1032 | reset;
  assign T_1035 = T_1033 == 1'h0;
  assign T_1037 = io_nasti_b_valid == 1'h0;
  assign T_1039 = io_nasti_b_bits_resp == GEN_13;
  assign T_1040 = T_1037 | T_1039;
  assign T_1041 = T_1040 | reset;
  assign T_1043 = T_1041 == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_15 = {1{$random}};
  tl_cnt_out = GEN_15[2:0];
  GEN_16 = {1{$random}};
  w_inflight = GEN_16[0:0];
  GEN_17 = {1{$random}};
  nasti_cnt_out = GEN_17[2:0];
  GEN_18 = {1{$random}};
  tl_cnt_in = GEN_18[2:0];
  GEN_19 = {1{$random}};
  GEN_8 = GEN_19[4:0];
  GEN_20 = {1{$random}};
  GEN_12 = GEN_20[0:0];
  GEN_21 = {1{$random}};
  GEN_14 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      tl_cnt_out <= 3'h0;
    end else begin
      tl_cnt_out <= GEN_0;
    end
    if(reset) begin
      w_inflight <= 1'h0;
    end else begin
      w_inflight <= GEN_4;
    end
    if(reset) begin
      nasti_cnt_out <= 3'h0;
    end else begin
      nasti_cnt_out <= GEN_1;
    end
    if(reset) begin
      tl_cnt_in <= 3'h0;
    end else begin
      tl_cnt_in <= GEN_5;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_966) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:609 assert(!gnt_arb.io.in(0).valid || roq.io.deq.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_966) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_972) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:610 assert(!gnt_arb.io.in(0).valid || get_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_972) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1027) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI tag error\n    at converters.scala:621 assert(!gnt_arb.io.in(1).valid || put_id_mapper.io.resp.matches, \"NASTI tag error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1027) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1035) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI read error\n    at converters.scala:623 assert(!io.nasti.r.valid || io.nasti.r.bits.resp === UInt(0), \"NASTI read error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1035) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1043) begin
          $fwrite(32'h80000002,"Assertion failed: NASTI write error\n    at converters.scala:624 assert(!io.nasti.b.valid || io.nasti.b.bits.resp === UInt(0), \"NASTI write error\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1043) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module Uncore(
  input   clk,
  input   reset,
  output  io_host_clk,
  output  io_host_clk_edge,
  output  io_host_in_ready,
  input   io_host_in_valid,
  input  [15:0] io_host_in_bits,
  input   io_host_out_ready,
  output  io_host_out_valid,
  output [15:0] io_host_out_bits,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  output  io_tiles_cached_0_acquire_ready,
  input   io_tiles_cached_0_acquire_valid,
  input  [25:0] io_tiles_cached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_cached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_cached_0_acquire_bits_addr_beat,
  input   io_tiles_cached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_cached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_cached_0_acquire_bits_union,
  input  [63:0] io_tiles_cached_0_acquire_bits_data,
  input   io_tiles_cached_0_probe_ready,
  output  io_tiles_cached_0_probe_valid,
  output [25:0] io_tiles_cached_0_probe_bits_addr_block,
  output [1:0] io_tiles_cached_0_probe_bits_p_type,
  output  io_tiles_cached_0_release_ready,
  input   io_tiles_cached_0_release_valid,
  input  [2:0] io_tiles_cached_0_release_bits_addr_beat,
  input  [25:0] io_tiles_cached_0_release_bits_addr_block,
  input  [1:0] io_tiles_cached_0_release_bits_client_xact_id,
  input   io_tiles_cached_0_release_bits_voluntary,
  input  [2:0] io_tiles_cached_0_release_bits_r_type,
  input  [63:0] io_tiles_cached_0_release_bits_data,
  input   io_tiles_cached_0_grant_ready,
  output  io_tiles_cached_0_grant_valid,
  output [2:0] io_tiles_cached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_cached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_cached_0_grant_bits_manager_xact_id,
  output  io_tiles_cached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_cached_0_grant_bits_g_type,
  output [63:0] io_tiles_cached_0_grant_bits_data,
  output  io_tiles_cached_0_grant_bits_manager_id,
  output  io_tiles_cached_0_finish_ready,
  input   io_tiles_cached_0_finish_valid,
  input  [2:0] io_tiles_cached_0_finish_bits_manager_xact_id,
  input   io_tiles_cached_0_finish_bits_manager_id,
  output  io_tiles_uncached_0_acquire_ready,
  input   io_tiles_uncached_0_acquire_valid,
  input  [25:0] io_tiles_uncached_0_acquire_bits_addr_block,
  input  [1:0] io_tiles_uncached_0_acquire_bits_client_xact_id,
  input  [2:0] io_tiles_uncached_0_acquire_bits_addr_beat,
  input   io_tiles_uncached_0_acquire_bits_is_builtin_type,
  input  [2:0] io_tiles_uncached_0_acquire_bits_a_type,
  input  [11:0] io_tiles_uncached_0_acquire_bits_union,
  input  [63:0] io_tiles_uncached_0_acquire_bits_data,
  input   io_tiles_uncached_0_grant_ready,
  output  io_tiles_uncached_0_grant_valid,
  output [2:0] io_tiles_uncached_0_grant_bits_addr_beat,
  output [1:0] io_tiles_uncached_0_grant_bits_client_xact_id,
  output [2:0] io_tiles_uncached_0_grant_bits_manager_xact_id,
  output  io_tiles_uncached_0_grant_bits_is_builtin_type,
  output [3:0] io_tiles_uncached_0_grant_bits_g_type,
  output [63:0] io_tiles_uncached_0_grant_bits_data,
  output  io_prci_0_reset,
  output  io_prci_0_id,
  output  io_prci_0_interrupts_mtip,
  output  io_prci_0_interrupts_meip,
  output  io_prci_0_interrupts_seip,
  output  io_prci_0_interrupts_debug,
  output  io_prci_0_interrupts_msip,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debugBus_req_ready,
  input   io_debugBus_req_valid,
  input  [4:0] io_debugBus_req_bits_addr,
  input  [1:0] io_debugBus_req_bits_op,
  input  [33:0] io_debugBus_req_bits_data,
  input   io_debugBus_resp_ready,
  output  io_debugBus_resp_valid,
  output [1:0] io_debugBus_resp_bits_resp,
  output [33:0] io_debugBus_resp_bits_data
);
  wire  htif_clk;
  wire  htif_reset;
  wire  htif_io_host_clk;
  wire  htif_io_host_clk_edge;
  wire  htif_io_host_in_ready;
  wire  htif_io_host_in_valid;
  wire [15:0] htif_io_host_in_bits;
  wire  htif_io_host_out_ready;
  wire  htif_io_host_out_valid;
  wire [15:0] htif_io_host_out_bits;
  wire  htif_io_cpu_0_reset;
  wire  htif_io_cpu_0_id;
  wire  htif_io_cpu_0_csr_req_ready;
  wire  htif_io_cpu_0_csr_req_valid;
  wire  htif_io_cpu_0_csr_req_bits_rw;
  wire [11:0] htif_io_cpu_0_csr_req_bits_addr;
  wire [63:0] htif_io_cpu_0_csr_req_bits_data;
  wire  htif_io_cpu_0_csr_resp_ready;
  wire  htif_io_cpu_0_csr_resp_valid;
  wire [63:0] htif_io_cpu_0_csr_resp_bits;
  wire  htif_io_mem_acquire_ready;
  wire  htif_io_mem_acquire_valid;
  wire [25:0] htif_io_mem_acquire_bits_addr_block;
  wire [1:0] htif_io_mem_acquire_bits_client_xact_id;
  wire [2:0] htif_io_mem_acquire_bits_addr_beat;
  wire  htif_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] htif_io_mem_acquire_bits_a_type;
  wire [11:0] htif_io_mem_acquire_bits_union;
  wire [63:0] htif_io_mem_acquire_bits_data;
  wire  htif_io_mem_grant_ready;
  wire  htif_io_mem_grant_valid;
  wire [2:0] htif_io_mem_grant_bits_addr_beat;
  wire [1:0] htif_io_mem_grant_bits_client_xact_id;
  wire [2:0] htif_io_mem_grant_bits_manager_xact_id;
  wire  htif_io_mem_grant_bits_is_builtin_type;
  wire [3:0] htif_io_mem_grant_bits_g_type;
  wire [63:0] htif_io_mem_grant_bits_data;
  wire  htif_io_scr_req_ready;
  wire  htif_io_scr_req_valid;
  wire  htif_io_scr_req_bits_rw;
  wire [5:0] htif_io_scr_req_bits_addr;
  wire [63:0] htif_io_scr_req_bits_data;
  wire  htif_io_scr_resp_ready;
  wire  htif_io_scr_resp_valid;
  wire [63:0] htif_io_scr_resp_bits;
  wire  outmemsys_clk;
  wire  outmemsys_reset;
  wire  outmemsys_io_tiles_cached_0_acquire_ready;
  wire  outmemsys_io_tiles_cached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_cached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_cached_0_probe_ready;
  wire  outmemsys_io_tiles_cached_0_probe_valid;
  wire [25:0] outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_probe_bits_p_type;
  wire  outmemsys_io_tiles_cached_0_release_ready;
  wire  outmemsys_io_tiles_cached_0_release_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] outmemsys_io_tiles_cached_0_release_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_cached_0_release_bits_client_xact_id;
  wire  outmemsys_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] outmemsys_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] outmemsys_io_tiles_cached_0_release_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_ready;
  wire  outmemsys_io_tiles_cached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_cached_0_grant_bits_data;
  wire  outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  wire  outmemsys_io_tiles_cached_0_finish_ready;
  wire  outmemsys_io_tiles_cached_0_finish_valid;
  wire [2:0] outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  outmemsys_io_tiles_cached_0_finish_bits_manager_id;
  wire  outmemsys_io_tiles_uncached_0_acquire_ready;
  wire  outmemsys_io_tiles_uncached_0_acquire_valid;
  wire [25:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] outmemsys_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] outmemsys_io_tiles_uncached_0_acquire_bits_data;
  wire  outmemsys_io_tiles_uncached_0_grant_ready;
  wire  outmemsys_io_tiles_uncached_0_grant_valid;
  wire [2:0] outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [2:0] outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] outmemsys_io_tiles_uncached_0_grant_bits_data;
  wire  outmemsys_io_htif_uncached_acquire_ready;
  wire  outmemsys_io_htif_uncached_acquire_valid;
  wire [25:0] outmemsys_io_htif_uncached_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_htif_uncached_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_htif_uncached_acquire_bits_addr_beat;
  wire  outmemsys_io_htif_uncached_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_htif_uncached_acquire_bits_a_type;
  wire [11:0] outmemsys_io_htif_uncached_acquire_bits_union;
  wire [63:0] outmemsys_io_htif_uncached_acquire_bits_data;
  wire  outmemsys_io_htif_uncached_grant_ready;
  wire  outmemsys_io_htif_uncached_grant_valid;
  wire [2:0] outmemsys_io_htif_uncached_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  wire [2:0] outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  wire  outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_htif_uncached_grant_bits_g_type;
  wire [63:0] outmemsys_io_htif_uncached_grant_bits_data;
  wire  outmemsys_io_incoherent_0;
  wire  outmemsys_io_mem_axi_0_aw_ready;
  wire  outmemsys_io_mem_axi_0_aw_valid;
  wire [31:0] outmemsys_io_mem_axi_0_aw_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_aw_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_aw_bits_burst;
  wire  outmemsys_io_mem_axi_0_aw_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_aw_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_aw_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_aw_bits_id;
  wire  outmemsys_io_mem_axi_0_aw_bits_user;
  wire  outmemsys_io_mem_axi_0_w_ready;
  wire  outmemsys_io_mem_axi_0_w_valid;
  wire [63:0] outmemsys_io_mem_axi_0_w_bits_data;
  wire  outmemsys_io_mem_axi_0_w_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_w_bits_id;
  wire [7:0] outmemsys_io_mem_axi_0_w_bits_strb;
  wire  outmemsys_io_mem_axi_0_w_bits_user;
  wire  outmemsys_io_mem_axi_0_b_ready;
  wire  outmemsys_io_mem_axi_0_b_valid;
  wire [1:0] outmemsys_io_mem_axi_0_b_bits_resp;
  wire [4:0] outmemsys_io_mem_axi_0_b_bits_id;
  wire  outmemsys_io_mem_axi_0_b_bits_user;
  wire  outmemsys_io_mem_axi_0_ar_ready;
  wire  outmemsys_io_mem_axi_0_ar_valid;
  wire [31:0] outmemsys_io_mem_axi_0_ar_bits_addr;
  wire [7:0] outmemsys_io_mem_axi_0_ar_bits_len;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_size;
  wire [1:0] outmemsys_io_mem_axi_0_ar_bits_burst;
  wire  outmemsys_io_mem_axi_0_ar_bits_lock;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_cache;
  wire [2:0] outmemsys_io_mem_axi_0_ar_bits_prot;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_qos;
  wire [3:0] outmemsys_io_mem_axi_0_ar_bits_region;
  wire [4:0] outmemsys_io_mem_axi_0_ar_bits_id;
  wire  outmemsys_io_mem_axi_0_ar_bits_user;
  wire  outmemsys_io_mem_axi_0_r_ready;
  wire  outmemsys_io_mem_axi_0_r_valid;
  wire [1:0] outmemsys_io_mem_axi_0_r_bits_resp;
  wire [63:0] outmemsys_io_mem_axi_0_r_bits_data;
  wire  outmemsys_io_mem_axi_0_r_bits_last;
  wire [4:0] outmemsys_io_mem_axi_0_r_bits_id;
  wire  outmemsys_io_mem_axi_0_r_bits_user;
  wire  outmemsys_io_mmio_acquire_ready;
  wire  outmemsys_io_mmio_acquire_valid;
  wire [25:0] outmemsys_io_mmio_acquire_bits_addr_block;
  wire [1:0] outmemsys_io_mmio_acquire_bits_client_xact_id;
  wire [2:0] outmemsys_io_mmio_acquire_bits_addr_beat;
  wire  outmemsys_io_mmio_acquire_bits_is_builtin_type;
  wire [2:0] outmemsys_io_mmio_acquire_bits_a_type;
  wire [11:0] outmemsys_io_mmio_acquire_bits_union;
  wire [63:0] outmemsys_io_mmio_acquire_bits_data;
  wire  outmemsys_io_mmio_grant_ready;
  wire  outmemsys_io_mmio_grant_valid;
  wire [2:0] outmemsys_io_mmio_grant_bits_addr_beat;
  wire [1:0] outmemsys_io_mmio_grant_bits_client_xact_id;
  wire  outmemsys_io_mmio_grant_bits_manager_xact_id;
  wire  outmemsys_io_mmio_grant_bits_is_builtin_type;
  wire [3:0] outmemsys_io_mmio_grant_bits_g_type;
  wire [63:0] outmemsys_io_mmio_grant_bits_data;
  wire  scrFile_clk;
  wire  scrFile_reset;
  wire  scrFile_io_smi_req_ready;
  wire  scrFile_io_smi_req_valid;
  wire  scrFile_io_smi_req_bits_rw;
  wire [5:0] scrFile_io_smi_req_bits_addr;
  wire [63:0] scrFile_io_smi_req_bits_data;
  wire  scrFile_io_smi_resp_ready;
  wire  scrFile_io_smi_resp_valid;
  wire [63:0] scrFile_io_smi_resp_bits;
  wire [63:0] scrFile_io_scr_rdata_0;
  wire [63:0] scrFile_io_scr_rdata_1;
  wire [63:0] scrFile_io_scr_rdata_2;
  wire [63:0] scrFile_io_scr_rdata_3;
  wire [63:0] scrFile_io_scr_rdata_4;
  wire [63:0] scrFile_io_scr_rdata_5;
  wire [63:0] scrFile_io_scr_rdata_6;
  wire [63:0] scrFile_io_scr_rdata_7;
  wire [63:0] scrFile_io_scr_rdata_8;
  wire [63:0] scrFile_io_scr_rdata_9;
  wire [63:0] scrFile_io_scr_rdata_10;
  wire [63:0] scrFile_io_scr_rdata_11;
  wire [63:0] scrFile_io_scr_rdata_12;
  wire [63:0] scrFile_io_scr_rdata_13;
  wire [63:0] scrFile_io_scr_rdata_14;
  wire [63:0] scrFile_io_scr_rdata_15;
  wire [63:0] scrFile_io_scr_rdata_16;
  wire [63:0] scrFile_io_scr_rdata_17;
  wire [63:0] scrFile_io_scr_rdata_18;
  wire [63:0] scrFile_io_scr_rdata_19;
  wire [63:0] scrFile_io_scr_rdata_20;
  wire [63:0] scrFile_io_scr_rdata_21;
  wire [63:0] scrFile_io_scr_rdata_22;
  wire [63:0] scrFile_io_scr_rdata_23;
  wire [63:0] scrFile_io_scr_rdata_24;
  wire [63:0] scrFile_io_scr_rdata_25;
  wire [63:0] scrFile_io_scr_rdata_26;
  wire [63:0] scrFile_io_scr_rdata_27;
  wire [63:0] scrFile_io_scr_rdata_28;
  wire [63:0] scrFile_io_scr_rdata_29;
  wire [63:0] scrFile_io_scr_rdata_30;
  wire [63:0] scrFile_io_scr_rdata_31;
  wire [63:0] scrFile_io_scr_rdata_32;
  wire [63:0] scrFile_io_scr_rdata_33;
  wire [63:0] scrFile_io_scr_rdata_34;
  wire [63:0] scrFile_io_scr_rdata_35;
  wire [63:0] scrFile_io_scr_rdata_36;
  wire [63:0] scrFile_io_scr_rdata_37;
  wire [63:0] scrFile_io_scr_rdata_38;
  wire [63:0] scrFile_io_scr_rdata_39;
  wire [63:0] scrFile_io_scr_rdata_40;
  wire [63:0] scrFile_io_scr_rdata_41;
  wire [63:0] scrFile_io_scr_rdata_42;
  wire [63:0] scrFile_io_scr_rdata_43;
  wire [63:0] scrFile_io_scr_rdata_44;
  wire [63:0] scrFile_io_scr_rdata_45;
  wire [63:0] scrFile_io_scr_rdata_46;
  wire [63:0] scrFile_io_scr_rdata_47;
  wire [63:0] scrFile_io_scr_rdata_48;
  wire [63:0] scrFile_io_scr_rdata_49;
  wire [63:0] scrFile_io_scr_rdata_50;
  wire [63:0] scrFile_io_scr_rdata_51;
  wire [63:0] scrFile_io_scr_rdata_52;
  wire [63:0] scrFile_io_scr_rdata_53;
  wire [63:0] scrFile_io_scr_rdata_54;
  wire [63:0] scrFile_io_scr_rdata_55;
  wire [63:0] scrFile_io_scr_rdata_56;
  wire [63:0] scrFile_io_scr_rdata_57;
  wire [63:0] scrFile_io_scr_rdata_58;
  wire [63:0] scrFile_io_scr_rdata_59;
  wire [63:0] scrFile_io_scr_rdata_60;
  wire [63:0] scrFile_io_scr_rdata_61;
  wire [63:0] scrFile_io_scr_rdata_62;
  wire [63:0] scrFile_io_scr_rdata_63;
  wire  scrFile_io_scr_wen;
  wire [5:0] scrFile_io_scr_waddr;
  wire [63:0] scrFile_io_scr_wdata;
  wire  TileLinkRecursiveInterconnect_8716_clk;
  wire  TileLinkRecursiveInterconnect_8716_reset;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_acquire_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_acquire_valid;
  wire [25:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_block;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_client_xact_id;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_beat;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_is_builtin_type;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_a_type;
  wire [11:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_union;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_data;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_grant_ready;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_grant_valid;
  wire [2:0] TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_addr_beat;
  wire [1:0] TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_client_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_manager_xact_id;
  wire  TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_is_builtin_type;
  wire [3:0] TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_g_type;
  wire [63:0] TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_data;
  wire  RTC_8717_clk;
  wire  RTC_8717_reset;
  wire  RTC_8717_io_tl_acquire_ready;
  wire  RTC_8717_io_tl_acquire_valid;
  wire [25:0] RTC_8717_io_tl_acquire_bits_addr_block;
  wire [1:0] RTC_8717_io_tl_acquire_bits_client_xact_id;
  wire [2:0] RTC_8717_io_tl_acquire_bits_addr_beat;
  wire  RTC_8717_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] RTC_8717_io_tl_acquire_bits_a_type;
  wire [11:0] RTC_8717_io_tl_acquire_bits_union;
  wire [63:0] RTC_8717_io_tl_acquire_bits_data;
  wire  RTC_8717_io_tl_grant_ready;
  wire  RTC_8717_io_tl_grant_valid;
  wire [2:0] RTC_8717_io_tl_grant_bits_addr_beat;
  wire [1:0] RTC_8717_io_tl_grant_bits_client_xact_id;
  wire  RTC_8717_io_tl_grant_bits_manager_xact_id;
  wire  RTC_8717_io_tl_grant_bits_is_builtin_type;
  wire [3:0] RTC_8717_io_tl_grant_bits_g_type;
  wire [63:0] RTC_8717_io_tl_grant_bits_data;
  wire  RTC_8717_io_irqs_0;
  wire  PLIC_8718_clk;
  wire  PLIC_8718_reset;
  wire  PLIC_8718_io_devices_0_valid;
  wire  PLIC_8718_io_devices_0_ready;
  wire  PLIC_8718_io_devices_0_complete;
  wire  PLIC_8718_io_devices_1_valid;
  wire  PLIC_8718_io_devices_1_ready;
  wire  PLIC_8718_io_devices_1_complete;
  wire  PLIC_8718_io_harts_0;
  wire  PLIC_8718_io_harts_1;
  wire  PLIC_8718_io_tl_acquire_ready;
  wire  PLIC_8718_io_tl_acquire_valid;
  wire [25:0] PLIC_8718_io_tl_acquire_bits_addr_block;
  wire [1:0] PLIC_8718_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PLIC_8718_io_tl_acquire_bits_addr_beat;
  wire  PLIC_8718_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PLIC_8718_io_tl_acquire_bits_a_type;
  wire [11:0] PLIC_8718_io_tl_acquire_bits_union;
  wire [63:0] PLIC_8718_io_tl_acquire_bits_data;
  wire  PLIC_8718_io_tl_grant_ready;
  wire  PLIC_8718_io_tl_grant_valid;
  wire [2:0] PLIC_8718_io_tl_grant_bits_addr_beat;
  wire [1:0] PLIC_8718_io_tl_grant_bits_client_xact_id;
  wire  PLIC_8718_io_tl_grant_bits_manager_xact_id;
  wire  PLIC_8718_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PLIC_8718_io_tl_grant_bits_g_type;
  wire [63:0] PLIC_8718_io_tl_grant_bits_data;
  wire  LevelGateway_8719_clk;
  wire  LevelGateway_8719_reset;
  wire  LevelGateway_8719_io_interrupt;
  wire  LevelGateway_8719_io_plic_valid;
  wire  LevelGateway_8719_io_plic_ready;
  wire  LevelGateway_8719_io_plic_complete;
  wire  LevelGateway_51_8720_clk;
  wire  LevelGateway_51_8720_reset;
  wire  LevelGateway_51_8720_io_interrupt;
  wire  LevelGateway_51_8720_io_plic_valid;
  wire  LevelGateway_51_8720_io_plic_ready;
  wire  LevelGateway_51_8720_io_plic_complete;
  wire  DebugModule_8721_clk;
  wire  DebugModule_8721_reset;
  wire  DebugModule_8721_io_db_req_ready;
  wire  DebugModule_8721_io_db_req_valid;
  wire [4:0] DebugModule_8721_io_db_req_bits_addr;
  wire [1:0] DebugModule_8721_io_db_req_bits_op;
  wire [33:0] DebugModule_8721_io_db_req_bits_data;
  wire  DebugModule_8721_io_db_resp_ready;
  wire  DebugModule_8721_io_db_resp_valid;
  wire [1:0] DebugModule_8721_io_db_resp_bits_resp;
  wire [33:0] DebugModule_8721_io_db_resp_bits_data;
  wire  DebugModule_8721_io_debugInterrupts_0;
  wire  DebugModule_8721_io_tl_acquire_ready;
  wire  DebugModule_8721_io_tl_acquire_valid;
  wire [25:0] DebugModule_8721_io_tl_acquire_bits_addr_block;
  wire [1:0] DebugModule_8721_io_tl_acquire_bits_client_xact_id;
  wire [2:0] DebugModule_8721_io_tl_acquire_bits_addr_beat;
  wire  DebugModule_8721_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] DebugModule_8721_io_tl_acquire_bits_a_type;
  wire [11:0] DebugModule_8721_io_tl_acquire_bits_union;
  wire [63:0] DebugModule_8721_io_tl_acquire_bits_data;
  wire  DebugModule_8721_io_tl_grant_ready;
  wire  DebugModule_8721_io_tl_grant_valid;
  wire [2:0] DebugModule_8721_io_tl_grant_bits_addr_beat;
  wire [1:0] DebugModule_8721_io_tl_grant_bits_client_xact_id;
  wire  DebugModule_8721_io_tl_grant_bits_manager_xact_id;
  wire  DebugModule_8721_io_tl_grant_bits_is_builtin_type;
  wire [3:0] DebugModule_8721_io_tl_grant_bits_g_type;
  wire [63:0] DebugModule_8721_io_tl_grant_bits_data;
  wire  DebugModule_8721_io_ndreset;
  wire  DebugModule_8721_io_fullreset;
  wire  PRCI_8722_clk;
  wire  PRCI_8722_reset;
  wire  PRCI_8722_io_interrupts_0_mtip;
  wire  PRCI_8722_io_interrupts_0_meip;
  wire  PRCI_8722_io_interrupts_0_seip;
  wire  PRCI_8722_io_interrupts_0_debug;
  wire  PRCI_8722_io_tl_acquire_ready;
  wire  PRCI_8722_io_tl_acquire_valid;
  wire [25:0] PRCI_8722_io_tl_acquire_bits_addr_block;
  wire [1:0] PRCI_8722_io_tl_acquire_bits_client_xact_id;
  wire [2:0] PRCI_8722_io_tl_acquire_bits_addr_beat;
  wire  PRCI_8722_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] PRCI_8722_io_tl_acquire_bits_a_type;
  wire [11:0] PRCI_8722_io_tl_acquire_bits_union;
  wire [63:0] PRCI_8722_io_tl_acquire_bits_data;
  wire  PRCI_8722_io_tl_grant_ready;
  wire  PRCI_8722_io_tl_grant_valid;
  wire [2:0] PRCI_8722_io_tl_grant_bits_addr_beat;
  wire [1:0] PRCI_8722_io_tl_grant_bits_client_xact_id;
  wire  PRCI_8722_io_tl_grant_bits_manager_xact_id;
  wire  PRCI_8722_io_tl_grant_bits_is_builtin_type;
  wire [3:0] PRCI_8722_io_tl_grant_bits_g_type;
  wire [63:0] PRCI_8722_io_tl_grant_bits_data;
  wire  PRCI_8722_io_tiles_0_reset;
  wire  PRCI_8722_io_tiles_0_id;
  wire  PRCI_8722_io_tiles_0_interrupts_mtip;
  wire  PRCI_8722_io_tiles_0_interrupts_meip;
  wire  PRCI_8722_io_tiles_0_interrupts_seip;
  wire  PRCI_8722_io_tiles_0_interrupts_debug;
  wire  PRCI_8722_io_tiles_0_interrupts_msip;
  reg  T_8725;
  reg [31:0] GEN_66;
  reg  T_8726;
  reg [31:0] GEN_67;
  wire  T_8727;
  wire  ROMSlave_8728_clk;
  wire  ROMSlave_8728_reset;
  wire  ROMSlave_8728_io_acquire_ready;
  wire  ROMSlave_8728_io_acquire_valid;
  wire [25:0] ROMSlave_8728_io_acquire_bits_addr_block;
  wire [1:0] ROMSlave_8728_io_acquire_bits_client_xact_id;
  wire [2:0] ROMSlave_8728_io_acquire_bits_addr_beat;
  wire  ROMSlave_8728_io_acquire_bits_is_builtin_type;
  wire [2:0] ROMSlave_8728_io_acquire_bits_a_type;
  wire [11:0] ROMSlave_8728_io_acquire_bits_union;
  wire [63:0] ROMSlave_8728_io_acquire_bits_data;
  wire  ROMSlave_8728_io_grant_ready;
  wire  ROMSlave_8728_io_grant_valid;
  wire [2:0] ROMSlave_8728_io_grant_bits_addr_beat;
  wire [1:0] ROMSlave_8728_io_grant_bits_client_xact_id;
  wire  ROMSlave_8728_io_grant_bits_manager_xact_id;
  wire  ROMSlave_8728_io_grant_bits_is_builtin_type;
  wire [3:0] ROMSlave_8728_io_grant_bits_g_type;
  wire [63:0] ROMSlave_8728_io_grant_bits_data;
  wire  NastiErrorSlave_8729_clk;
  wire  NastiErrorSlave_8729_reset;
  wire  NastiErrorSlave_8729_io_aw_ready;
  wire  NastiErrorSlave_8729_io_aw_valid;
  wire [31:0] NastiErrorSlave_8729_io_aw_bits_addr;
  wire [7:0] NastiErrorSlave_8729_io_aw_bits_len;
  wire [2:0] NastiErrorSlave_8729_io_aw_bits_size;
  wire [1:0] NastiErrorSlave_8729_io_aw_bits_burst;
  wire  NastiErrorSlave_8729_io_aw_bits_lock;
  wire [3:0] NastiErrorSlave_8729_io_aw_bits_cache;
  wire [2:0] NastiErrorSlave_8729_io_aw_bits_prot;
  wire [3:0] NastiErrorSlave_8729_io_aw_bits_qos;
  wire [3:0] NastiErrorSlave_8729_io_aw_bits_region;
  wire [4:0] NastiErrorSlave_8729_io_aw_bits_id;
  wire  NastiErrorSlave_8729_io_aw_bits_user;
  wire  NastiErrorSlave_8729_io_w_ready;
  wire  NastiErrorSlave_8729_io_w_valid;
  wire [63:0] NastiErrorSlave_8729_io_w_bits_data;
  wire  NastiErrorSlave_8729_io_w_bits_last;
  wire [4:0] NastiErrorSlave_8729_io_w_bits_id;
  wire [7:0] NastiErrorSlave_8729_io_w_bits_strb;
  wire  NastiErrorSlave_8729_io_w_bits_user;
  wire  NastiErrorSlave_8729_io_b_ready;
  wire  NastiErrorSlave_8729_io_b_valid;
  wire [1:0] NastiErrorSlave_8729_io_b_bits_resp;
  wire [4:0] NastiErrorSlave_8729_io_b_bits_id;
  wire  NastiErrorSlave_8729_io_b_bits_user;
  wire  NastiErrorSlave_8729_io_ar_ready;
  wire  NastiErrorSlave_8729_io_ar_valid;
  wire [31:0] NastiErrorSlave_8729_io_ar_bits_addr;
  wire [7:0] NastiErrorSlave_8729_io_ar_bits_len;
  wire [2:0] NastiErrorSlave_8729_io_ar_bits_size;
  wire [1:0] NastiErrorSlave_8729_io_ar_bits_burst;
  wire  NastiErrorSlave_8729_io_ar_bits_lock;
  wire [3:0] NastiErrorSlave_8729_io_ar_bits_cache;
  wire [2:0] NastiErrorSlave_8729_io_ar_bits_prot;
  wire [3:0] NastiErrorSlave_8729_io_ar_bits_qos;
  wire [3:0] NastiErrorSlave_8729_io_ar_bits_region;
  wire [4:0] NastiErrorSlave_8729_io_ar_bits_id;
  wire  NastiErrorSlave_8729_io_ar_bits_user;
  wire  NastiErrorSlave_8729_io_r_ready;
  wire  NastiErrorSlave_8729_io_r_valid;
  wire [1:0] NastiErrorSlave_8729_io_r_bits_resp;
  wire [63:0] NastiErrorSlave_8729_io_r_bits_data;
  wire  NastiErrorSlave_8729_io_r_bits_last;
  wire [4:0] NastiErrorSlave_8729_io_r_bits_id;
  wire  NastiErrorSlave_8729_io_r_bits_user;
  wire  NastiIOTileLinkIOConverter_56_8730_clk;
  wire  NastiIOTileLinkIOConverter_56_8730_reset;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_valid;
  wire [25:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_block;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_client_xact_id;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_beat;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_is_builtin_type;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_a_type;
  wire [11:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_union;
  wire [63:0] NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_data;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_grant_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_grant_valid;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_addr_beat;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_client_xact_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_manager_xact_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_is_builtin_type;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_g_type;
  wire [63:0] NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_data;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_valid;
  wire [31:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_burst;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_user;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_w_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_w_valid;
  wire [63:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_data;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_id;
  wire [7:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_strb;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_user;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_b_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_b_valid;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_resp;
  wire [4:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_user;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_valid;
  wire [31:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_addr;
  wire [7:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_len;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_size;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_burst;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_lock;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_cache;
  wire [2:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_prot;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_qos;
  wire [3:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_region;
  wire [4:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_user;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_r_ready;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_r_valid;
  wire [1:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_resp;
  wire [63:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_data;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_last;
  wire [4:0] NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_id;
  wire  NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_user;
  wire  Queue_61_8743_clk;
  wire  Queue_61_8743_reset;
  wire  Queue_61_8743_io_enq_ready;
  wire  Queue_61_8743_io_enq_valid;
  wire [31:0] Queue_61_8743_io_enq_bits_addr;
  wire [7:0] Queue_61_8743_io_enq_bits_len;
  wire [2:0] Queue_61_8743_io_enq_bits_size;
  wire [1:0] Queue_61_8743_io_enq_bits_burst;
  wire  Queue_61_8743_io_enq_bits_lock;
  wire [3:0] Queue_61_8743_io_enq_bits_cache;
  wire [2:0] Queue_61_8743_io_enq_bits_prot;
  wire [3:0] Queue_61_8743_io_enq_bits_qos;
  wire [3:0] Queue_61_8743_io_enq_bits_region;
  wire [4:0] Queue_61_8743_io_enq_bits_id;
  wire  Queue_61_8743_io_enq_bits_user;
  wire  Queue_61_8743_io_deq_ready;
  wire  Queue_61_8743_io_deq_valid;
  wire [31:0] Queue_61_8743_io_deq_bits_addr;
  wire [7:0] Queue_61_8743_io_deq_bits_len;
  wire [2:0] Queue_61_8743_io_deq_bits_size;
  wire [1:0] Queue_61_8743_io_deq_bits_burst;
  wire  Queue_61_8743_io_deq_bits_lock;
  wire [3:0] Queue_61_8743_io_deq_bits_cache;
  wire [2:0] Queue_61_8743_io_deq_bits_prot;
  wire [3:0] Queue_61_8743_io_deq_bits_qos;
  wire [3:0] Queue_61_8743_io_deq_bits_region;
  wire [4:0] Queue_61_8743_io_deq_bits_id;
  wire  Queue_61_8743_io_deq_bits_user;
  wire  Queue_61_8743_io_count;
  wire  Queue_62_8756_clk;
  wire  Queue_62_8756_reset;
  wire  Queue_62_8756_io_enq_ready;
  wire  Queue_62_8756_io_enq_valid;
  wire [31:0] Queue_62_8756_io_enq_bits_addr;
  wire [7:0] Queue_62_8756_io_enq_bits_len;
  wire [2:0] Queue_62_8756_io_enq_bits_size;
  wire [1:0] Queue_62_8756_io_enq_bits_burst;
  wire  Queue_62_8756_io_enq_bits_lock;
  wire [3:0] Queue_62_8756_io_enq_bits_cache;
  wire [2:0] Queue_62_8756_io_enq_bits_prot;
  wire [3:0] Queue_62_8756_io_enq_bits_qos;
  wire [3:0] Queue_62_8756_io_enq_bits_region;
  wire [4:0] Queue_62_8756_io_enq_bits_id;
  wire  Queue_62_8756_io_enq_bits_user;
  wire  Queue_62_8756_io_deq_ready;
  wire  Queue_62_8756_io_deq_valid;
  wire [31:0] Queue_62_8756_io_deq_bits_addr;
  wire [7:0] Queue_62_8756_io_deq_bits_len;
  wire [2:0] Queue_62_8756_io_deq_bits_size;
  wire [1:0] Queue_62_8756_io_deq_bits_burst;
  wire  Queue_62_8756_io_deq_bits_lock;
  wire [3:0] Queue_62_8756_io_deq_bits_cache;
  wire [2:0] Queue_62_8756_io_deq_bits_prot;
  wire [3:0] Queue_62_8756_io_deq_bits_qos;
  wire [3:0] Queue_62_8756_io_deq_bits_region;
  wire [4:0] Queue_62_8756_io_deq_bits_id;
  wire  Queue_62_8756_io_deq_bits_user;
  wire  Queue_62_8756_io_count;
  wire  Queue_63_8763_clk;
  wire  Queue_63_8763_reset;
  wire  Queue_63_8763_io_enq_ready;
  wire  Queue_63_8763_io_enq_valid;
  wire [63:0] Queue_63_8763_io_enq_bits_data;
  wire  Queue_63_8763_io_enq_bits_last;
  wire [4:0] Queue_63_8763_io_enq_bits_id;
  wire [7:0] Queue_63_8763_io_enq_bits_strb;
  wire  Queue_63_8763_io_enq_bits_user;
  wire  Queue_63_8763_io_deq_ready;
  wire  Queue_63_8763_io_deq_valid;
  wire [63:0] Queue_63_8763_io_deq_bits_data;
  wire  Queue_63_8763_io_deq_bits_last;
  wire [4:0] Queue_63_8763_io_deq_bits_id;
  wire [7:0] Queue_63_8763_io_deq_bits_strb;
  wire  Queue_63_8763_io_deq_bits_user;
  wire [1:0] Queue_63_8763_io_count;
  wire  Queue_64_8770_clk;
  wire  Queue_64_8770_reset;
  wire  Queue_64_8770_io_enq_ready;
  wire  Queue_64_8770_io_enq_valid;
  wire [1:0] Queue_64_8770_io_enq_bits_resp;
  wire [63:0] Queue_64_8770_io_enq_bits_data;
  wire  Queue_64_8770_io_enq_bits_last;
  wire [4:0] Queue_64_8770_io_enq_bits_id;
  wire  Queue_64_8770_io_enq_bits_user;
  wire  Queue_64_8770_io_deq_ready;
  wire  Queue_64_8770_io_deq_valid;
  wire [1:0] Queue_64_8770_io_deq_bits_resp;
  wire [63:0] Queue_64_8770_io_deq_bits_data;
  wire  Queue_64_8770_io_deq_bits_last;
  wire [4:0] Queue_64_8770_io_deq_bits_id;
  wire  Queue_64_8770_io_deq_bits_user;
  wire [1:0] Queue_64_8770_io_count;
  wire  Queue_65_8775_clk;
  wire  Queue_65_8775_reset;
  wire  Queue_65_8775_io_enq_ready;
  wire  Queue_65_8775_io_enq_valid;
  wire [1:0] Queue_65_8775_io_enq_bits_resp;
  wire [4:0] Queue_65_8775_io_enq_bits_id;
  wire  Queue_65_8775_io_enq_bits_user;
  wire  Queue_65_8775_io_deq_ready;
  wire  Queue_65_8775_io_deq_valid;
  wire [1:0] Queue_65_8775_io_deq_bits_resp;
  wire [4:0] Queue_65_8775_io_deq_bits_id;
  wire  Queue_65_8775_io_deq_bits_user;
  wire  Queue_65_8775_io_count;
  reg  GEN_0;
  reg [31:0] GEN_68;
  reg [63:0] GEN_1;
  reg [63:0] GEN_69;
  reg [63:0] GEN_2;
  reg [63:0] GEN_70;
  reg [63:0] GEN_3;
  reg [63:0] GEN_71;
  reg [63:0] GEN_4;
  reg [63:0] GEN_72;
  reg [63:0] GEN_5;
  reg [63:0] GEN_73;
  reg [63:0] GEN_6;
  reg [63:0] GEN_74;
  reg [63:0] GEN_7;
  reg [63:0] GEN_75;
  reg [63:0] GEN_8;
  reg [63:0] GEN_76;
  reg [63:0] GEN_9;
  reg [63:0] GEN_77;
  reg [63:0] GEN_10;
  reg [63:0] GEN_78;
  reg [63:0] GEN_11;
  reg [63:0] GEN_79;
  reg [63:0] GEN_12;
  reg [63:0] GEN_80;
  reg [63:0] GEN_13;
  reg [63:0] GEN_81;
  reg [63:0] GEN_14;
  reg [63:0] GEN_82;
  reg [63:0] GEN_15;
  reg [63:0] GEN_83;
  reg [63:0] GEN_16;
  reg [63:0] GEN_84;
  reg [63:0] GEN_17;
  reg [63:0] GEN_85;
  reg [63:0] GEN_18;
  reg [63:0] GEN_86;
  reg [63:0] GEN_19;
  reg [63:0] GEN_87;
  reg [63:0] GEN_20;
  reg [63:0] GEN_88;
  reg [63:0] GEN_21;
  reg [63:0] GEN_89;
  reg [63:0] GEN_22;
  reg [63:0] GEN_90;
  reg [63:0] GEN_23;
  reg [63:0] GEN_91;
  reg [63:0] GEN_24;
  reg [63:0] GEN_92;
  reg [63:0] GEN_25;
  reg [63:0] GEN_93;
  reg [63:0] GEN_26;
  reg [63:0] GEN_94;
  reg [63:0] GEN_27;
  reg [63:0] GEN_95;
  reg [63:0] GEN_28;
  reg [63:0] GEN_96;
  reg [63:0] GEN_29;
  reg [63:0] GEN_97;
  reg [63:0] GEN_30;
  reg [63:0] GEN_98;
  reg [63:0] GEN_31;
  reg [63:0] GEN_99;
  reg [63:0] GEN_32;
  reg [63:0] GEN_100;
  reg [63:0] GEN_33;
  reg [63:0] GEN_101;
  reg [63:0] GEN_34;
  reg [63:0] GEN_102;
  reg [63:0] GEN_35;
  reg [63:0] GEN_103;
  reg [63:0] GEN_36;
  reg [63:0] GEN_104;
  reg [63:0] GEN_37;
  reg [63:0] GEN_105;
  reg [63:0] GEN_38;
  reg [63:0] GEN_106;
  reg [63:0] GEN_39;
  reg [63:0] GEN_107;
  reg [63:0] GEN_40;
  reg [63:0] GEN_108;
  reg [63:0] GEN_41;
  reg [63:0] GEN_109;
  reg [63:0] GEN_42;
  reg [63:0] GEN_110;
  reg [63:0] GEN_43;
  reg [63:0] GEN_111;
  reg [63:0] GEN_44;
  reg [63:0] GEN_112;
  reg [63:0] GEN_45;
  reg [63:0] GEN_113;
  reg [63:0] GEN_46;
  reg [63:0] GEN_114;
  reg [63:0] GEN_47;
  reg [63:0] GEN_115;
  reg [63:0] GEN_48;
  reg [63:0] GEN_116;
  reg [63:0] GEN_49;
  reg [63:0] GEN_117;
  reg [63:0] GEN_50;
  reg [63:0] GEN_118;
  reg [63:0] GEN_51;
  reg [63:0] GEN_119;
  reg [63:0] GEN_52;
  reg [63:0] GEN_120;
  reg [63:0] GEN_53;
  reg [63:0] GEN_121;
  reg [63:0] GEN_54;
  reg [63:0] GEN_122;
  reg [63:0] GEN_55;
  reg [63:0] GEN_123;
  reg [63:0] GEN_56;
  reg [63:0] GEN_124;
  reg [63:0] GEN_57;
  reg [63:0] GEN_125;
  reg [63:0] GEN_58;
  reg [63:0] GEN_126;
  reg [63:0] GEN_59;
  reg [63:0] GEN_127;
  reg [63:0] GEN_60;
  reg [63:0] GEN_128;
  reg [63:0] GEN_61;
  reg [63:0] GEN_129;
  reg [63:0] GEN_62;
  reg [63:0] GEN_130;
  reg [63:0] GEN_63;
  reg [63:0] GEN_131;
  reg [63:0] GEN_64;
  reg [63:0] GEN_132;
  reg [63:0] GEN_65;
  reg [63:0] GEN_133;
  Htif htif (
    .clk(htif_clk),
    .reset(htif_reset),
    .io_host_clk(htif_io_host_clk),
    .io_host_clk_edge(htif_io_host_clk_edge),
    .io_host_in_ready(htif_io_host_in_ready),
    .io_host_in_valid(htif_io_host_in_valid),
    .io_host_in_bits(htif_io_host_in_bits),
    .io_host_out_ready(htif_io_host_out_ready),
    .io_host_out_valid(htif_io_host_out_valid),
    .io_host_out_bits(htif_io_host_out_bits),
    .io_cpu_0_reset(htif_io_cpu_0_reset),
    .io_cpu_0_id(htif_io_cpu_0_id),
    .io_cpu_0_csr_req_ready(htif_io_cpu_0_csr_req_ready),
    .io_cpu_0_csr_req_valid(htif_io_cpu_0_csr_req_valid),
    .io_cpu_0_csr_req_bits_rw(htif_io_cpu_0_csr_req_bits_rw),
    .io_cpu_0_csr_req_bits_addr(htif_io_cpu_0_csr_req_bits_addr),
    .io_cpu_0_csr_req_bits_data(htif_io_cpu_0_csr_req_bits_data),
    .io_cpu_0_csr_resp_ready(htif_io_cpu_0_csr_resp_ready),
    .io_cpu_0_csr_resp_valid(htif_io_cpu_0_csr_resp_valid),
    .io_cpu_0_csr_resp_bits(htif_io_cpu_0_csr_resp_bits),
    .io_mem_acquire_ready(htif_io_mem_acquire_ready),
    .io_mem_acquire_valid(htif_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(htif_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(htif_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(htif_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(htif_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(htif_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(htif_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(htif_io_mem_acquire_bits_data),
    .io_mem_grant_ready(htif_io_mem_grant_ready),
    .io_mem_grant_valid(htif_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(htif_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(htif_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(htif_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(htif_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(htif_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(htif_io_mem_grant_bits_data),
    .io_scr_req_ready(htif_io_scr_req_ready),
    .io_scr_req_valid(htif_io_scr_req_valid),
    .io_scr_req_bits_rw(htif_io_scr_req_bits_rw),
    .io_scr_req_bits_addr(htif_io_scr_req_bits_addr),
    .io_scr_req_bits_data(htif_io_scr_req_bits_data),
    .io_scr_resp_ready(htif_io_scr_resp_ready),
    .io_scr_resp_valid(htif_io_scr_resp_valid),
    .io_scr_resp_bits(htif_io_scr_resp_bits)
  );
  OuterMemorySystem outmemsys (
    .clk(outmemsys_clk),
    .reset(outmemsys_reset),
    .io_tiles_cached_0_acquire_ready(outmemsys_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(outmemsys_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(outmemsys_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(outmemsys_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(outmemsys_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(outmemsys_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(outmemsys_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(outmemsys_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(outmemsys_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(outmemsys_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(outmemsys_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(outmemsys_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(outmemsys_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(outmemsys_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(outmemsys_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(outmemsys_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(outmemsys_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(outmemsys_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(outmemsys_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(outmemsys_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(outmemsys_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(outmemsys_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(outmemsys_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(outmemsys_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(outmemsys_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(outmemsys_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(outmemsys_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(outmemsys_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(outmemsys_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(outmemsys_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(outmemsys_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(outmemsys_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(outmemsys_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(outmemsys_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(outmemsys_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(outmemsys_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(outmemsys_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(outmemsys_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(outmemsys_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(outmemsys_io_tiles_uncached_0_grant_bits_data),
    .io_htif_uncached_acquire_ready(outmemsys_io_htif_uncached_acquire_ready),
    .io_htif_uncached_acquire_valid(outmemsys_io_htif_uncached_acquire_valid),
    .io_htif_uncached_acquire_bits_addr_block(outmemsys_io_htif_uncached_acquire_bits_addr_block),
    .io_htif_uncached_acquire_bits_client_xact_id(outmemsys_io_htif_uncached_acquire_bits_client_xact_id),
    .io_htif_uncached_acquire_bits_addr_beat(outmemsys_io_htif_uncached_acquire_bits_addr_beat),
    .io_htif_uncached_acquire_bits_is_builtin_type(outmemsys_io_htif_uncached_acquire_bits_is_builtin_type),
    .io_htif_uncached_acquire_bits_a_type(outmemsys_io_htif_uncached_acquire_bits_a_type),
    .io_htif_uncached_acquire_bits_union(outmemsys_io_htif_uncached_acquire_bits_union),
    .io_htif_uncached_acquire_bits_data(outmemsys_io_htif_uncached_acquire_bits_data),
    .io_htif_uncached_grant_ready(outmemsys_io_htif_uncached_grant_ready),
    .io_htif_uncached_grant_valid(outmemsys_io_htif_uncached_grant_valid),
    .io_htif_uncached_grant_bits_addr_beat(outmemsys_io_htif_uncached_grant_bits_addr_beat),
    .io_htif_uncached_grant_bits_client_xact_id(outmemsys_io_htif_uncached_grant_bits_client_xact_id),
    .io_htif_uncached_grant_bits_manager_xact_id(outmemsys_io_htif_uncached_grant_bits_manager_xact_id),
    .io_htif_uncached_grant_bits_is_builtin_type(outmemsys_io_htif_uncached_grant_bits_is_builtin_type),
    .io_htif_uncached_grant_bits_g_type(outmemsys_io_htif_uncached_grant_bits_g_type),
    .io_htif_uncached_grant_bits_data(outmemsys_io_htif_uncached_grant_bits_data),
    .io_incoherent_0(outmemsys_io_incoherent_0),
    .io_mem_axi_0_aw_ready(outmemsys_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(outmemsys_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(outmemsys_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(outmemsys_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(outmemsys_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(outmemsys_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(outmemsys_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(outmemsys_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(outmemsys_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(outmemsys_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(outmemsys_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(outmemsys_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(outmemsys_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(outmemsys_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(outmemsys_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(outmemsys_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(outmemsys_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(outmemsys_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(outmemsys_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(outmemsys_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(outmemsys_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(outmemsys_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(outmemsys_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(outmemsys_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(outmemsys_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(outmemsys_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(outmemsys_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(outmemsys_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(outmemsys_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(outmemsys_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(outmemsys_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(outmemsys_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(outmemsys_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(outmemsys_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(outmemsys_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(outmemsys_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(outmemsys_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(outmemsys_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(outmemsys_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(outmemsys_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(outmemsys_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(outmemsys_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(outmemsys_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(outmemsys_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(outmemsys_io_mem_axi_0_r_bits_user),
    .io_mmio_acquire_ready(outmemsys_io_mmio_acquire_ready),
    .io_mmio_acquire_valid(outmemsys_io_mmio_acquire_valid),
    .io_mmio_acquire_bits_addr_block(outmemsys_io_mmio_acquire_bits_addr_block),
    .io_mmio_acquire_bits_client_xact_id(outmemsys_io_mmio_acquire_bits_client_xact_id),
    .io_mmio_acquire_bits_addr_beat(outmemsys_io_mmio_acquire_bits_addr_beat),
    .io_mmio_acquire_bits_is_builtin_type(outmemsys_io_mmio_acquire_bits_is_builtin_type),
    .io_mmio_acquire_bits_a_type(outmemsys_io_mmio_acquire_bits_a_type),
    .io_mmio_acquire_bits_union(outmemsys_io_mmio_acquire_bits_union),
    .io_mmio_acquire_bits_data(outmemsys_io_mmio_acquire_bits_data),
    .io_mmio_grant_ready(outmemsys_io_mmio_grant_ready),
    .io_mmio_grant_valid(outmemsys_io_mmio_grant_valid),
    .io_mmio_grant_bits_addr_beat(outmemsys_io_mmio_grant_bits_addr_beat),
    .io_mmio_grant_bits_client_xact_id(outmemsys_io_mmio_grant_bits_client_xact_id),
    .io_mmio_grant_bits_manager_xact_id(outmemsys_io_mmio_grant_bits_manager_xact_id),
    .io_mmio_grant_bits_is_builtin_type(outmemsys_io_mmio_grant_bits_is_builtin_type),
    .io_mmio_grant_bits_g_type(outmemsys_io_mmio_grant_bits_g_type),
    .io_mmio_grant_bits_data(outmemsys_io_mmio_grant_bits_data)
  );
  SCRFile scrFile (
    .clk(scrFile_clk),
    .reset(scrFile_reset),
    .io_smi_req_ready(scrFile_io_smi_req_ready),
    .io_smi_req_valid(scrFile_io_smi_req_valid),
    .io_smi_req_bits_rw(scrFile_io_smi_req_bits_rw),
    .io_smi_req_bits_addr(scrFile_io_smi_req_bits_addr),
    .io_smi_req_bits_data(scrFile_io_smi_req_bits_data),
    .io_smi_resp_ready(scrFile_io_smi_resp_ready),
    .io_smi_resp_valid(scrFile_io_smi_resp_valid),
    .io_smi_resp_bits(scrFile_io_smi_resp_bits),
    .io_scr_rdata_0(scrFile_io_scr_rdata_0),
    .io_scr_rdata_1(scrFile_io_scr_rdata_1),
    .io_scr_rdata_2(scrFile_io_scr_rdata_2),
    .io_scr_rdata_3(scrFile_io_scr_rdata_3),
    .io_scr_rdata_4(scrFile_io_scr_rdata_4),
    .io_scr_rdata_5(scrFile_io_scr_rdata_5),
    .io_scr_rdata_6(scrFile_io_scr_rdata_6),
    .io_scr_rdata_7(scrFile_io_scr_rdata_7),
    .io_scr_rdata_8(scrFile_io_scr_rdata_8),
    .io_scr_rdata_9(scrFile_io_scr_rdata_9),
    .io_scr_rdata_10(scrFile_io_scr_rdata_10),
    .io_scr_rdata_11(scrFile_io_scr_rdata_11),
    .io_scr_rdata_12(scrFile_io_scr_rdata_12),
    .io_scr_rdata_13(scrFile_io_scr_rdata_13),
    .io_scr_rdata_14(scrFile_io_scr_rdata_14),
    .io_scr_rdata_15(scrFile_io_scr_rdata_15),
    .io_scr_rdata_16(scrFile_io_scr_rdata_16),
    .io_scr_rdata_17(scrFile_io_scr_rdata_17),
    .io_scr_rdata_18(scrFile_io_scr_rdata_18),
    .io_scr_rdata_19(scrFile_io_scr_rdata_19),
    .io_scr_rdata_20(scrFile_io_scr_rdata_20),
    .io_scr_rdata_21(scrFile_io_scr_rdata_21),
    .io_scr_rdata_22(scrFile_io_scr_rdata_22),
    .io_scr_rdata_23(scrFile_io_scr_rdata_23),
    .io_scr_rdata_24(scrFile_io_scr_rdata_24),
    .io_scr_rdata_25(scrFile_io_scr_rdata_25),
    .io_scr_rdata_26(scrFile_io_scr_rdata_26),
    .io_scr_rdata_27(scrFile_io_scr_rdata_27),
    .io_scr_rdata_28(scrFile_io_scr_rdata_28),
    .io_scr_rdata_29(scrFile_io_scr_rdata_29),
    .io_scr_rdata_30(scrFile_io_scr_rdata_30),
    .io_scr_rdata_31(scrFile_io_scr_rdata_31),
    .io_scr_rdata_32(scrFile_io_scr_rdata_32),
    .io_scr_rdata_33(scrFile_io_scr_rdata_33),
    .io_scr_rdata_34(scrFile_io_scr_rdata_34),
    .io_scr_rdata_35(scrFile_io_scr_rdata_35),
    .io_scr_rdata_36(scrFile_io_scr_rdata_36),
    .io_scr_rdata_37(scrFile_io_scr_rdata_37),
    .io_scr_rdata_38(scrFile_io_scr_rdata_38),
    .io_scr_rdata_39(scrFile_io_scr_rdata_39),
    .io_scr_rdata_40(scrFile_io_scr_rdata_40),
    .io_scr_rdata_41(scrFile_io_scr_rdata_41),
    .io_scr_rdata_42(scrFile_io_scr_rdata_42),
    .io_scr_rdata_43(scrFile_io_scr_rdata_43),
    .io_scr_rdata_44(scrFile_io_scr_rdata_44),
    .io_scr_rdata_45(scrFile_io_scr_rdata_45),
    .io_scr_rdata_46(scrFile_io_scr_rdata_46),
    .io_scr_rdata_47(scrFile_io_scr_rdata_47),
    .io_scr_rdata_48(scrFile_io_scr_rdata_48),
    .io_scr_rdata_49(scrFile_io_scr_rdata_49),
    .io_scr_rdata_50(scrFile_io_scr_rdata_50),
    .io_scr_rdata_51(scrFile_io_scr_rdata_51),
    .io_scr_rdata_52(scrFile_io_scr_rdata_52),
    .io_scr_rdata_53(scrFile_io_scr_rdata_53),
    .io_scr_rdata_54(scrFile_io_scr_rdata_54),
    .io_scr_rdata_55(scrFile_io_scr_rdata_55),
    .io_scr_rdata_56(scrFile_io_scr_rdata_56),
    .io_scr_rdata_57(scrFile_io_scr_rdata_57),
    .io_scr_rdata_58(scrFile_io_scr_rdata_58),
    .io_scr_rdata_59(scrFile_io_scr_rdata_59),
    .io_scr_rdata_60(scrFile_io_scr_rdata_60),
    .io_scr_rdata_61(scrFile_io_scr_rdata_61),
    .io_scr_rdata_62(scrFile_io_scr_rdata_62),
    .io_scr_rdata_63(scrFile_io_scr_rdata_63),
    .io_scr_wen(scrFile_io_scr_wen),
    .io_scr_waddr(scrFile_io_scr_waddr),
    .io_scr_wdata(scrFile_io_scr_wdata)
  );
  TileLinkRecursiveInterconnect TileLinkRecursiveInterconnect_8716 (
    .clk(TileLinkRecursiveInterconnect_8716_clk),
    .reset(TileLinkRecursiveInterconnect_8716_reset),
    .io_in_0_acquire_ready(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(TileLinkRecursiveInterconnect_8716_io_in_0_grant_ready),
    .io_in_0_grant_valid(TileLinkRecursiveInterconnect_8716_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_data),
    .io_out_0_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_ready),
    .io_out_0_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_valid),
    .io_out_0_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_block),
    .io_out_0_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_client_xact_id),
    .io_out_0_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_beat),
    .io_out_0_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_is_builtin_type),
    .io_out_0_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_a_type),
    .io_out_0_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_union),
    .io_out_0_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_data),
    .io_out_0_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_0_grant_ready),
    .io_out_0_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_0_grant_valid),
    .io_out_0_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_addr_beat),
    .io_out_0_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_client_xact_id),
    .io_out_0_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_manager_xact_id),
    .io_out_0_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_is_builtin_type),
    .io_out_0_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_g_type),
    .io_out_0_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_data),
    .io_out_1_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_ready),
    .io_out_1_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_valid),
    .io_out_1_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_block),
    .io_out_1_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_client_xact_id),
    .io_out_1_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_beat),
    .io_out_1_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_is_builtin_type),
    .io_out_1_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_a_type),
    .io_out_1_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_union),
    .io_out_1_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_data),
    .io_out_1_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_1_grant_ready),
    .io_out_1_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_1_grant_valid),
    .io_out_1_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_addr_beat),
    .io_out_1_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_client_xact_id),
    .io_out_1_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_manager_xact_id),
    .io_out_1_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_is_builtin_type),
    .io_out_1_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_g_type),
    .io_out_1_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_data),
    .io_out_2_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_ready),
    .io_out_2_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_valid),
    .io_out_2_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_block),
    .io_out_2_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_client_xact_id),
    .io_out_2_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_beat),
    .io_out_2_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_is_builtin_type),
    .io_out_2_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_a_type),
    .io_out_2_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_union),
    .io_out_2_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_data),
    .io_out_2_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_2_grant_ready),
    .io_out_2_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_2_grant_valid),
    .io_out_2_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_addr_beat),
    .io_out_2_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_client_xact_id),
    .io_out_2_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_manager_xact_id),
    .io_out_2_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_is_builtin_type),
    .io_out_2_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_g_type),
    .io_out_2_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_data),
    .io_out_3_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_ready),
    .io_out_3_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_valid),
    .io_out_3_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_block),
    .io_out_3_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_client_xact_id),
    .io_out_3_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_beat),
    .io_out_3_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_is_builtin_type),
    .io_out_3_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_a_type),
    .io_out_3_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_union),
    .io_out_3_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_data),
    .io_out_3_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_3_grant_ready),
    .io_out_3_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_3_grant_valid),
    .io_out_3_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_addr_beat),
    .io_out_3_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_client_xact_id),
    .io_out_3_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_manager_xact_id),
    .io_out_3_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_is_builtin_type),
    .io_out_3_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_g_type),
    .io_out_3_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_data),
    .io_out_4_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_ready),
    .io_out_4_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_valid),
    .io_out_4_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_block),
    .io_out_4_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_client_xact_id),
    .io_out_4_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_beat),
    .io_out_4_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_is_builtin_type),
    .io_out_4_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_a_type),
    .io_out_4_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_union),
    .io_out_4_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_data),
    .io_out_4_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_4_grant_ready),
    .io_out_4_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_4_grant_valid),
    .io_out_4_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_addr_beat),
    .io_out_4_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_client_xact_id),
    .io_out_4_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_manager_xact_id),
    .io_out_4_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_is_builtin_type),
    .io_out_4_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_g_type),
    .io_out_4_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_data),
    .io_out_5_acquire_ready(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_ready),
    .io_out_5_acquire_valid(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_valid),
    .io_out_5_acquire_bits_addr_block(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_block),
    .io_out_5_acquire_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_client_xact_id),
    .io_out_5_acquire_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_beat),
    .io_out_5_acquire_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_is_builtin_type),
    .io_out_5_acquire_bits_a_type(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_a_type),
    .io_out_5_acquire_bits_union(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_union),
    .io_out_5_acquire_bits_data(TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_data),
    .io_out_5_grant_ready(TileLinkRecursiveInterconnect_8716_io_out_5_grant_ready),
    .io_out_5_grant_valid(TileLinkRecursiveInterconnect_8716_io_out_5_grant_valid),
    .io_out_5_grant_bits_addr_beat(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_addr_beat),
    .io_out_5_grant_bits_client_xact_id(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_client_xact_id),
    .io_out_5_grant_bits_manager_xact_id(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_manager_xact_id),
    .io_out_5_grant_bits_is_builtin_type(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_is_builtin_type),
    .io_out_5_grant_bits_g_type(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_g_type),
    .io_out_5_grant_bits_data(TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_data)
  );
  RTC RTC_8717 (
    .clk(RTC_8717_clk),
    .reset(RTC_8717_reset),
    .io_tl_acquire_ready(RTC_8717_io_tl_acquire_ready),
    .io_tl_acquire_valid(RTC_8717_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(RTC_8717_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(RTC_8717_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(RTC_8717_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(RTC_8717_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(RTC_8717_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(RTC_8717_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(RTC_8717_io_tl_acquire_bits_data),
    .io_tl_grant_ready(RTC_8717_io_tl_grant_ready),
    .io_tl_grant_valid(RTC_8717_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(RTC_8717_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(RTC_8717_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(RTC_8717_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(RTC_8717_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(RTC_8717_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(RTC_8717_io_tl_grant_bits_data),
    .io_irqs_0(RTC_8717_io_irqs_0)
  );
  PLIC PLIC_8718 (
    .clk(PLIC_8718_clk),
    .reset(PLIC_8718_reset),
    .io_devices_0_valid(PLIC_8718_io_devices_0_valid),
    .io_devices_0_ready(PLIC_8718_io_devices_0_ready),
    .io_devices_0_complete(PLIC_8718_io_devices_0_complete),
    .io_devices_1_valid(PLIC_8718_io_devices_1_valid),
    .io_devices_1_ready(PLIC_8718_io_devices_1_ready),
    .io_devices_1_complete(PLIC_8718_io_devices_1_complete),
    .io_harts_0(PLIC_8718_io_harts_0),
    .io_harts_1(PLIC_8718_io_harts_1),
    .io_tl_acquire_ready(PLIC_8718_io_tl_acquire_ready),
    .io_tl_acquire_valid(PLIC_8718_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PLIC_8718_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PLIC_8718_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PLIC_8718_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PLIC_8718_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PLIC_8718_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PLIC_8718_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PLIC_8718_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PLIC_8718_io_tl_grant_ready),
    .io_tl_grant_valid(PLIC_8718_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PLIC_8718_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PLIC_8718_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PLIC_8718_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PLIC_8718_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PLIC_8718_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PLIC_8718_io_tl_grant_bits_data)
  );
  LevelGateway LevelGateway_8719 (
    .clk(LevelGateway_8719_clk),
    .reset(LevelGateway_8719_reset),
    .io_interrupt(LevelGateway_8719_io_interrupt),
    .io_plic_valid(LevelGateway_8719_io_plic_valid),
    .io_plic_ready(LevelGateway_8719_io_plic_ready),
    .io_plic_complete(LevelGateway_8719_io_plic_complete)
  );
  LevelGateway LevelGateway_51_8720 (
    .clk(LevelGateway_51_8720_clk),
    .reset(LevelGateway_51_8720_reset),
    .io_interrupt(LevelGateway_51_8720_io_interrupt),
    .io_plic_valid(LevelGateway_51_8720_io_plic_valid),
    .io_plic_ready(LevelGateway_51_8720_io_plic_ready),
    .io_plic_complete(LevelGateway_51_8720_io_plic_complete)
  );
  DebugModule DebugModule_8721 (
    .clk(DebugModule_8721_clk),
    .reset(DebugModule_8721_reset),
    .io_db_req_ready(DebugModule_8721_io_db_req_ready),
    .io_db_req_valid(DebugModule_8721_io_db_req_valid),
    .io_db_req_bits_addr(DebugModule_8721_io_db_req_bits_addr),
    .io_db_req_bits_op(DebugModule_8721_io_db_req_bits_op),
    .io_db_req_bits_data(DebugModule_8721_io_db_req_bits_data),
    .io_db_resp_ready(DebugModule_8721_io_db_resp_ready),
    .io_db_resp_valid(DebugModule_8721_io_db_resp_valid),
    .io_db_resp_bits_resp(DebugModule_8721_io_db_resp_bits_resp),
    .io_db_resp_bits_data(DebugModule_8721_io_db_resp_bits_data),
    .io_debugInterrupts_0(DebugModule_8721_io_debugInterrupts_0),
    .io_tl_acquire_ready(DebugModule_8721_io_tl_acquire_ready),
    .io_tl_acquire_valid(DebugModule_8721_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(DebugModule_8721_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(DebugModule_8721_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(DebugModule_8721_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(DebugModule_8721_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(DebugModule_8721_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(DebugModule_8721_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(DebugModule_8721_io_tl_acquire_bits_data),
    .io_tl_grant_ready(DebugModule_8721_io_tl_grant_ready),
    .io_tl_grant_valid(DebugModule_8721_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(DebugModule_8721_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(DebugModule_8721_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(DebugModule_8721_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(DebugModule_8721_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(DebugModule_8721_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(DebugModule_8721_io_tl_grant_bits_data),
    .io_ndreset(DebugModule_8721_io_ndreset),
    .io_fullreset(DebugModule_8721_io_fullreset)
  );
  PRCI PRCI_8722 (
    .clk(PRCI_8722_clk),
    .reset(PRCI_8722_reset),
    .io_interrupts_0_mtip(PRCI_8722_io_interrupts_0_mtip),
    .io_interrupts_0_meip(PRCI_8722_io_interrupts_0_meip),
    .io_interrupts_0_seip(PRCI_8722_io_interrupts_0_seip),
    .io_interrupts_0_debug(PRCI_8722_io_interrupts_0_debug),
    .io_tl_acquire_ready(PRCI_8722_io_tl_acquire_ready),
    .io_tl_acquire_valid(PRCI_8722_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(PRCI_8722_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(PRCI_8722_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(PRCI_8722_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(PRCI_8722_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(PRCI_8722_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(PRCI_8722_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(PRCI_8722_io_tl_acquire_bits_data),
    .io_tl_grant_ready(PRCI_8722_io_tl_grant_ready),
    .io_tl_grant_valid(PRCI_8722_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(PRCI_8722_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(PRCI_8722_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(PRCI_8722_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(PRCI_8722_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(PRCI_8722_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(PRCI_8722_io_tl_grant_bits_data),
    .io_tiles_0_reset(PRCI_8722_io_tiles_0_reset),
    .io_tiles_0_id(PRCI_8722_io_tiles_0_id),
    .io_tiles_0_interrupts_mtip(PRCI_8722_io_tiles_0_interrupts_mtip),
    .io_tiles_0_interrupts_meip(PRCI_8722_io_tiles_0_interrupts_meip),
    .io_tiles_0_interrupts_seip(PRCI_8722_io_tiles_0_interrupts_seip),
    .io_tiles_0_interrupts_debug(PRCI_8722_io_tiles_0_interrupts_debug),
    .io_tiles_0_interrupts_msip(PRCI_8722_io_tiles_0_interrupts_msip)
  );
  ROMSlave ROMSlave_8728 (
    .clk(ROMSlave_8728_clk),
    .reset(ROMSlave_8728_reset),
    .io_acquire_ready(ROMSlave_8728_io_acquire_ready),
    .io_acquire_valid(ROMSlave_8728_io_acquire_valid),
    .io_acquire_bits_addr_block(ROMSlave_8728_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(ROMSlave_8728_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(ROMSlave_8728_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(ROMSlave_8728_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(ROMSlave_8728_io_acquire_bits_a_type),
    .io_acquire_bits_union(ROMSlave_8728_io_acquire_bits_union),
    .io_acquire_bits_data(ROMSlave_8728_io_acquire_bits_data),
    .io_grant_ready(ROMSlave_8728_io_grant_ready),
    .io_grant_valid(ROMSlave_8728_io_grant_valid),
    .io_grant_bits_addr_beat(ROMSlave_8728_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(ROMSlave_8728_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(ROMSlave_8728_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(ROMSlave_8728_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(ROMSlave_8728_io_grant_bits_g_type),
    .io_grant_bits_data(ROMSlave_8728_io_grant_bits_data)
  );
  NastiErrorSlave NastiErrorSlave_8729 (
    .clk(NastiErrorSlave_8729_clk),
    .reset(NastiErrorSlave_8729_reset),
    .io_aw_ready(NastiErrorSlave_8729_io_aw_ready),
    .io_aw_valid(NastiErrorSlave_8729_io_aw_valid),
    .io_aw_bits_addr(NastiErrorSlave_8729_io_aw_bits_addr),
    .io_aw_bits_len(NastiErrorSlave_8729_io_aw_bits_len),
    .io_aw_bits_size(NastiErrorSlave_8729_io_aw_bits_size),
    .io_aw_bits_burst(NastiErrorSlave_8729_io_aw_bits_burst),
    .io_aw_bits_lock(NastiErrorSlave_8729_io_aw_bits_lock),
    .io_aw_bits_cache(NastiErrorSlave_8729_io_aw_bits_cache),
    .io_aw_bits_prot(NastiErrorSlave_8729_io_aw_bits_prot),
    .io_aw_bits_qos(NastiErrorSlave_8729_io_aw_bits_qos),
    .io_aw_bits_region(NastiErrorSlave_8729_io_aw_bits_region),
    .io_aw_bits_id(NastiErrorSlave_8729_io_aw_bits_id),
    .io_aw_bits_user(NastiErrorSlave_8729_io_aw_bits_user),
    .io_w_ready(NastiErrorSlave_8729_io_w_ready),
    .io_w_valid(NastiErrorSlave_8729_io_w_valid),
    .io_w_bits_data(NastiErrorSlave_8729_io_w_bits_data),
    .io_w_bits_last(NastiErrorSlave_8729_io_w_bits_last),
    .io_w_bits_id(NastiErrorSlave_8729_io_w_bits_id),
    .io_w_bits_strb(NastiErrorSlave_8729_io_w_bits_strb),
    .io_w_bits_user(NastiErrorSlave_8729_io_w_bits_user),
    .io_b_ready(NastiErrorSlave_8729_io_b_ready),
    .io_b_valid(NastiErrorSlave_8729_io_b_valid),
    .io_b_bits_resp(NastiErrorSlave_8729_io_b_bits_resp),
    .io_b_bits_id(NastiErrorSlave_8729_io_b_bits_id),
    .io_b_bits_user(NastiErrorSlave_8729_io_b_bits_user),
    .io_ar_ready(NastiErrorSlave_8729_io_ar_ready),
    .io_ar_valid(NastiErrorSlave_8729_io_ar_valid),
    .io_ar_bits_addr(NastiErrorSlave_8729_io_ar_bits_addr),
    .io_ar_bits_len(NastiErrorSlave_8729_io_ar_bits_len),
    .io_ar_bits_size(NastiErrorSlave_8729_io_ar_bits_size),
    .io_ar_bits_burst(NastiErrorSlave_8729_io_ar_bits_burst),
    .io_ar_bits_lock(NastiErrorSlave_8729_io_ar_bits_lock),
    .io_ar_bits_cache(NastiErrorSlave_8729_io_ar_bits_cache),
    .io_ar_bits_prot(NastiErrorSlave_8729_io_ar_bits_prot),
    .io_ar_bits_qos(NastiErrorSlave_8729_io_ar_bits_qos),
    .io_ar_bits_region(NastiErrorSlave_8729_io_ar_bits_region),
    .io_ar_bits_id(NastiErrorSlave_8729_io_ar_bits_id),
    .io_ar_bits_user(NastiErrorSlave_8729_io_ar_bits_user),
    .io_r_ready(NastiErrorSlave_8729_io_r_ready),
    .io_r_valid(NastiErrorSlave_8729_io_r_valid),
    .io_r_bits_resp(NastiErrorSlave_8729_io_r_bits_resp),
    .io_r_bits_data(NastiErrorSlave_8729_io_r_bits_data),
    .io_r_bits_last(NastiErrorSlave_8729_io_r_bits_last),
    .io_r_bits_id(NastiErrorSlave_8729_io_r_bits_id),
    .io_r_bits_user(NastiErrorSlave_8729_io_r_bits_user)
  );
  NastiIOTileLinkIOConverter_56 NastiIOTileLinkIOConverter_56_8730 (
    .clk(NastiIOTileLinkIOConverter_56_8730_clk),
    .reset(NastiIOTileLinkIOConverter_56_8730_reset),
    .io_tl_acquire_ready(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_ready),
    .io_tl_acquire_valid(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_valid),
    .io_tl_acquire_bits_addr_block(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_block),
    .io_tl_acquire_bits_client_xact_id(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_client_xact_id),
    .io_tl_acquire_bits_addr_beat(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_beat),
    .io_tl_acquire_bits_is_builtin_type(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_is_builtin_type),
    .io_tl_acquire_bits_a_type(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_a_type),
    .io_tl_acquire_bits_union(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_union),
    .io_tl_acquire_bits_data(NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_data),
    .io_tl_grant_ready(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_ready),
    .io_tl_grant_valid(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_valid),
    .io_tl_grant_bits_addr_beat(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_addr_beat),
    .io_tl_grant_bits_client_xact_id(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_client_xact_id),
    .io_tl_grant_bits_manager_xact_id(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_manager_xact_id),
    .io_tl_grant_bits_is_builtin_type(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_is_builtin_type),
    .io_tl_grant_bits_g_type(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_g_type),
    .io_tl_grant_bits_data(NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_data),
    .io_nasti_aw_ready(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_ready),
    .io_nasti_aw_valid(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_addr),
    .io_nasti_aw_bits_len(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_len),
    .io_nasti_aw_bits_size(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_size),
    .io_nasti_aw_bits_burst(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_burst),
    .io_nasti_aw_bits_lock(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_lock),
    .io_nasti_aw_bits_cache(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_cache),
    .io_nasti_aw_bits_prot(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_prot),
    .io_nasti_aw_bits_qos(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_qos),
    .io_nasti_aw_bits_region(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_region),
    .io_nasti_aw_bits_id(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_id),
    .io_nasti_aw_bits_user(NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_user),
    .io_nasti_w_ready(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_ready),
    .io_nasti_w_valid(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_valid),
    .io_nasti_w_bits_data(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_last),
    .io_nasti_w_bits_id(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_id),
    .io_nasti_w_bits_strb(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_strb),
    .io_nasti_w_bits_user(NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_user),
    .io_nasti_b_ready(NastiIOTileLinkIOConverter_56_8730_io_nasti_b_ready),
    .io_nasti_b_valid(NastiIOTileLinkIOConverter_56_8730_io_nasti_b_valid),
    .io_nasti_b_bits_resp(NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_resp),
    .io_nasti_b_bits_id(NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_id),
    .io_nasti_b_bits_user(NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_user),
    .io_nasti_ar_ready(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_ready),
    .io_nasti_ar_valid(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_addr),
    .io_nasti_ar_bits_len(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_len),
    .io_nasti_ar_bits_size(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_size),
    .io_nasti_ar_bits_burst(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_burst),
    .io_nasti_ar_bits_lock(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_lock),
    .io_nasti_ar_bits_cache(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_cache),
    .io_nasti_ar_bits_prot(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_prot),
    .io_nasti_ar_bits_qos(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_qos),
    .io_nasti_ar_bits_region(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_region),
    .io_nasti_ar_bits_id(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_id),
    .io_nasti_ar_bits_user(NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_user),
    .io_nasti_r_ready(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_ready),
    .io_nasti_r_valid(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_valid),
    .io_nasti_r_bits_resp(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_resp),
    .io_nasti_r_bits_data(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_last),
    .io_nasti_r_bits_id(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_id),
    .io_nasti_r_bits_user(NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_user)
  );
  Queue_39 Queue_61_8743 (
    .clk(Queue_61_8743_clk),
    .reset(Queue_61_8743_reset),
    .io_enq_ready(Queue_61_8743_io_enq_ready),
    .io_enq_valid(Queue_61_8743_io_enq_valid),
    .io_enq_bits_addr(Queue_61_8743_io_enq_bits_addr),
    .io_enq_bits_len(Queue_61_8743_io_enq_bits_len),
    .io_enq_bits_size(Queue_61_8743_io_enq_bits_size),
    .io_enq_bits_burst(Queue_61_8743_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_61_8743_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_61_8743_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_61_8743_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_61_8743_io_enq_bits_qos),
    .io_enq_bits_region(Queue_61_8743_io_enq_bits_region),
    .io_enq_bits_id(Queue_61_8743_io_enq_bits_id),
    .io_enq_bits_user(Queue_61_8743_io_enq_bits_user),
    .io_deq_ready(Queue_61_8743_io_deq_ready),
    .io_deq_valid(Queue_61_8743_io_deq_valid),
    .io_deq_bits_addr(Queue_61_8743_io_deq_bits_addr),
    .io_deq_bits_len(Queue_61_8743_io_deq_bits_len),
    .io_deq_bits_size(Queue_61_8743_io_deq_bits_size),
    .io_deq_bits_burst(Queue_61_8743_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_61_8743_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_61_8743_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_61_8743_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_61_8743_io_deq_bits_qos),
    .io_deq_bits_region(Queue_61_8743_io_deq_bits_region),
    .io_deq_bits_id(Queue_61_8743_io_deq_bits_id),
    .io_deq_bits_user(Queue_61_8743_io_deq_bits_user),
    .io_count(Queue_61_8743_io_count)
  );
  Queue_39 Queue_62_8756 (
    .clk(Queue_62_8756_clk),
    .reset(Queue_62_8756_reset),
    .io_enq_ready(Queue_62_8756_io_enq_ready),
    .io_enq_valid(Queue_62_8756_io_enq_valid),
    .io_enq_bits_addr(Queue_62_8756_io_enq_bits_addr),
    .io_enq_bits_len(Queue_62_8756_io_enq_bits_len),
    .io_enq_bits_size(Queue_62_8756_io_enq_bits_size),
    .io_enq_bits_burst(Queue_62_8756_io_enq_bits_burst),
    .io_enq_bits_lock(Queue_62_8756_io_enq_bits_lock),
    .io_enq_bits_cache(Queue_62_8756_io_enq_bits_cache),
    .io_enq_bits_prot(Queue_62_8756_io_enq_bits_prot),
    .io_enq_bits_qos(Queue_62_8756_io_enq_bits_qos),
    .io_enq_bits_region(Queue_62_8756_io_enq_bits_region),
    .io_enq_bits_id(Queue_62_8756_io_enq_bits_id),
    .io_enq_bits_user(Queue_62_8756_io_enq_bits_user),
    .io_deq_ready(Queue_62_8756_io_deq_ready),
    .io_deq_valid(Queue_62_8756_io_deq_valid),
    .io_deq_bits_addr(Queue_62_8756_io_deq_bits_addr),
    .io_deq_bits_len(Queue_62_8756_io_deq_bits_len),
    .io_deq_bits_size(Queue_62_8756_io_deq_bits_size),
    .io_deq_bits_burst(Queue_62_8756_io_deq_bits_burst),
    .io_deq_bits_lock(Queue_62_8756_io_deq_bits_lock),
    .io_deq_bits_cache(Queue_62_8756_io_deq_bits_cache),
    .io_deq_bits_prot(Queue_62_8756_io_deq_bits_prot),
    .io_deq_bits_qos(Queue_62_8756_io_deq_bits_qos),
    .io_deq_bits_region(Queue_62_8756_io_deq_bits_region),
    .io_deq_bits_id(Queue_62_8756_io_deq_bits_id),
    .io_deq_bits_user(Queue_62_8756_io_deq_bits_user),
    .io_count(Queue_62_8756_io_count)
  );
  Queue_41 Queue_63_8763 (
    .clk(Queue_63_8763_clk),
    .reset(Queue_63_8763_reset),
    .io_enq_ready(Queue_63_8763_io_enq_ready),
    .io_enq_valid(Queue_63_8763_io_enq_valid),
    .io_enq_bits_data(Queue_63_8763_io_enq_bits_data),
    .io_enq_bits_last(Queue_63_8763_io_enq_bits_last),
    .io_enq_bits_id(Queue_63_8763_io_enq_bits_id),
    .io_enq_bits_strb(Queue_63_8763_io_enq_bits_strb),
    .io_enq_bits_user(Queue_63_8763_io_enq_bits_user),
    .io_deq_ready(Queue_63_8763_io_deq_ready),
    .io_deq_valid(Queue_63_8763_io_deq_valid),
    .io_deq_bits_data(Queue_63_8763_io_deq_bits_data),
    .io_deq_bits_last(Queue_63_8763_io_deq_bits_last),
    .io_deq_bits_id(Queue_63_8763_io_deq_bits_id),
    .io_deq_bits_strb(Queue_63_8763_io_deq_bits_strb),
    .io_deq_bits_user(Queue_63_8763_io_deq_bits_user),
    .io_count(Queue_63_8763_io_count)
  );
  Queue_42 Queue_64_8770 (
    .clk(Queue_64_8770_clk),
    .reset(Queue_64_8770_reset),
    .io_enq_ready(Queue_64_8770_io_enq_ready),
    .io_enq_valid(Queue_64_8770_io_enq_valid),
    .io_enq_bits_resp(Queue_64_8770_io_enq_bits_resp),
    .io_enq_bits_data(Queue_64_8770_io_enq_bits_data),
    .io_enq_bits_last(Queue_64_8770_io_enq_bits_last),
    .io_enq_bits_id(Queue_64_8770_io_enq_bits_id),
    .io_enq_bits_user(Queue_64_8770_io_enq_bits_user),
    .io_deq_ready(Queue_64_8770_io_deq_ready),
    .io_deq_valid(Queue_64_8770_io_deq_valid),
    .io_deq_bits_resp(Queue_64_8770_io_deq_bits_resp),
    .io_deq_bits_data(Queue_64_8770_io_deq_bits_data),
    .io_deq_bits_last(Queue_64_8770_io_deq_bits_last),
    .io_deq_bits_id(Queue_64_8770_io_deq_bits_id),
    .io_deq_bits_user(Queue_64_8770_io_deq_bits_user),
    .io_count(Queue_64_8770_io_count)
  );
  Queue_43 Queue_65_8775 (
    .clk(Queue_65_8775_clk),
    .reset(Queue_65_8775_reset),
    .io_enq_ready(Queue_65_8775_io_enq_ready),
    .io_enq_valid(Queue_65_8775_io_enq_valid),
    .io_enq_bits_resp(Queue_65_8775_io_enq_bits_resp),
    .io_enq_bits_id(Queue_65_8775_io_enq_bits_id),
    .io_enq_bits_user(Queue_65_8775_io_enq_bits_user),
    .io_deq_ready(Queue_65_8775_io_deq_ready),
    .io_deq_valid(Queue_65_8775_io_deq_valid),
    .io_deq_bits_resp(Queue_65_8775_io_deq_bits_resp),
    .io_deq_bits_id(Queue_65_8775_io_deq_bits_id),
    .io_deq_bits_user(Queue_65_8775_io_deq_bits_user),
    .io_count(Queue_65_8775_io_count)
  );
  assign io_host_clk = htif_io_host_clk;
  assign io_host_clk_edge = htif_io_host_clk_edge;
  assign io_host_in_ready = htif_io_host_in_ready;
  assign io_host_out_valid = htif_io_host_out_valid;
  assign io_host_out_bits = htif_io_host_out_bits;
  assign io_mem_axi_0_aw_valid = outmemsys_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = outmemsys_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = outmemsys_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = outmemsys_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = outmemsys_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = outmemsys_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = outmemsys_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = outmemsys_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = outmemsys_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = outmemsys_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = outmemsys_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = outmemsys_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = outmemsys_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = outmemsys_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = outmemsys_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = outmemsys_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = outmemsys_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = outmemsys_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = outmemsys_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = outmemsys_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = outmemsys_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = outmemsys_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = outmemsys_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = outmemsys_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = outmemsys_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = outmemsys_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = outmemsys_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = outmemsys_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = outmemsys_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = outmemsys_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = outmemsys_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = outmemsys_io_mem_axi_0_r_ready;
  assign io_tiles_cached_0_acquire_ready = outmemsys_io_tiles_cached_0_acquire_ready;
  assign io_tiles_cached_0_probe_valid = outmemsys_io_tiles_cached_0_probe_valid;
  assign io_tiles_cached_0_probe_bits_addr_block = outmemsys_io_tiles_cached_0_probe_bits_addr_block;
  assign io_tiles_cached_0_probe_bits_p_type = outmemsys_io_tiles_cached_0_probe_bits_p_type;
  assign io_tiles_cached_0_release_ready = outmemsys_io_tiles_cached_0_release_ready;
  assign io_tiles_cached_0_grant_valid = outmemsys_io_tiles_cached_0_grant_valid;
  assign io_tiles_cached_0_grant_bits_addr_beat = outmemsys_io_tiles_cached_0_grant_bits_addr_beat;
  assign io_tiles_cached_0_grant_bits_client_xact_id = outmemsys_io_tiles_cached_0_grant_bits_client_xact_id;
  assign io_tiles_cached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign io_tiles_cached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign io_tiles_cached_0_grant_bits_g_type = outmemsys_io_tiles_cached_0_grant_bits_g_type;
  assign io_tiles_cached_0_grant_bits_data = outmemsys_io_tiles_cached_0_grant_bits_data;
  assign io_tiles_cached_0_grant_bits_manager_id = outmemsys_io_tiles_cached_0_grant_bits_manager_id;
  assign io_tiles_cached_0_finish_ready = outmemsys_io_tiles_cached_0_finish_ready;
  assign io_tiles_uncached_0_acquire_ready = outmemsys_io_tiles_uncached_0_acquire_ready;
  assign io_tiles_uncached_0_grant_valid = outmemsys_io_tiles_uncached_0_grant_valid;
  assign io_tiles_uncached_0_grant_bits_addr_beat = outmemsys_io_tiles_uncached_0_grant_bits_addr_beat;
  assign io_tiles_uncached_0_grant_bits_client_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign io_tiles_uncached_0_grant_bits_manager_xact_id = outmemsys_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign io_tiles_uncached_0_grant_bits_is_builtin_type = outmemsys_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign io_tiles_uncached_0_grant_bits_g_type = outmemsys_io_tiles_uncached_0_grant_bits_g_type;
  assign io_tiles_uncached_0_grant_bits_data = outmemsys_io_tiles_uncached_0_grant_bits_data;
  assign io_prci_0_reset = T_8727;
  assign io_prci_0_id = PRCI_8722_io_tiles_0_id;
  assign io_prci_0_interrupts_mtip = PRCI_8722_io_tiles_0_interrupts_mtip;
  assign io_prci_0_interrupts_meip = PRCI_8722_io_tiles_0_interrupts_meip;
  assign io_prci_0_interrupts_seip = PRCI_8722_io_tiles_0_interrupts_seip;
  assign io_prci_0_interrupts_debug = PRCI_8722_io_tiles_0_interrupts_debug;
  assign io_prci_0_interrupts_msip = PRCI_8722_io_tiles_0_interrupts_msip;
  assign io_debugBus_req_ready = DebugModule_8721_io_db_req_ready;
  assign io_debugBus_resp_valid = DebugModule_8721_io_db_resp_valid;
  assign io_debugBus_resp_bits_resp = DebugModule_8721_io_db_resp_bits_resp;
  assign io_debugBus_resp_bits_data = DebugModule_8721_io_db_resp_bits_data;
  assign htif_clk = clk;
  assign htif_reset = reset;
  assign htif_io_host_in_valid = io_host_in_valid;
  assign htif_io_host_in_bits = io_host_in_bits;
  assign htif_io_host_out_ready = io_host_out_ready;
  assign htif_io_cpu_0_csr_req_ready = GEN_0;
  assign htif_io_cpu_0_csr_resp_valid = 1'h0;
  assign htif_io_cpu_0_csr_resp_bits = GEN_1;
  assign htif_io_mem_acquire_ready = outmemsys_io_htif_uncached_acquire_ready;
  assign htif_io_mem_grant_valid = outmemsys_io_htif_uncached_grant_valid;
  assign htif_io_mem_grant_bits_addr_beat = outmemsys_io_htif_uncached_grant_bits_addr_beat;
  assign htif_io_mem_grant_bits_client_xact_id = outmemsys_io_htif_uncached_grant_bits_client_xact_id;
  assign htif_io_mem_grant_bits_manager_xact_id = outmemsys_io_htif_uncached_grant_bits_manager_xact_id;
  assign htif_io_mem_grant_bits_is_builtin_type = outmemsys_io_htif_uncached_grant_bits_is_builtin_type;
  assign htif_io_mem_grant_bits_g_type = outmemsys_io_htif_uncached_grant_bits_g_type;
  assign htif_io_mem_grant_bits_data = outmemsys_io_htif_uncached_grant_bits_data;
  assign htif_io_scr_req_ready = scrFile_io_smi_req_ready;
  assign htif_io_scr_resp_valid = scrFile_io_smi_resp_valid;
  assign htif_io_scr_resp_bits = scrFile_io_smi_resp_bits;
  assign outmemsys_clk = clk;
  assign outmemsys_reset = reset;
  assign outmemsys_io_tiles_cached_0_acquire_valid = io_tiles_cached_0_acquire_valid;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_block = io_tiles_cached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_acquire_bits_client_xact_id = io_tiles_cached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_acquire_bits_addr_beat = io_tiles_cached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_acquire_bits_is_builtin_type = io_tiles_cached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_a_type = io_tiles_cached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_cached_0_acquire_bits_union = io_tiles_cached_0_acquire_bits_union;
  assign outmemsys_io_tiles_cached_0_acquire_bits_data = io_tiles_cached_0_acquire_bits_data;
  assign outmemsys_io_tiles_cached_0_probe_ready = io_tiles_cached_0_probe_ready;
  assign outmemsys_io_tiles_cached_0_release_valid = io_tiles_cached_0_release_valid;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_beat = io_tiles_cached_0_release_bits_addr_beat;
  assign outmemsys_io_tiles_cached_0_release_bits_addr_block = io_tiles_cached_0_release_bits_addr_block;
  assign outmemsys_io_tiles_cached_0_release_bits_client_xact_id = io_tiles_cached_0_release_bits_client_xact_id;
  assign outmemsys_io_tiles_cached_0_release_bits_voluntary = io_tiles_cached_0_release_bits_voluntary;
  assign outmemsys_io_tiles_cached_0_release_bits_r_type = io_tiles_cached_0_release_bits_r_type;
  assign outmemsys_io_tiles_cached_0_release_bits_data = io_tiles_cached_0_release_bits_data;
  assign outmemsys_io_tiles_cached_0_grant_ready = io_tiles_cached_0_grant_ready;
  assign outmemsys_io_tiles_cached_0_finish_valid = io_tiles_cached_0_finish_valid;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_xact_id = io_tiles_cached_0_finish_bits_manager_xact_id;
  assign outmemsys_io_tiles_cached_0_finish_bits_manager_id = io_tiles_cached_0_finish_bits_manager_id;
  assign outmemsys_io_tiles_uncached_0_acquire_valid = io_tiles_uncached_0_acquire_valid;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_block = io_tiles_uncached_0_acquire_bits_addr_block;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_client_xact_id = io_tiles_uncached_0_acquire_bits_client_xact_id;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_addr_beat = io_tiles_uncached_0_acquire_bits_addr_beat;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_is_builtin_type = io_tiles_uncached_0_acquire_bits_is_builtin_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_a_type = io_tiles_uncached_0_acquire_bits_a_type;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_union = io_tiles_uncached_0_acquire_bits_union;
  assign outmemsys_io_tiles_uncached_0_acquire_bits_data = io_tiles_uncached_0_acquire_bits_data;
  assign outmemsys_io_tiles_uncached_0_grant_ready = io_tiles_uncached_0_grant_ready;
  assign outmemsys_io_htif_uncached_acquire_valid = htif_io_mem_acquire_valid;
  assign outmemsys_io_htif_uncached_acquire_bits_addr_block = htif_io_mem_acquire_bits_addr_block;
  assign outmemsys_io_htif_uncached_acquire_bits_client_xact_id = htif_io_mem_acquire_bits_client_xact_id;
  assign outmemsys_io_htif_uncached_acquire_bits_addr_beat = htif_io_mem_acquire_bits_addr_beat;
  assign outmemsys_io_htif_uncached_acquire_bits_is_builtin_type = htif_io_mem_acquire_bits_is_builtin_type;
  assign outmemsys_io_htif_uncached_acquire_bits_a_type = htif_io_mem_acquire_bits_a_type;
  assign outmemsys_io_htif_uncached_acquire_bits_union = htif_io_mem_acquire_bits_union;
  assign outmemsys_io_htif_uncached_acquire_bits_data = htif_io_mem_acquire_bits_data;
  assign outmemsys_io_htif_uncached_grant_ready = htif_io_mem_grant_ready;
  assign outmemsys_io_incoherent_0 = htif_io_cpu_0_reset;
  assign outmemsys_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign outmemsys_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign outmemsys_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign outmemsys_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign outmemsys_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign outmemsys_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign outmemsys_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign outmemsys_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign outmemsys_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign outmemsys_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign outmemsys_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign outmemsys_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign outmemsys_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign outmemsys_io_mmio_acquire_ready = TileLinkRecursiveInterconnect_8716_io_in_0_acquire_ready;
  assign outmemsys_io_mmio_grant_valid = TileLinkRecursiveInterconnect_8716_io_in_0_grant_valid;
  assign outmemsys_io_mmio_grant_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_addr_beat;
  assign outmemsys_io_mmio_grant_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_client_xact_id;
  assign outmemsys_io_mmio_grant_bits_manager_xact_id = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_manager_xact_id;
  assign outmemsys_io_mmio_grant_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_is_builtin_type;
  assign outmemsys_io_mmio_grant_bits_g_type = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_g_type;
  assign outmemsys_io_mmio_grant_bits_data = TileLinkRecursiveInterconnect_8716_io_in_0_grant_bits_data;
  assign scrFile_clk = clk;
  assign scrFile_reset = reset;
  assign scrFile_io_smi_req_valid = htif_io_scr_req_valid;
  assign scrFile_io_smi_req_bits_rw = htif_io_scr_req_bits_rw;
  assign scrFile_io_smi_req_bits_addr = htif_io_scr_req_bits_addr;
  assign scrFile_io_smi_req_bits_data = htif_io_scr_req_bits_data;
  assign scrFile_io_smi_resp_ready = htif_io_scr_resp_ready;
  assign scrFile_io_scr_rdata_0 = GEN_2;
  assign scrFile_io_scr_rdata_1 = GEN_3;
  assign scrFile_io_scr_rdata_2 = GEN_4;
  assign scrFile_io_scr_rdata_3 = GEN_5;
  assign scrFile_io_scr_rdata_4 = GEN_6;
  assign scrFile_io_scr_rdata_5 = GEN_7;
  assign scrFile_io_scr_rdata_6 = GEN_8;
  assign scrFile_io_scr_rdata_7 = GEN_9;
  assign scrFile_io_scr_rdata_8 = GEN_10;
  assign scrFile_io_scr_rdata_9 = GEN_11;
  assign scrFile_io_scr_rdata_10 = GEN_12;
  assign scrFile_io_scr_rdata_11 = GEN_13;
  assign scrFile_io_scr_rdata_12 = GEN_14;
  assign scrFile_io_scr_rdata_13 = GEN_15;
  assign scrFile_io_scr_rdata_14 = GEN_16;
  assign scrFile_io_scr_rdata_15 = GEN_17;
  assign scrFile_io_scr_rdata_16 = GEN_18;
  assign scrFile_io_scr_rdata_17 = GEN_19;
  assign scrFile_io_scr_rdata_18 = GEN_20;
  assign scrFile_io_scr_rdata_19 = GEN_21;
  assign scrFile_io_scr_rdata_20 = GEN_22;
  assign scrFile_io_scr_rdata_21 = GEN_23;
  assign scrFile_io_scr_rdata_22 = GEN_24;
  assign scrFile_io_scr_rdata_23 = GEN_25;
  assign scrFile_io_scr_rdata_24 = GEN_26;
  assign scrFile_io_scr_rdata_25 = GEN_27;
  assign scrFile_io_scr_rdata_26 = GEN_28;
  assign scrFile_io_scr_rdata_27 = GEN_29;
  assign scrFile_io_scr_rdata_28 = GEN_30;
  assign scrFile_io_scr_rdata_29 = GEN_31;
  assign scrFile_io_scr_rdata_30 = GEN_32;
  assign scrFile_io_scr_rdata_31 = GEN_33;
  assign scrFile_io_scr_rdata_32 = GEN_34;
  assign scrFile_io_scr_rdata_33 = GEN_35;
  assign scrFile_io_scr_rdata_34 = GEN_36;
  assign scrFile_io_scr_rdata_35 = GEN_37;
  assign scrFile_io_scr_rdata_36 = GEN_38;
  assign scrFile_io_scr_rdata_37 = GEN_39;
  assign scrFile_io_scr_rdata_38 = GEN_40;
  assign scrFile_io_scr_rdata_39 = GEN_41;
  assign scrFile_io_scr_rdata_40 = GEN_42;
  assign scrFile_io_scr_rdata_41 = GEN_43;
  assign scrFile_io_scr_rdata_42 = GEN_44;
  assign scrFile_io_scr_rdata_43 = GEN_45;
  assign scrFile_io_scr_rdata_44 = GEN_46;
  assign scrFile_io_scr_rdata_45 = GEN_47;
  assign scrFile_io_scr_rdata_46 = GEN_48;
  assign scrFile_io_scr_rdata_47 = GEN_49;
  assign scrFile_io_scr_rdata_48 = GEN_50;
  assign scrFile_io_scr_rdata_49 = GEN_51;
  assign scrFile_io_scr_rdata_50 = GEN_52;
  assign scrFile_io_scr_rdata_51 = GEN_53;
  assign scrFile_io_scr_rdata_52 = GEN_54;
  assign scrFile_io_scr_rdata_53 = GEN_55;
  assign scrFile_io_scr_rdata_54 = GEN_56;
  assign scrFile_io_scr_rdata_55 = GEN_57;
  assign scrFile_io_scr_rdata_56 = GEN_58;
  assign scrFile_io_scr_rdata_57 = GEN_59;
  assign scrFile_io_scr_rdata_58 = GEN_60;
  assign scrFile_io_scr_rdata_59 = GEN_61;
  assign scrFile_io_scr_rdata_60 = GEN_62;
  assign scrFile_io_scr_rdata_61 = GEN_63;
  assign scrFile_io_scr_rdata_62 = GEN_64;
  assign scrFile_io_scr_rdata_63 = GEN_65;
  assign TileLinkRecursiveInterconnect_8716_clk = clk;
  assign TileLinkRecursiveInterconnect_8716_reset = reset;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_valid = outmemsys_io_mmio_acquire_valid;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_block = outmemsys_io_mmio_acquire_bits_addr_block;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_client_xact_id = outmemsys_io_mmio_acquire_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_addr_beat = outmemsys_io_mmio_acquire_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_is_builtin_type = outmemsys_io_mmio_acquire_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_a_type = outmemsys_io_mmio_acquire_bits_a_type;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_union = outmemsys_io_mmio_acquire_bits_union;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_acquire_bits_data = outmemsys_io_mmio_acquire_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_in_0_grant_ready = outmemsys_io_mmio_grant_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_acquire_ready = DebugModule_8721_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_valid = DebugModule_8721_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_addr_beat = DebugModule_8721_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_client_xact_id = DebugModule_8721_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_manager_xact_id = DebugModule_8721_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_is_builtin_type = DebugModule_8721_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_g_type = DebugModule_8721_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_0_grant_bits_data = DebugModule_8721_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_acquire_ready = ROMSlave_8728_io_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_valid = ROMSlave_8728_io_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_addr_beat = ROMSlave_8728_io_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_client_xact_id = ROMSlave_8728_io_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_manager_xact_id = ROMSlave_8728_io_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_is_builtin_type = ROMSlave_8728_io_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_g_type = ROMSlave_8728_io_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_1_grant_bits_data = ROMSlave_8728_io_grant_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_acquire_ready = RTC_8717_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_valid = RTC_8717_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_addr_beat = RTC_8717_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_client_xact_id = RTC_8717_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_manager_xact_id = RTC_8717_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_is_builtin_type = RTC_8717_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_g_type = RTC_8717_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_2_grant_bits_data = RTC_8717_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_acquire_ready = PLIC_8718_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_valid = PLIC_8718_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_addr_beat = PLIC_8718_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_client_xact_id = PLIC_8718_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_manager_xact_id = PLIC_8718_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_is_builtin_type = PLIC_8718_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_g_type = PLIC_8718_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_3_grant_bits_data = PLIC_8718_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_acquire_ready = PRCI_8722_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_valid = PRCI_8722_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_addr_beat = PRCI_8722_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_client_xact_id = PRCI_8722_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_manager_xact_id = PRCI_8722_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_is_builtin_type = PRCI_8722_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_g_type = PRCI_8722_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_4_grant_bits_data = PRCI_8722_io_tl_grant_bits_data;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_acquire_ready = NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_ready;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_valid = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_valid;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_addr_beat = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_addr_beat;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_client_xact_id = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_client_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_manager_xact_id = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_manager_xact_id;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_is_builtin_type = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_is_builtin_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_g_type = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_g_type;
  assign TileLinkRecursiveInterconnect_8716_io_out_5_grant_bits_data = NastiIOTileLinkIOConverter_56_8730_io_tl_grant_bits_data;
  assign RTC_8717_clk = clk;
  assign RTC_8717_reset = reset;
  assign RTC_8717_io_tl_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_valid;
  assign RTC_8717_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_block;
  assign RTC_8717_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_client_xact_id;
  assign RTC_8717_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_addr_beat;
  assign RTC_8717_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_is_builtin_type;
  assign RTC_8717_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_a_type;
  assign RTC_8717_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_union;
  assign RTC_8717_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_2_acquire_bits_data;
  assign RTC_8717_io_tl_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_2_grant_ready;
  assign PLIC_8718_clk = clk;
  assign PLIC_8718_reset = reset;
  assign PLIC_8718_io_devices_0_valid = LevelGateway_8719_io_plic_valid;
  assign PLIC_8718_io_devices_1_valid = LevelGateway_51_8720_io_plic_valid;
  assign PLIC_8718_io_tl_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_valid;
  assign PLIC_8718_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_block;
  assign PLIC_8718_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_client_xact_id;
  assign PLIC_8718_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_addr_beat;
  assign PLIC_8718_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_is_builtin_type;
  assign PLIC_8718_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_a_type;
  assign PLIC_8718_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_union;
  assign PLIC_8718_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_3_acquire_bits_data;
  assign PLIC_8718_io_tl_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_3_grant_ready;
  assign LevelGateway_8719_clk = clk;
  assign LevelGateway_8719_reset = reset;
  assign LevelGateway_8719_io_interrupt = io_interrupts_0;
  assign LevelGateway_8719_io_plic_ready = PLIC_8718_io_devices_0_ready;
  assign LevelGateway_8719_io_plic_complete = PLIC_8718_io_devices_0_complete;
  assign LevelGateway_51_8720_clk = clk;
  assign LevelGateway_51_8720_reset = reset;
  assign LevelGateway_51_8720_io_interrupt = io_interrupts_1;
  assign LevelGateway_51_8720_io_plic_ready = PLIC_8718_io_devices_1_ready;
  assign LevelGateway_51_8720_io_plic_complete = PLIC_8718_io_devices_1_complete;
  assign DebugModule_8721_clk = clk;
  assign DebugModule_8721_reset = reset;
  assign DebugModule_8721_io_db_req_valid = io_debugBus_req_valid;
  assign DebugModule_8721_io_db_req_bits_addr = io_debugBus_req_bits_addr;
  assign DebugModule_8721_io_db_req_bits_op = io_debugBus_req_bits_op;
  assign DebugModule_8721_io_db_req_bits_data = io_debugBus_req_bits_data;
  assign DebugModule_8721_io_db_resp_ready = io_debugBus_resp_ready;
  assign DebugModule_8721_io_tl_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_valid;
  assign DebugModule_8721_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_block;
  assign DebugModule_8721_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_client_xact_id;
  assign DebugModule_8721_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_addr_beat;
  assign DebugModule_8721_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_is_builtin_type;
  assign DebugModule_8721_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_a_type;
  assign DebugModule_8721_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_union;
  assign DebugModule_8721_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_0_acquire_bits_data;
  assign DebugModule_8721_io_tl_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_0_grant_ready;
  assign PRCI_8722_clk = clk;
  assign PRCI_8722_reset = reset;
  assign PRCI_8722_io_interrupts_0_mtip = RTC_8717_io_irqs_0;
  assign PRCI_8722_io_interrupts_0_meip = PLIC_8718_io_harts_0;
  assign PRCI_8722_io_interrupts_0_seip = PLIC_8718_io_harts_1;
  assign PRCI_8722_io_interrupts_0_debug = DebugModule_8721_io_debugInterrupts_0;
  assign PRCI_8722_io_tl_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_valid;
  assign PRCI_8722_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_block;
  assign PRCI_8722_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_client_xact_id;
  assign PRCI_8722_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_addr_beat;
  assign PRCI_8722_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_is_builtin_type;
  assign PRCI_8722_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_a_type;
  assign PRCI_8722_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_union;
  assign PRCI_8722_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_4_acquire_bits_data;
  assign PRCI_8722_io_tl_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_4_grant_ready;
  assign T_8727 = reset | T_8726;
  assign ROMSlave_8728_clk = clk;
  assign ROMSlave_8728_reset = reset;
  assign ROMSlave_8728_io_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_valid;
  assign ROMSlave_8728_io_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_block;
  assign ROMSlave_8728_io_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_client_xact_id;
  assign ROMSlave_8728_io_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_addr_beat;
  assign ROMSlave_8728_io_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_is_builtin_type;
  assign ROMSlave_8728_io_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_a_type;
  assign ROMSlave_8728_io_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_union;
  assign ROMSlave_8728_io_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_1_acquire_bits_data;
  assign ROMSlave_8728_io_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_1_grant_ready;
  assign NastiErrorSlave_8729_clk = clk;
  assign NastiErrorSlave_8729_reset = reset;
  assign NastiErrorSlave_8729_io_aw_valid = Queue_62_8756_io_deq_valid;
  assign NastiErrorSlave_8729_io_aw_bits_addr = Queue_62_8756_io_deq_bits_addr;
  assign NastiErrorSlave_8729_io_aw_bits_len = Queue_62_8756_io_deq_bits_len;
  assign NastiErrorSlave_8729_io_aw_bits_size = Queue_62_8756_io_deq_bits_size;
  assign NastiErrorSlave_8729_io_aw_bits_burst = Queue_62_8756_io_deq_bits_burst;
  assign NastiErrorSlave_8729_io_aw_bits_lock = Queue_62_8756_io_deq_bits_lock;
  assign NastiErrorSlave_8729_io_aw_bits_cache = Queue_62_8756_io_deq_bits_cache;
  assign NastiErrorSlave_8729_io_aw_bits_prot = Queue_62_8756_io_deq_bits_prot;
  assign NastiErrorSlave_8729_io_aw_bits_qos = Queue_62_8756_io_deq_bits_qos;
  assign NastiErrorSlave_8729_io_aw_bits_region = Queue_62_8756_io_deq_bits_region;
  assign NastiErrorSlave_8729_io_aw_bits_id = Queue_62_8756_io_deq_bits_id;
  assign NastiErrorSlave_8729_io_aw_bits_user = Queue_62_8756_io_deq_bits_user;
  assign NastiErrorSlave_8729_io_w_valid = Queue_63_8763_io_deq_valid;
  assign NastiErrorSlave_8729_io_w_bits_data = Queue_63_8763_io_deq_bits_data;
  assign NastiErrorSlave_8729_io_w_bits_last = Queue_63_8763_io_deq_bits_last;
  assign NastiErrorSlave_8729_io_w_bits_id = Queue_63_8763_io_deq_bits_id;
  assign NastiErrorSlave_8729_io_w_bits_strb = Queue_63_8763_io_deq_bits_strb;
  assign NastiErrorSlave_8729_io_w_bits_user = Queue_63_8763_io_deq_bits_user;
  assign NastiErrorSlave_8729_io_b_ready = Queue_65_8775_io_enq_ready;
  assign NastiErrorSlave_8729_io_ar_valid = Queue_61_8743_io_deq_valid;
  assign NastiErrorSlave_8729_io_ar_bits_addr = Queue_61_8743_io_deq_bits_addr;
  assign NastiErrorSlave_8729_io_ar_bits_len = Queue_61_8743_io_deq_bits_len;
  assign NastiErrorSlave_8729_io_ar_bits_size = Queue_61_8743_io_deq_bits_size;
  assign NastiErrorSlave_8729_io_ar_bits_burst = Queue_61_8743_io_deq_bits_burst;
  assign NastiErrorSlave_8729_io_ar_bits_lock = Queue_61_8743_io_deq_bits_lock;
  assign NastiErrorSlave_8729_io_ar_bits_cache = Queue_61_8743_io_deq_bits_cache;
  assign NastiErrorSlave_8729_io_ar_bits_prot = Queue_61_8743_io_deq_bits_prot;
  assign NastiErrorSlave_8729_io_ar_bits_qos = Queue_61_8743_io_deq_bits_qos;
  assign NastiErrorSlave_8729_io_ar_bits_region = Queue_61_8743_io_deq_bits_region;
  assign NastiErrorSlave_8729_io_ar_bits_id = Queue_61_8743_io_deq_bits_id;
  assign NastiErrorSlave_8729_io_ar_bits_user = Queue_61_8743_io_deq_bits_user;
  assign NastiErrorSlave_8729_io_r_ready = Queue_64_8770_io_enq_ready;
  assign NastiIOTileLinkIOConverter_56_8730_clk = clk;
  assign NastiIOTileLinkIOConverter_56_8730_reset = reset;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_valid = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_valid;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_block = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_block;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_client_xact_id = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_client_xact_id;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_addr_beat = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_addr_beat;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_is_builtin_type = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_is_builtin_type;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_a_type = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_a_type;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_union = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_union;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_acquire_bits_data = TileLinkRecursiveInterconnect_8716_io_out_5_acquire_bits_data;
  assign NastiIOTileLinkIOConverter_56_8730_io_tl_grant_ready = TileLinkRecursiveInterconnect_8716_io_out_5_grant_ready;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_ready = Queue_62_8756_io_enq_ready;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_w_ready = Queue_63_8763_io_enq_ready;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_b_valid = Queue_65_8775_io_deq_valid;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_resp = Queue_65_8775_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_id = Queue_65_8775_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_b_bits_user = Queue_65_8775_io_deq_bits_user;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_ready = Queue_61_8743_io_enq_ready;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_valid = Queue_64_8770_io_deq_valid;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_resp = Queue_64_8770_io_deq_bits_resp;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_data = Queue_64_8770_io_deq_bits_data;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_last = Queue_64_8770_io_deq_bits_last;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_id = Queue_64_8770_io_deq_bits_id;
  assign NastiIOTileLinkIOConverter_56_8730_io_nasti_r_bits_user = Queue_64_8770_io_deq_bits_user;
  assign Queue_61_8743_clk = clk;
  assign Queue_61_8743_reset = reset;
  assign Queue_61_8743_io_enq_valid = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_valid;
  assign Queue_61_8743_io_enq_bits_addr = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_addr;
  assign Queue_61_8743_io_enq_bits_len = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_len;
  assign Queue_61_8743_io_enq_bits_size = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_size;
  assign Queue_61_8743_io_enq_bits_burst = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_burst;
  assign Queue_61_8743_io_enq_bits_lock = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_lock;
  assign Queue_61_8743_io_enq_bits_cache = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_cache;
  assign Queue_61_8743_io_enq_bits_prot = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_prot;
  assign Queue_61_8743_io_enq_bits_qos = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_qos;
  assign Queue_61_8743_io_enq_bits_region = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_region;
  assign Queue_61_8743_io_enq_bits_id = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_id;
  assign Queue_61_8743_io_enq_bits_user = NastiIOTileLinkIOConverter_56_8730_io_nasti_ar_bits_user;
  assign Queue_61_8743_io_deq_ready = NastiErrorSlave_8729_io_ar_ready;
  assign Queue_62_8756_clk = clk;
  assign Queue_62_8756_reset = reset;
  assign Queue_62_8756_io_enq_valid = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_valid;
  assign Queue_62_8756_io_enq_bits_addr = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_addr;
  assign Queue_62_8756_io_enq_bits_len = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_len;
  assign Queue_62_8756_io_enq_bits_size = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_size;
  assign Queue_62_8756_io_enq_bits_burst = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_burst;
  assign Queue_62_8756_io_enq_bits_lock = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_lock;
  assign Queue_62_8756_io_enq_bits_cache = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_cache;
  assign Queue_62_8756_io_enq_bits_prot = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_prot;
  assign Queue_62_8756_io_enq_bits_qos = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_qos;
  assign Queue_62_8756_io_enq_bits_region = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_region;
  assign Queue_62_8756_io_enq_bits_id = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_id;
  assign Queue_62_8756_io_enq_bits_user = NastiIOTileLinkIOConverter_56_8730_io_nasti_aw_bits_user;
  assign Queue_62_8756_io_deq_ready = NastiErrorSlave_8729_io_aw_ready;
  assign Queue_63_8763_clk = clk;
  assign Queue_63_8763_reset = reset;
  assign Queue_63_8763_io_enq_valid = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_valid;
  assign Queue_63_8763_io_enq_bits_data = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_data;
  assign Queue_63_8763_io_enq_bits_last = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_last;
  assign Queue_63_8763_io_enq_bits_id = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_id;
  assign Queue_63_8763_io_enq_bits_strb = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_strb;
  assign Queue_63_8763_io_enq_bits_user = NastiIOTileLinkIOConverter_56_8730_io_nasti_w_bits_user;
  assign Queue_63_8763_io_deq_ready = NastiErrorSlave_8729_io_w_ready;
  assign Queue_64_8770_clk = clk;
  assign Queue_64_8770_reset = reset;
  assign Queue_64_8770_io_enq_valid = NastiErrorSlave_8729_io_r_valid;
  assign Queue_64_8770_io_enq_bits_resp = NastiErrorSlave_8729_io_r_bits_resp;
  assign Queue_64_8770_io_enq_bits_data = NastiErrorSlave_8729_io_r_bits_data;
  assign Queue_64_8770_io_enq_bits_last = NastiErrorSlave_8729_io_r_bits_last;
  assign Queue_64_8770_io_enq_bits_id = NastiErrorSlave_8729_io_r_bits_id;
  assign Queue_64_8770_io_enq_bits_user = NastiErrorSlave_8729_io_r_bits_user;
  assign Queue_64_8770_io_deq_ready = NastiIOTileLinkIOConverter_56_8730_io_nasti_r_ready;
  assign Queue_65_8775_clk = clk;
  assign Queue_65_8775_reset = reset;
  assign Queue_65_8775_io_enq_valid = NastiErrorSlave_8729_io_b_valid;
  assign Queue_65_8775_io_enq_bits_resp = NastiErrorSlave_8729_io_b_bits_resp;
  assign Queue_65_8775_io_enq_bits_id = NastiErrorSlave_8729_io_b_bits_id;
  assign Queue_65_8775_io_enq_bits_user = NastiErrorSlave_8729_io_b_bits_user;
  assign Queue_65_8775_io_deq_ready = NastiIOTileLinkIOConverter_56_8730_io_nasti_b_ready;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_66 = {1{$random}};
  T_8725 = GEN_66[0:0];
  GEN_67 = {1{$random}};
  T_8726 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  GEN_0 = GEN_68[0:0];
  GEN_69 = {2{$random}};
  GEN_1 = GEN_69[63:0];
  GEN_70 = {2{$random}};
  GEN_2 = GEN_70[63:0];
  GEN_71 = {2{$random}};
  GEN_3 = GEN_71[63:0];
  GEN_72 = {2{$random}};
  GEN_4 = GEN_72[63:0];
  GEN_73 = {2{$random}};
  GEN_5 = GEN_73[63:0];
  GEN_74 = {2{$random}};
  GEN_6 = GEN_74[63:0];
  GEN_75 = {2{$random}};
  GEN_7 = GEN_75[63:0];
  GEN_76 = {2{$random}};
  GEN_8 = GEN_76[63:0];
  GEN_77 = {2{$random}};
  GEN_9 = GEN_77[63:0];
  GEN_78 = {2{$random}};
  GEN_10 = GEN_78[63:0];
  GEN_79 = {2{$random}};
  GEN_11 = GEN_79[63:0];
  GEN_80 = {2{$random}};
  GEN_12 = GEN_80[63:0];
  GEN_81 = {2{$random}};
  GEN_13 = GEN_81[63:0];
  GEN_82 = {2{$random}};
  GEN_14 = GEN_82[63:0];
  GEN_83 = {2{$random}};
  GEN_15 = GEN_83[63:0];
  GEN_84 = {2{$random}};
  GEN_16 = GEN_84[63:0];
  GEN_85 = {2{$random}};
  GEN_17 = GEN_85[63:0];
  GEN_86 = {2{$random}};
  GEN_18 = GEN_86[63:0];
  GEN_87 = {2{$random}};
  GEN_19 = GEN_87[63:0];
  GEN_88 = {2{$random}};
  GEN_20 = GEN_88[63:0];
  GEN_89 = {2{$random}};
  GEN_21 = GEN_89[63:0];
  GEN_90 = {2{$random}};
  GEN_22 = GEN_90[63:0];
  GEN_91 = {2{$random}};
  GEN_23 = GEN_91[63:0];
  GEN_92 = {2{$random}};
  GEN_24 = GEN_92[63:0];
  GEN_93 = {2{$random}};
  GEN_25 = GEN_93[63:0];
  GEN_94 = {2{$random}};
  GEN_26 = GEN_94[63:0];
  GEN_95 = {2{$random}};
  GEN_27 = GEN_95[63:0];
  GEN_96 = {2{$random}};
  GEN_28 = GEN_96[63:0];
  GEN_97 = {2{$random}};
  GEN_29 = GEN_97[63:0];
  GEN_98 = {2{$random}};
  GEN_30 = GEN_98[63:0];
  GEN_99 = {2{$random}};
  GEN_31 = GEN_99[63:0];
  GEN_100 = {2{$random}};
  GEN_32 = GEN_100[63:0];
  GEN_101 = {2{$random}};
  GEN_33 = GEN_101[63:0];
  GEN_102 = {2{$random}};
  GEN_34 = GEN_102[63:0];
  GEN_103 = {2{$random}};
  GEN_35 = GEN_103[63:0];
  GEN_104 = {2{$random}};
  GEN_36 = GEN_104[63:0];
  GEN_105 = {2{$random}};
  GEN_37 = GEN_105[63:0];
  GEN_106 = {2{$random}};
  GEN_38 = GEN_106[63:0];
  GEN_107 = {2{$random}};
  GEN_39 = GEN_107[63:0];
  GEN_108 = {2{$random}};
  GEN_40 = GEN_108[63:0];
  GEN_109 = {2{$random}};
  GEN_41 = GEN_109[63:0];
  GEN_110 = {2{$random}};
  GEN_42 = GEN_110[63:0];
  GEN_111 = {2{$random}};
  GEN_43 = GEN_111[63:0];
  GEN_112 = {2{$random}};
  GEN_44 = GEN_112[63:0];
  GEN_113 = {2{$random}};
  GEN_45 = GEN_113[63:0];
  GEN_114 = {2{$random}};
  GEN_46 = GEN_114[63:0];
  GEN_115 = {2{$random}};
  GEN_47 = GEN_115[63:0];
  GEN_116 = {2{$random}};
  GEN_48 = GEN_116[63:0];
  GEN_117 = {2{$random}};
  GEN_49 = GEN_117[63:0];
  GEN_118 = {2{$random}};
  GEN_50 = GEN_118[63:0];
  GEN_119 = {2{$random}};
  GEN_51 = GEN_119[63:0];
  GEN_120 = {2{$random}};
  GEN_52 = GEN_120[63:0];
  GEN_121 = {2{$random}};
  GEN_53 = GEN_121[63:0];
  GEN_122 = {2{$random}};
  GEN_54 = GEN_122[63:0];
  GEN_123 = {2{$random}};
  GEN_55 = GEN_123[63:0];
  GEN_124 = {2{$random}};
  GEN_56 = GEN_124[63:0];
  GEN_125 = {2{$random}};
  GEN_57 = GEN_125[63:0];
  GEN_126 = {2{$random}};
  GEN_58 = GEN_126[63:0];
  GEN_127 = {2{$random}};
  GEN_59 = GEN_127[63:0];
  GEN_128 = {2{$random}};
  GEN_60 = GEN_128[63:0];
  GEN_129 = {2{$random}};
  GEN_61 = GEN_129[63:0];
  GEN_130 = {2{$random}};
  GEN_62 = GEN_130[63:0];
  GEN_131 = {2{$random}};
  GEN_63 = GEN_131[63:0];
  GEN_132 = {2{$random}};
  GEN_64 = GEN_132[63:0];
  GEN_133 = {2{$random}};
  GEN_65 = GEN_133[63:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_8725 <= 1'h1;
    end else begin
      T_8725 <= htif_io_cpu_0_reset;
    end
    if(reset) begin
      T_8726 <= 1'h1;
    end else begin
      T_8726 <= T_8725;
    end
  end
endmodule
module CSRFile(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_msip,
  input  [11:0] io_rw_addr,
  input  [2:0] io_rw_cmd,
  output [63:0] io_rw_rdata,
  input  [63:0] io_rw_wdata,
  output  io_csr_stall,
  output  io_csr_xcpt,
  output  io_eret,
  output [1:0] io_prv,
  output  io_status_debug,
  output [1:0] io_status_prv,
  output  io_status_sd,
  output [30:0] io_status_zero3,
  output  io_status_sd_rv32,
  output [1:0] io_status_zero2,
  output [4:0] io_status_vm,
  output [4:0] io_status_zero1,
  output  io_status_pum,
  output  io_status_mprv,
  output [1:0] io_status_xs,
  output [1:0] io_status_fs,
  output [1:0] io_status_mpp,
  output [1:0] io_status_hpp,
  output  io_status_spp,
  output  io_status_mpie,
  output  io_status_hpie,
  output  io_status_spie,
  output  io_status_upie,
  output  io_status_mie,
  output  io_status_hie,
  output  io_status_sie,
  output  io_status_uie,
  output [31:0] io_ptbr,
  output [39:0] io_evec,
  input   io_exception,
  input   io_retire,
  input   io_uarch_counters_0,
  input   io_uarch_counters_1,
  input   io_uarch_counters_2,
  input   io_uarch_counters_3,
  input   io_uarch_counters_4,
  input   io_uarch_counters_5,
  input   io_uarch_counters_6,
  input   io_uarch_counters_7,
  input   io_uarch_counters_8,
  input   io_uarch_counters_9,
  input   io_uarch_counters_10,
  input   io_uarch_counters_11,
  input   io_uarch_counters_12,
  input   io_uarch_counters_13,
  input   io_uarch_counters_14,
  input   io_uarch_counters_15,
  input  [63:0] io_cause,
  input  [39:0] io_pc,
  input  [39:0] io_badaddr,
  output  io_fatc,
  output [63:0] io_time,
  output [2:0] io_fcsr_rm,
  input   io_fcsr_flags_valid,
  input  [4:0] io_fcsr_flags_bits,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  output  io_rocc_status_debug,
  output [1:0] io_rocc_status_prv,
  output  io_rocc_status_sd,
  output [30:0] io_rocc_status_zero3,
  output  io_rocc_status_sd_rv32,
  output [1:0] io_rocc_status_zero2,
  output [4:0] io_rocc_status_vm,
  output [4:0] io_rocc_status_zero1,
  output  io_rocc_status_pum,
  output  io_rocc_status_mprv,
  output [1:0] io_rocc_status_xs,
  output [1:0] io_rocc_status_fs,
  output [1:0] io_rocc_status_mpp,
  output [1:0] io_rocc_status_hpp,
  output  io_rocc_status_spp,
  output  io_rocc_status_mpie,
  output  io_rocc_status_hpie,
  output  io_rocc_status_spie,
  output  io_rocc_status_upie,
  output  io_rocc_status_mie,
  output  io_rocc_status_hie,
  output  io_rocc_status_sie,
  output  io_rocc_status_uie,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [63:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id,
  output  io_interrupt,
  output [63:0] io_interrupt_cause,
  output [3:0] io_bp_0_control_tdrtype,
  output [4:0] io_bp_0_control_bpamaskmax,
  output [35:0] io_bp_0_control_reserved,
  output [7:0] io_bp_0_control_bpaction,
  output [3:0] io_bp_0_control_bpmatch,
  output  io_bp_0_control_m,
  output  io_bp_0_control_h,
  output  io_bp_0_control_s,
  output  io_bp_0_control_u,
  output  io_bp_0_control_r,
  output  io_bp_0_control_w,
  output  io_bp_0_control_x,
  output [38:0] io_bp_0_address
);
  wire  T_4951_debug;
  wire [1:0] T_4951_prv;
  wire  T_4951_sd;
  wire [30:0] T_4951_zero3;
  wire  T_4951_sd_rv32;
  wire [1:0] T_4951_zero2;
  wire [4:0] T_4951_vm;
  wire [4:0] T_4951_zero1;
  wire  T_4951_pum;
  wire  T_4951_mprv;
  wire [1:0] T_4951_xs;
  wire [1:0] T_4951_fs;
  wire [1:0] T_4951_mpp;
  wire [1:0] T_4951_hpp;
  wire  T_4951_spp;
  wire  T_4951_mpie;
  wire  T_4951_hpie;
  wire  T_4951_spie;
  wire  T_4951_upie;
  wire  T_4951_mie;
  wire  T_4951_hie;
  wire  T_4951_sie;
  wire  T_4951_uie;
  wire [66:0] T_4976;
  wire  T_4977;
  wire  T_4978;
  wire  T_4979;
  wire  T_4980;
  wire  T_4981;
  wire  T_4982;
  wire  T_4983;
  wire  T_4984;
  wire  T_4985;
  wire [1:0] T_4986;
  wire [1:0] T_4987;
  wire [1:0] T_4988;
  wire [1:0] T_4989;
  wire  T_4990;
  wire  T_4991;
  wire [4:0] T_4992;
  wire [4:0] T_4993;
  wire [1:0] T_4994;
  wire  T_4995;
  wire [30:0] T_4996;
  wire  T_4997;
  wire [1:0] T_4998;
  wire  T_4999;
  wire  reset_mstatus_debug;
  wire [1:0] reset_mstatus_prv;
  wire  reset_mstatus_sd;
  wire [30:0] reset_mstatus_zero3;
  wire  reset_mstatus_sd_rv32;
  wire [1:0] reset_mstatus_zero2;
  wire [4:0] reset_mstatus_vm;
  wire [4:0] reset_mstatus_zero1;
  wire  reset_mstatus_pum;
  wire  reset_mstatus_mprv;
  wire [1:0] reset_mstatus_xs;
  wire [1:0] reset_mstatus_fs;
  wire [1:0] reset_mstatus_mpp;
  wire [1:0] reset_mstatus_hpp;
  wire  reset_mstatus_spp;
  wire  reset_mstatus_mpie;
  wire  reset_mstatus_hpie;
  wire  reset_mstatus_spie;
  wire  reset_mstatus_upie;
  wire  reset_mstatus_mie;
  wire  reset_mstatus_hie;
  wire  reset_mstatus_sie;
  wire  reset_mstatus_uie;
  reg  reg_mstatus_debug;
  reg [31:0] GEN_237;
  reg [1:0] reg_mstatus_prv;
  reg [31:0] GEN_238;
  reg  reg_mstatus_sd;
  reg [31:0] GEN_239;
  reg [30:0] reg_mstatus_zero3;
  reg [31:0] GEN_240;
  reg  reg_mstatus_sd_rv32;
  reg [31:0] GEN_241;
  reg [1:0] reg_mstatus_zero2;
  reg [31:0] GEN_242;
  reg [4:0] reg_mstatus_vm;
  reg [31:0] GEN_243;
  reg [4:0] reg_mstatus_zero1;
  reg [31:0] GEN_244;
  reg  reg_mstatus_pum;
  reg [31:0] GEN_245;
  reg  reg_mstatus_mprv;
  reg [31:0] GEN_246;
  reg [1:0] reg_mstatus_xs;
  reg [31:0] GEN_247;
  reg [1:0] reg_mstatus_fs;
  reg [31:0] GEN_253;
  reg [1:0] reg_mstatus_mpp;
  reg [31:0] GEN_254;
  reg [1:0] reg_mstatus_hpp;
  reg [31:0] GEN_255;
  reg  reg_mstatus_spp;
  reg [31:0] GEN_256;
  reg  reg_mstatus_mpie;
  reg [31:0] GEN_257;
  reg  reg_mstatus_hpie;
  reg [31:0] GEN_258;
  reg  reg_mstatus_spie;
  reg [31:0] GEN_259;
  reg  reg_mstatus_upie;
  reg [31:0] GEN_260;
  reg  reg_mstatus_mie;
  reg [31:0] GEN_261;
  reg  reg_mstatus_hie;
  reg [31:0] GEN_262;
  reg  reg_mstatus_sie;
  reg [31:0] GEN_263;
  reg  reg_mstatus_uie;
  reg [31:0] GEN_264;
  wire [1:0] T_5085_xdebugver;
  wire  T_5085_ndreset;
  wire  T_5085_fullreset;
  wire [11:0] T_5085_hwbpcount;
  wire  T_5085_ebreakm;
  wire  T_5085_ebreakh;
  wire  T_5085_ebreaks;
  wire  T_5085_ebreaku;
  wire  T_5085_zero2;
  wire  T_5085_stopcycle;
  wire  T_5085_stoptime;
  wire [2:0] T_5085_cause;
  wire  T_5085_debugint;
  wire  T_5085_zero1;
  wire  T_5085_halt;
  wire  T_5085_step;
  wire [1:0] T_5085_prv;
  wire [31:0] T_5104;
  wire [1:0] T_5105;
  wire  T_5106;
  wire  T_5107;
  wire  T_5108;
  wire  T_5109;
  wire [2:0] T_5110;
  wire  T_5111;
  wire  T_5112;
  wire  T_5113;
  wire  T_5114;
  wire  T_5115;
  wire  T_5116;
  wire  T_5117;
  wire [11:0] T_5118;
  wire  T_5119;
  wire  T_5120;
  wire [1:0] T_5121;
  wire [1:0] reset_dcsr_xdebugver;
  wire  reset_dcsr_ndreset;
  wire  reset_dcsr_fullreset;
  wire [11:0] reset_dcsr_hwbpcount;
  wire  reset_dcsr_ebreakm;
  wire  reset_dcsr_ebreakh;
  wire  reset_dcsr_ebreaks;
  wire  reset_dcsr_ebreaku;
  wire  reset_dcsr_zero2;
  wire  reset_dcsr_stopcycle;
  wire  reset_dcsr_stoptime;
  wire [2:0] reset_dcsr_cause;
  wire  reset_dcsr_debugint;
  wire  reset_dcsr_zero1;
  wire  reset_dcsr_halt;
  wire  reset_dcsr_step;
  wire [1:0] reset_dcsr_prv;
  reg [1:0] reg_dcsr_xdebugver;
  reg [31:0] GEN_265;
  reg  reg_dcsr_ndreset;
  reg [31:0] GEN_277;
  reg  reg_dcsr_fullreset;
  reg [31:0] GEN_278;
  reg [11:0] reg_dcsr_hwbpcount;
  reg [31:0] GEN_279;
  reg  reg_dcsr_ebreakm;
  reg [31:0] GEN_280;
  reg  reg_dcsr_ebreakh;
  reg [31:0] GEN_281;
  reg  reg_dcsr_ebreaks;
  reg [31:0] GEN_282;
  reg  reg_dcsr_ebreaku;
  reg [31:0] GEN_283;
  reg  reg_dcsr_zero2;
  reg [31:0] GEN_284;
  reg  reg_dcsr_stopcycle;
  reg [31:0] GEN_286;
  reg  reg_dcsr_stoptime;
  reg [31:0] GEN_288;
  reg [2:0] reg_dcsr_cause;
  reg [31:0] GEN_289;
  reg  reg_dcsr_debugint;
  reg [31:0] GEN_290;
  reg  reg_dcsr_zero1;
  reg [31:0] GEN_292;
  reg  reg_dcsr_halt;
  reg [31:0] GEN_294;
  reg  reg_dcsr_step;
  reg [31:0] GEN_296;
  reg [1:0] reg_dcsr_prv;
  reg [31:0] GEN_298;
  wire  T_5187_rocc;
  wire  T_5187_meip;
  wire  T_5187_heip;
  wire  T_5187_seip;
  wire  T_5187_ueip;
  wire  T_5187_mtip;
  wire  T_5187_htip;
  wire  T_5187_stip;
  wire  T_5187_utip;
  wire  T_5187_msip;
  wire  T_5187_hsip;
  wire  T_5187_ssip;
  wire  T_5187_usip;
  wire [12:0] T_5202;
  wire  T_5203;
  wire  T_5204;
  wire  T_5205;
  wire  T_5206;
  wire  T_5207;
  wire  T_5208;
  wire  T_5209;
  wire  T_5210;
  wire  T_5211;
  wire  T_5212;
  wire  T_5213;
  wire  T_5214;
  wire  T_5215;
  wire  T_5216_rocc;
  wire  T_5216_meip;
  wire  T_5216_heip;
  wire  T_5216_seip;
  wire  T_5216_ueip;
  wire  T_5216_mtip;
  wire  T_5216_htip;
  wire  T_5216_stip;
  wire  T_5216_utip;
  wire  T_5216_msip;
  wire  T_5216_hsip;
  wire  T_5216_ssip;
  wire  T_5216_usip;
  wire  T_5237_rocc;
  wire  T_5237_meip;
  wire  T_5237_heip;
  wire  T_5237_seip;
  wire  T_5237_ueip;
  wire  T_5237_mtip;
  wire  T_5237_htip;
  wire  T_5237_stip;
  wire  T_5237_utip;
  wire  T_5237_msip;
  wire  T_5237_hsip;
  wire  T_5237_ssip;
  wire  T_5237_usip;
  wire [1:0] T_5254;
  wire [2:0] T_5255;
  wire [1:0] T_5256;
  wire [2:0] T_5257;
  wire [5:0] T_5258;
  wire [1:0] T_5259;
  wire [2:0] T_5260;
  wire [1:0] T_5261;
  wire [1:0] T_5262;
  wire [3:0] T_5263;
  wire [6:0] T_5264;
  wire [12:0] supported_interrupts;
  wire [1:0] T_5265;
  wire [2:0] T_5266;
  wire [1:0] T_5267;
  wire [2:0] T_5268;
  wire [5:0] T_5269;
  wire [1:0] T_5270;
  wire [2:0] T_5271;
  wire [1:0] T_5272;
  wire [1:0] T_5273;
  wire [3:0] T_5274;
  wire [6:0] T_5275;
  wire [12:0] delegable_interrupts;
  reg  reg_debug;
  reg [31:0] GEN_300;
  reg [39:0] reg_dpc;
  reg [63:0] GEN_302;
  reg [63:0] reg_dscratch;
  reg [63:0] GEN_303;
  reg  reg_tdrselect_tdrmode;
  reg [31:0] GEN_304;
  reg [61:0] reg_tdrselect_reserved;
  reg [63:0] GEN_305;
  reg  reg_tdrselect_tdrindex;
  reg [31:0] GEN_306;
  reg [3:0] reg_bp_0_control_tdrtype;
  reg [31:0] GEN_307;
  reg [4:0] reg_bp_0_control_bpamaskmax;
  reg [31:0] GEN_308;
  reg [35:0] reg_bp_0_control_reserved;
  reg [63:0] GEN_309;
  reg [7:0] reg_bp_0_control_bpaction;
  reg [31:0] GEN_310;
  reg [3:0] reg_bp_0_control_bpmatch;
  reg [31:0] GEN_311;
  reg  reg_bp_0_control_m;
  reg [31:0] GEN_312;
  reg  reg_bp_0_control_h;
  reg [31:0] GEN_313;
  reg  reg_bp_0_control_s;
  reg [31:0] GEN_314;
  reg  reg_bp_0_control_u;
  reg [31:0] GEN_315;
  reg  reg_bp_0_control_r;
  reg [31:0] GEN_316;
  reg  reg_bp_0_control_w;
  reg [31:0] GEN_317;
  reg  reg_bp_0_control_x;
  reg [31:0] GEN_318;
  reg [38:0] reg_bp_0_address;
  reg [63:0] GEN_319;
  reg [3:0] reg_bp_1_control_tdrtype;
  reg [31:0] GEN_320;
  reg [4:0] reg_bp_1_control_bpamaskmax;
  reg [31:0] GEN_321;
  reg [35:0] reg_bp_1_control_reserved;
  reg [63:0] GEN_322;
  reg [7:0] reg_bp_1_control_bpaction;
  reg [31:0] GEN_323;
  reg [3:0] reg_bp_1_control_bpmatch;
  reg [31:0] GEN_324;
  reg  reg_bp_1_control_m;
  reg [31:0] GEN_325;
  reg  reg_bp_1_control_h;
  reg [31:0] GEN_326;
  reg  reg_bp_1_control_s;
  reg [31:0] GEN_327;
  reg  reg_bp_1_control_u;
  reg [31:0] GEN_329;
  reg  reg_bp_1_control_r;
  reg [31:0] GEN_330;
  reg  reg_bp_1_control_w;
  reg [31:0] GEN_332;
  reg  reg_bp_1_control_x;
  reg [31:0] GEN_333;
  reg [38:0] reg_bp_1_address;
  reg [63:0] GEN_334;
  reg [63:0] reg_mie;
  reg [63:0] GEN_335;
  reg [63:0] reg_mideleg;
  reg [63:0] GEN_336;
  reg [63:0] reg_medeleg;
  reg [63:0] GEN_338;
  reg  reg_mip_rocc;
  reg [31:0] GEN_339;
  reg  reg_mip_meip;
  reg [31:0] GEN_341;
  reg  reg_mip_heip;
  reg [31:0] GEN_342;
  reg  reg_mip_seip;
  reg [31:0] GEN_344;
  reg  reg_mip_ueip;
  reg [31:0] GEN_345;
  reg  reg_mip_mtip;
  reg [31:0] GEN_347;
  reg  reg_mip_htip;
  reg [31:0] GEN_348;
  reg  reg_mip_stip;
  reg [31:0] GEN_350;
  reg  reg_mip_utip;
  reg [31:0] GEN_351;
  reg  reg_mip_msip;
  reg [31:0] GEN_353;
  reg  reg_mip_hsip;
  reg [31:0] GEN_354;
  reg  reg_mip_ssip;
  reg [31:0] GEN_356;
  reg  reg_mip_usip;
  reg [31:0] GEN_357;
  reg [39:0] reg_mepc;
  reg [63:0] GEN_358;
  reg [63:0] reg_mcause;
  reg [63:0] GEN_359;
  reg [39:0] reg_mbadaddr;
  reg [63:0] GEN_360;
  reg [63:0] reg_mscratch;
  reg [63:0] GEN_361;
  reg [31:0] reg_mtvec;
  reg [31:0] GEN_362;
  reg [39:0] reg_sepc;
  reg [63:0] GEN_363;
  reg [63:0] reg_scause;
  reg [63:0] GEN_364;
  reg [39:0] reg_sbadaddr;
  reg [63:0] GEN_365;
  reg [63:0] reg_sscratch;
  reg [63:0] GEN_366;
  reg [38:0] reg_stvec;
  reg [63:0] GEN_367;
  reg [19:0] reg_sptbr;
  reg [31:0] GEN_368;
  reg  reg_wfi;
  reg [31:0] GEN_369;
  reg [5:0] T_5476;
  reg [31:0] GEN_370;
  wire [6:0] GEN_597;
  wire [7:0] T_5480;
  wire [6:0] T_5481;
  wire [5:0] T_5482;
  wire [5:0] GEN_27;
  reg [57:0] T_5484;
  reg [63:0] GEN_371;
  wire  T_5485;
  wire  T_5486;
  wire [57:0] GEN_598;
  wire [58:0] T_5488;
  wire [57:0] T_5489;
  wire [57:0] GEN_28;
  reg [5:0] T_5492;
  reg [31:0] GEN_372;
  wire [6:0] GEN_599;
  wire [7:0] T_5496;
  wire [6:0] T_5497;
  wire [5:0] T_5498;
  wire [5:0] GEN_29;
  reg [57:0] T_5500;
  reg [63:0] GEN_373;
  wire  T_5501;
  wire  T_5502;
  wire [58:0] T_5504;
  wire [57:0] T_5505;
  wire [57:0] GEN_30;
  reg [5:0] T_5508;
  reg [31:0] GEN_374;
  wire [6:0] GEN_601;
  wire [7:0] T_5512;
  wire [6:0] T_5513;
  wire [5:0] T_5514;
  wire [5:0] GEN_31;
  reg [57:0] T_5516;
  reg [63:0] GEN_375;
  wire  T_5517;
  wire  T_5518;
  wire [58:0] T_5520;
  wire [57:0] T_5521;
  wire [57:0] GEN_32;
  reg [5:0] T_5524;
  reg [31:0] GEN_376;
  wire [6:0] GEN_603;
  wire [7:0] T_5528;
  wire [6:0] T_5529;
  wire [5:0] T_5530;
  wire [5:0] GEN_33;
  reg [57:0] T_5532;
  reg [63:0] GEN_377;
  wire  T_5533;
  wire  T_5534;
  wire [58:0] T_5536;
  wire [57:0] T_5537;
  wire [57:0] GEN_34;
  reg [5:0] T_5540;
  reg [31:0] GEN_378;
  wire [6:0] GEN_605;
  wire [7:0] T_5544;
  wire [6:0] T_5545;
  wire [5:0] T_5546;
  wire [5:0] GEN_35;
  reg [57:0] T_5548;
  reg [63:0] GEN_379;
  wire  T_5549;
  wire  T_5550;
  wire [58:0] T_5552;
  wire [57:0] T_5553;
  wire [57:0] GEN_36;
  reg [5:0] T_5556;
  reg [31:0] GEN_380;
  wire [6:0] GEN_607;
  wire [7:0] T_5560;
  wire [6:0] T_5561;
  wire [5:0] T_5562;
  wire [5:0] GEN_37;
  reg [57:0] T_5564;
  reg [63:0] GEN_381;
  wire  T_5565;
  wire  T_5566;
  wire [58:0] T_5568;
  wire [57:0] T_5569;
  wire [57:0] GEN_38;
  reg [5:0] T_5572;
  reg [31:0] GEN_383;
  wire [6:0] GEN_609;
  wire [7:0] T_5576;
  wire [6:0] T_5577;
  wire [5:0] T_5578;
  wire [5:0] GEN_39;
  reg [57:0] T_5580;
  reg [63:0] GEN_384;
  wire  T_5581;
  wire  T_5582;
  wire [58:0] T_5584;
  wire [57:0] T_5585;
  wire [57:0] GEN_40;
  reg [5:0] T_5588;
  reg [31:0] GEN_386;
  wire [6:0] GEN_611;
  wire [7:0] T_5592;
  wire [6:0] T_5593;
  wire [5:0] T_5594;
  wire [5:0] GEN_41;
  reg [57:0] T_5596;
  reg [63:0] GEN_387;
  wire  T_5597;
  wire  T_5598;
  wire [58:0] T_5600;
  wire [57:0] T_5601;
  wire [57:0] GEN_42;
  reg [5:0] T_5604;
  reg [31:0] GEN_388;
  wire [6:0] GEN_613;
  wire [7:0] T_5608;
  wire [6:0] T_5609;
  wire [5:0] T_5610;
  wire [5:0] GEN_43;
  reg [57:0] T_5612;
  reg [63:0] GEN_389;
  wire  T_5613;
  wire  T_5614;
  wire [58:0] T_5616;
  wire [57:0] T_5617;
  wire [57:0] GEN_44;
  reg [5:0] T_5620;
  reg [31:0] GEN_390;
  wire [6:0] GEN_615;
  wire [7:0] T_5624;
  wire [6:0] T_5625;
  wire [5:0] T_5626;
  wire [5:0] GEN_45;
  reg [57:0] T_5628;
  reg [63:0] GEN_392;
  wire  T_5629;
  wire  T_5630;
  wire [58:0] T_5632;
  wire [57:0] T_5633;
  wire [57:0] GEN_46;
  reg [5:0] T_5636;
  reg [31:0] GEN_393;
  wire [6:0] GEN_617;
  wire [7:0] T_5640;
  wire [6:0] T_5641;
  wire [5:0] T_5642;
  wire [5:0] GEN_47;
  reg [57:0] T_5644;
  reg [63:0] GEN_395;
  wire  T_5645;
  wire  T_5646;
  wire [58:0] T_5648;
  wire [57:0] T_5649;
  wire [57:0] GEN_48;
  reg [5:0] T_5652;
  reg [31:0] GEN_396;
  wire [6:0] GEN_619;
  wire [7:0] T_5656;
  wire [6:0] T_5657;
  wire [5:0] T_5658;
  wire [5:0] GEN_49;
  reg [57:0] T_5660;
  reg [63:0] GEN_398;
  wire  T_5661;
  wire  T_5662;
  wire [58:0] T_5664;
  wire [57:0] T_5665;
  wire [57:0] GEN_50;
  reg [5:0] T_5668;
  reg [31:0] GEN_399;
  wire [6:0] GEN_621;
  wire [7:0] T_5672;
  wire [6:0] T_5673;
  wire [5:0] T_5674;
  wire [5:0] GEN_51;
  reg [57:0] T_5676;
  reg [63:0] GEN_401;
  wire  T_5677;
  wire  T_5678;
  wire [58:0] T_5680;
  wire [57:0] T_5681;
  wire [57:0] GEN_52;
  reg [5:0] T_5684;
  reg [31:0] GEN_402;
  wire [6:0] GEN_623;
  wire [7:0] T_5688;
  wire [6:0] T_5689;
  wire [5:0] T_5690;
  wire [5:0] GEN_53;
  reg [57:0] T_5692;
  reg [63:0] GEN_404;
  wire  T_5693;
  wire  T_5694;
  wire [58:0] T_5696;
  wire [57:0] T_5697;
  wire [57:0] GEN_54;
  reg [5:0] T_5700;
  reg [31:0] GEN_405;
  wire [6:0] GEN_625;
  wire [7:0] T_5704;
  wire [6:0] T_5705;
  wire [5:0] T_5706;
  wire [5:0] GEN_55;
  reg [57:0] T_5708;
  reg [63:0] GEN_406;
  wire  T_5709;
  wire  T_5710;
  wire [58:0] T_5712;
  wire [57:0] T_5713;
  wire [57:0] GEN_56;
  reg [5:0] T_5716;
  reg [31:0] GEN_408;
  wire [6:0] GEN_627;
  wire [7:0] T_5720;
  wire [6:0] T_5721;
  wire [5:0] T_5722;
  wire [5:0] GEN_57;
  reg [57:0] T_5724;
  reg [63:0] GEN_409;
  wire  T_5725;
  wire  T_5726;
  wire [58:0] T_5728;
  wire [57:0] T_5729;
  wire [57:0] GEN_58;
  reg [4:0] reg_fflags;
  reg [31:0] GEN_410;
  reg [2:0] reg_frm;
  reg [31:0] GEN_411;
  reg [5:0] T_5734;
  reg [31:0] GEN_412;
  wire [6:0] GEN_629;
  wire [7:0] T_5738;
  wire [6:0] T_5739;
  wire [5:0] T_5740;
  wire [5:0] GEN_59;
  reg [57:0] T_5742;
  reg [63:0] GEN_413;
  wire  T_5743;
  wire  T_5744;
  wire [58:0] T_5746;
  wire [57:0] T_5747;
  wire [57:0] GEN_60;
  wire [63:0] T_5748;
  reg [5:0] T_5751;
  reg [31:0] GEN_414;
  wire [6:0] GEN_631;
  wire [7:0] T_5755;
  wire [6:0] T_5756;
  wire [5:0] T_5757;
  reg [57:0] T_5759;
  reg [63:0] GEN_415;
  wire  T_5760;
  wire [58:0] T_5763;
  wire [57:0] T_5764;
  wire [57:0] GEN_62;
  wire [63:0] reg_cycle;
  wire  mip_rocc;
  wire  mip_meip;
  wire  mip_heip;
  wire  mip_seip;
  wire  mip_ueip;
  wire  mip_mtip;
  wire  mip_htip;
  wire  mip_stip;
  wire  mip_utip;
  wire  mip_msip;
  wire  mip_hsip;
  wire  mip_ssip;
  wire  mip_usip;
  wire [1:0] T_5778;
  wire [2:0] T_5779;
  wire [1:0] T_5780;
  wire [2:0] T_5781;
  wire [5:0] T_5782;
  wire [1:0] T_5783;
  wire [2:0] T_5784;
  wire [1:0] T_5785;
  wire [1:0] T_5786;
  wire [3:0] T_5787;
  wire [6:0] T_5788;
  wire [12:0] T_5789;
  wire [12:0] read_mip;
  wire [63:0] GEN_633;
  wire [63:0] pending_interrupts;
  wire  T_5791;
  wire  T_5793;
  wire  T_5795;
  wire  T_5796;
  wire  T_5797;
  wire  T_5798;
  wire [63:0] T_5799;
  wire [63:0] T_5800;
  wire [63:0] m_interrupts;
  wire [1:0] GEN_634;
  wire  T_5805;
  wire  T_5807;
  wire  T_5808;
  wire  T_5809;
  wire  T_5810;
  wire [63:0] T_5811;
  wire [63:0] s_interrupts;
  wire [63:0] all_interrupts;
  wire  T_5814;
  wire  T_5815;
  wire  T_5816;
  wire  T_5817;
  wire  T_5818;
  wire  T_5819;
  wire  T_5820;
  wire  T_5821;
  wire  T_5822;
  wire  T_5823;
  wire  T_5824;
  wire  T_5825;
  wire  T_5826;
  wire  T_5827;
  wire  T_5828;
  wire  T_5829;
  wire  T_5830;
  wire  T_5831;
  wire  T_5832;
  wire  T_5833;
  wire  T_5834;
  wire  T_5835;
  wire  T_5836;
  wire  T_5837;
  wire  T_5838;
  wire  T_5839;
  wire  T_5840;
  wire  T_5841;
  wire  T_5842;
  wire  T_5843;
  wire  T_5844;
  wire  T_5845;
  wire  T_5846;
  wire  T_5847;
  wire  T_5848;
  wire  T_5849;
  wire  T_5850;
  wire  T_5851;
  wire  T_5852;
  wire  T_5853;
  wire  T_5854;
  wire  T_5855;
  wire  T_5856;
  wire  T_5857;
  wire  T_5858;
  wire  T_5859;
  wire  T_5860;
  wire  T_5861;
  wire  T_5862;
  wire  T_5863;
  wire  T_5864;
  wire  T_5865;
  wire  T_5866;
  wire  T_5867;
  wire  T_5868;
  wire  T_5869;
  wire  T_5870;
  wire  T_5871;
  wire  T_5872;
  wire  T_5873;
  wire  T_5874;
  wire  T_5875;
  wire  T_5876;
  wire [5:0] T_5942;
  wire [5:0] T_5943;
  wire [5:0] T_5944;
  wire [5:0] T_5945;
  wire [5:0] T_5946;
  wire [5:0] T_5947;
  wire [5:0] T_5948;
  wire [5:0] T_5949;
  wire [5:0] T_5950;
  wire [5:0] T_5951;
  wire [5:0] T_5952;
  wire [5:0] T_5953;
  wire [5:0] T_5954;
  wire [5:0] T_5955;
  wire [5:0] T_5956;
  wire [5:0] T_5957;
  wire [5:0] T_5958;
  wire [5:0] T_5959;
  wire [5:0] T_5960;
  wire [5:0] T_5961;
  wire [5:0] T_5962;
  wire [5:0] T_5963;
  wire [5:0] T_5964;
  wire [5:0] T_5965;
  wire [5:0] T_5966;
  wire [5:0] T_5967;
  wire [5:0] T_5968;
  wire [5:0] T_5969;
  wire [5:0] T_5970;
  wire [5:0] T_5971;
  wire [5:0] T_5972;
  wire [5:0] T_5973;
  wire [5:0] T_5974;
  wire [5:0] T_5975;
  wire [5:0] T_5976;
  wire [5:0] T_5977;
  wire [5:0] T_5978;
  wire [5:0] T_5979;
  wire [5:0] T_5980;
  wire [5:0] T_5981;
  wire [5:0] T_5982;
  wire [5:0] T_5983;
  wire [5:0] T_5984;
  wire [5:0] T_5985;
  wire [5:0] T_5986;
  wire [5:0] T_5987;
  wire [5:0] T_5988;
  wire [5:0] T_5989;
  wire [5:0] T_5990;
  wire [5:0] T_5991;
  wire [5:0] T_5992;
  wire [5:0] T_5993;
  wire [5:0] T_5994;
  wire [5:0] T_5995;
  wire [5:0] T_5996;
  wire [5:0] T_5997;
  wire [5:0] T_5998;
  wire [5:0] T_5999;
  wire [5:0] T_6000;
  wire [5:0] T_6001;
  wire [5:0] T_6002;
  wire [5:0] T_6003;
  wire [5:0] T_6004;
  wire [63:0] GEN_636;
  wire [64:0] T_6005;
  wire [63:0] interruptCause;
  wire [63:0] GEN_637;
  wire  T_6007;
  wire  T_6012;
  wire  GEN_63;
  wire [63:0] GEN_64;
  wire  system_insn;
  wire  T_6015;
  wire  T_6017;
  wire  cpu_ren;
  wire [1:0] T_6018;
  wire [1:0] T_6019;
  wire [2:0] T_6020;
  wire [4:0] T_6021;
  wire [1:0] T_6022;
  wire [2:0] T_6023;
  wire [3:0] T_6024;
  wire [4:0] T_6025;
  wire [7:0] T_6026;
  wire [12:0] T_6027;
  wire [2:0] T_6028;
  wire [4:0] T_6029;
  wire [9:0] T_6030;
  wire [10:0] T_6031;
  wire [15:0] T_6032;
  wire [31:0] T_6033;
  wire [33:0] T_6034;
  wire [2:0] T_6035;
  wire [3:0] T_6036;
  wire [37:0] T_6037;
  wire [53:0] T_6038;
  wire [66:0] T_6039;
  wire [63:0] read_mstatus;
  wire [62:0] T_6040;
  wire [63:0] T_6041;
  wire  GEN_0;
  wire  GEN_65;
  wire  GEN_1;
  wire  GEN_66;
  wire [1:0] T_6056;
  wire  GEN_2;
  wire  GEN_67;
  wire [2:0] T_6057;
  wire  GEN_3;
  wire  GEN_68;
  wire  GEN_4;
  wire  GEN_69;
  wire [1:0] T_6058;
  wire  GEN_5;
  wire  GEN_70;
  wire [2:0] T_6059;
  wire [5:0] T_6060;
  wire [7:0] GEN_6;
  wire [7:0] GEN_71;
  wire [3:0] GEN_7;
  wire [3:0] GEN_72;
  wire [11:0] T_6061;
  wire  GEN_8;
  wire  GEN_73;
  wire [12:0] T_6062;
  wire [3:0] GEN_9;
  wire [3:0] GEN_74;
  wire [4:0] GEN_10;
  wire [4:0] GEN_75;
  wire [8:0] T_6063;
  wire [35:0] GEN_11;
  wire [35:0] GEN_76;
  wire [44:0] T_6064;
  wire [57:0] T_6065;
  wire [63:0] T_6066;
  wire  T_6089;
  wire [23:0] GEN_638;
  wire [24:0] T_6091;
  wire [23:0] T_6092;
  wire [63:0] T_6093;
  wire  T_6094;
  wire [23:0] GEN_639;
  wire [24:0] T_6096;
  wire [23:0] T_6097;
  wire [63:0] T_6098;
  wire [2:0] T_6099;
  wire [1:0] T_6100;
  wire [4:0] T_6101;
  wire [3:0] T_6102;
  wire [1:0] T_6103;
  wire [5:0] T_6104;
  wire [10:0] T_6105;
  wire [1:0] T_6106;
  wire [1:0] T_6107;
  wire [3:0] T_6108;
  wire [12:0] T_6109;
  wire [2:0] T_6110;
  wire [3:0] T_6111;
  wire [16:0] T_6112;
  wire [20:0] T_6113;
  wire [31:0] T_6114;
  wire [7:0] T_6115;
  wire [63:0] T_6116;
  wire [63:0] T_6117;
  wire  T_6118_debug;
  wire [1:0] T_6118_prv;
  wire  T_6118_sd;
  wire [30:0] T_6118_zero3;
  wire  T_6118_sd_rv32;
  wire [1:0] T_6118_zero2;
  wire [4:0] T_6118_vm;
  wire [4:0] T_6118_zero1;
  wire  T_6118_pum;
  wire  T_6118_mprv;
  wire [1:0] T_6118_xs;
  wire [1:0] T_6118_fs;
  wire [1:0] T_6118_mpp;
  wire [1:0] T_6118_hpp;
  wire  T_6118_spp;
  wire  T_6118_mpie;
  wire  T_6118_hpie;
  wire  T_6118_spie;
  wire  T_6118_upie;
  wire  T_6118_mie;
  wire  T_6118_hie;
  wire  T_6118_sie;
  wire  T_6118_uie;
  wire [1:0] T_6150;
  wire [1:0] T_6151;
  wire [2:0] T_6152;
  wire [4:0] T_6153;
  wire [1:0] T_6154;
  wire [2:0] T_6155;
  wire [3:0] T_6156;
  wire [4:0] T_6157;
  wire [7:0] T_6158;
  wire [12:0] T_6159;
  wire [2:0] T_6160;
  wire [4:0] T_6161;
  wire [9:0] T_6162;
  wire [10:0] T_6163;
  wire [15:0] T_6164;
  wire [31:0] T_6165;
  wire [33:0] T_6166;
  wire [2:0] T_6167;
  wire [3:0] T_6168;
  wire [37:0] T_6169;
  wire [53:0] T_6170;
  wire [66:0] T_6171;
  wire [63:0] T_6172;
  wire  T_6173;
  wire [23:0] GEN_641;
  wire [24:0] T_6175;
  wire [23:0] T_6176;
  wire [63:0] T_6177;
  wire  T_6179;
  wire [23:0] GEN_642;
  wire [24:0] T_6181;
  wire [23:0] T_6182;
  wire [63:0] T_6183;
  wire  T_6184;
  wire [24:0] GEN_643;
  wire [25:0] T_6186;
  wire [24:0] T_6187;
  wire [63:0] T_6188;
  wire [11:0] GEN_644;
  wire  T_6194;
  wire [11:0] GEN_645;
  wire  T_6196;
  wire [11:0] GEN_646;
  wire  T_6198;
  wire  T_6200;
  wire  T_6202;
  wire  T_6204;
  wire  T_6206;
  wire  T_6208;
  wire [11:0] GEN_647;
  wire  T_6210;
  wire [11:0] GEN_648;
  wire  T_6212;
  wire [11:0] GEN_649;
  wire  T_6214;
  wire [11:0] GEN_650;
  wire  T_6216;
  wire  T_6218;
  wire [11:0] GEN_651;
  wire  T_6220;
  wire [11:0] GEN_652;
  wire  T_6222;
  wire [11:0] GEN_653;
  wire  T_6224;
  wire [11:0] GEN_654;
  wire  T_6226;
  wire [11:0] GEN_655;
  wire  T_6228;
  wire [11:0] GEN_656;
  wire  T_6230;
  wire [11:0] GEN_657;
  wire  T_6232;
  wire [11:0] GEN_658;
  wire  T_6234;
  wire [11:0] GEN_659;
  wire  T_6236;
  wire [11:0] GEN_660;
  wire  T_6238;
  wire  T_6240;
  wire [11:0] GEN_661;
  wire  T_6242;
  wire [11:0] GEN_662;
  wire  T_6244;
  wire [11:0] GEN_663;
  wire  T_6246;
  wire [11:0] GEN_664;
  wire  T_6248;
  wire [11:0] GEN_665;
  wire  T_6250;
  wire [11:0] GEN_666;
  wire  T_6252;
  wire [11:0] GEN_667;
  wire  T_6254;
  wire [11:0] GEN_668;
  wire  T_6256;
  wire [11:0] GEN_669;
  wire  T_6258;
  wire [11:0] GEN_670;
  wire  T_6260;
  wire [11:0] GEN_671;
  wire  T_6262;
  wire [11:0] GEN_672;
  wire  T_6264;
  wire [11:0] GEN_673;
  wire  T_6266;
  wire [11:0] GEN_674;
  wire  T_6268;
  wire [11:0] GEN_675;
  wire  T_6270;
  wire [11:0] GEN_676;
  wire  T_6272;
  wire [11:0] GEN_677;
  wire  T_6274;
  wire [11:0] GEN_678;
  wire  T_6276;
  wire [11:0] GEN_679;
  wire  T_6278;
  wire [11:0] GEN_680;
  wire  T_6280;
  wire  T_6281;
  wire  T_6282;
  wire  T_6283;
  wire  T_6284;
  wire  T_6285;
  wire  T_6286;
  wire  T_6287;
  wire  T_6288;
  wire  T_6289;
  wire  T_6290;
  wire  T_6291;
  wire  T_6292;
  wire  T_6293;
  wire  T_6294;
  wire  T_6295;
  wire  T_6296;
  wire  T_6297;
  wire  T_6298;
  wire  T_6299;
  wire  T_6300;
  wire  T_6301;
  wire  T_6302;
  wire  T_6303;
  wire  T_6304;
  wire  T_6305;
  wire  T_6306;
  wire  T_6307;
  wire  T_6308;
  wire  T_6309;
  wire  T_6310;
  wire  T_6311;
  wire  T_6312;
  wire  T_6313;
  wire  T_6314;
  wire  T_6315;
  wire  T_6316;
  wire  T_6317;
  wire  T_6318;
  wire  T_6319;
  wire  T_6320;
  wire  T_6321;
  wire  T_6322;
  wire  addr_valid;
  wire  T_6323;
  wire  fp_csr;
  wire  T_6325;
  wire [1:0] T_6326;
  wire [1:0] T_6327;
  wire [1:0] GEN_681;
  wire  T_6329;
  wire [1:0] T_6330;
  wire [2:0] csr_addr_priv;
  wire [2:0] T_6331;
  wire  priv_sufficient;
  wire [1:0] T_6332;
  wire [1:0] T_6333;
  wire  read_only;
  wire  T_6335;
  wire  T_6336;
  wire  cpu_wen;
  wire  T_6338;
  wire  wen;
  wire  T_6339;
  wire  T_6340;
  wire  T_6341;
  wire [63:0] T_6343;
  wire  T_6344;
  wire [63:0] T_6346;
  wire [63:0] T_6347;
  wire [63:0] T_6350;
  wire [63:0] T_6351;
  wire [63:0] wdata;
  wire  do_system_insn;
  wire [2:0] T_6353;
  wire [7:0] GEN_683;
  wire [7:0] opcode;
  wire  T_6354;
  wire  insn_call;
  wire  T_6355;
  wire  insn_break;
  wire  T_6356;
  wire  insn_ret;
  wire  T_6357;
  wire  insn_sfence_vm;
  wire  T_6358;
  wire  insn_wfi;
  wire  T_6359;
  wire  T_6361;
  wire  T_6363;
  wire  T_6364;
  wire  T_6366;
  wire  T_6368;
  wire  T_6369;
  wire  T_6370;
  wire  T_6371;
  wire  T_6372;
  wire  T_6375;
  wire  T_6376;
  wire  T_6377;
  wire  csr_xcpt;
  wire  GEN_77;
  wire [12:0] GEN_685;
  wire  T_6380;
  wire  GEN_78;
  wire  T_6383;
  wire [3:0] GEN_686;
  wire [4:0] T_6385;
  wire [3:0] T_6386;
  wire [1:0] T_6389;
  wire [3:0] T_6390;
  wire [63:0] cause;
  wire [5:0] cause_lsbs;
  wire  T_6391;
  wire [5:0] GEN_687;
  wire  T_6393;
  wire  causeIsDebugInt;
  wire [63:0] GEN_688;
  wire  T_6395;
  wire [1:0] T_6396;
  wire [1:0] T_6397;
  wire [3:0] T_6398;
  wire [3:0] T_6399;
  wire  T_6400;
  wire  causeIsDebugBreak;
  wire  T_6402;
  wire  T_6403;
  wire [63:0] T_6409;
  wire  T_6410;
  wire [63:0] T_6411;
  wire  T_6412;
  wire  T_6413;
  wire  delegate;
  wire [11:0] debugTVec;
  wire [39:0] T_6417;
  wire [39:0] T_6418;
  wire [39:0] tvec;
  wire  T_6420;
  wire  T_6422;
  wire [39:0] T_6424;
  wire [39:0] epc;
  wire  T_6425;
  wire [39:0] T_6426;
  wire [1:0] T_6427;
  wire  T_6429;
  wire [1:0] T_6430;
  wire  T_6432;
  wire  T_6433;
  wire [39:0] T_6435;
  wire [39:0] GEN_691;
  wire [39:0] T_6437;
  wire [39:0] T_6438;
  wire [63:0] T_6439;
  wire  T_6440;
  wire [1:0] T_6444;
  wire  GEN_79;
  wire [39:0] GEN_80;
  wire [2:0] GEN_81;
  wire [1:0] GEN_82;
  wire  T_6446;
  wire  T_6447;
  wire [39:0] GEN_83;
  wire [63:0] GEN_84;
  wire [39:0] GEN_85;
  wire  GEN_86;
  wire [1:0] GEN_87;
  wire  GEN_88;
  wire [1:0] GEN_89;
  wire  T_6453;
  wire  T_6454;
  wire [39:0] GEN_90;
  wire [63:0] GEN_91;
  wire [39:0] GEN_92;
  wire  GEN_93;
  wire [1:0] GEN_94;
  wire  GEN_95;
  wire [1:0] GEN_96;
  wire  GEN_97;
  wire [39:0] GEN_98;
  wire [2:0] GEN_99;
  wire [1:0] GEN_100;
  wire [39:0] GEN_101;
  wire [63:0] GEN_102;
  wire [39:0] GEN_103;
  wire  GEN_104;
  wire [1:0] GEN_105;
  wire  GEN_106;
  wire [1:0] GEN_107;
  wire [39:0] GEN_108;
  wire [63:0] GEN_109;
  wire [39:0] GEN_110;
  wire  GEN_111;
  wire [1:0] GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire [1:0] GEN_117;
  wire [1:0] GEN_118;
  wire  T_6466;
  wire  T_6467;
  wire [1:0] GEN_119;
  wire  GEN_120;
  wire  T_6472;
  wire  T_6473;
  wire  T_6474;
  wire  GEN_121;
  wire  T_6476;
  wire  T_6479;
  wire  T_6480;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire [1:0] GEN_126;
  wire [1:0] GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire [1:0] GEN_130;
  wire [1:0] GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire [1:0] GEN_135;
  wire [1:0] T_6485;
  wire [1:0] GEN_692;
  wire [2:0] T_6486;
  wire [1:0] T_6487;
  wire [2:0] T_6488;
  wire [2:0] GEN_693;
  wire [3:0] T_6489;
  wire [2:0] T_6490;
  wire [2:0] GEN_694;
  wire  T_6492;
  wire  T_6493;
  wire  T_6495;
  wire [63:0] T_6497;
  wire [63:0] T_6499;
  wire [38:0] GEN_12;
  wire [38:0] GEN_136;
  wire [38:0] T_6501;
  wire [63:0] T_6509;
  wire [63:0] T_6511;
  wire [63:0] T_6521;
  wire [63:0] T_6523;
  wire [31:0] T_6525;
  wire [12:0] T_6527;
  wire [63:0] T_6529;
  wire [63:0] T_6531;
  wire [63:0] T_6533;
  wire [63:0] T_6535;
  wire [63:0] T_6537;
  wire [63:0] T_6539;
  wire [63:0] T_6541;
  wire  T_6543;
  wire [31:0] T_6545;
  wire [39:0] T_6547;
  wire [63:0] T_6549;
  wire [4:0] T_6551;
  wire [2:0] T_6553;
  wire [7:0] T_6555;
  wire [63:0] T_6557;
  wire [63:0] T_6559;
  wire [63:0] T_6561;
  wire [63:0] T_6563;
  wire [63:0] T_6565;
  wire [63:0] T_6567;
  wire [19:0] T_6569;
  wire [63:0] T_6573;
  wire [63:0] T_6575;
  wire [63:0] T_6585;
  wire [63:0] GEN_695;
  wire [63:0] T_6586;
  wire [63:0] T_6587;
  wire [63:0] T_6588;
  wire [63:0] T_6589;
  wire [63:0] T_6590;
  wire [63:0] T_6591;
  wire [63:0] T_6592;
  wire [63:0] T_6593;
  wire [63:0] T_6594;
  wire [63:0] T_6595;
  wire [63:0] T_6596;
  wire [63:0] T_6597;
  wire [63:0] GEN_703;
  wire [63:0] T_6598;
  wire [63:0] GEN_704;
  wire [63:0] T_6599;
  wire [63:0] T_6600;
  wire [63:0] T_6601;
  wire [63:0] T_6602;
  wire [63:0] T_6603;
  wire [63:0] T_6604;
  wire [63:0] T_6605;
  wire [63:0] T_6606;
  wire [63:0] GEN_705;
  wire [63:0] T_6607;
  wire [63:0] GEN_706;
  wire [63:0] T_6608;
  wire [63:0] GEN_707;
  wire [63:0] T_6609;
  wire [63:0] T_6610;
  wire [63:0] GEN_708;
  wire [63:0] T_6611;
  wire [63:0] GEN_709;
  wire [63:0] T_6612;
  wire [63:0] GEN_710;
  wire [63:0] T_6613;
  wire [63:0] T_6614;
  wire [63:0] T_6615;
  wire [63:0] T_6616;
  wire [63:0] T_6617;
  wire [63:0] T_6618;
  wire [63:0] T_6619;
  wire [63:0] GEN_711;
  wire [63:0] T_6620;
  wire [63:0] T_6621;
  wire [63:0] T_6622;
  wire [63:0] T_6623;
  wire [63:0] T_6624;
  wire [63:0] T_6625;
  wire [63:0] T_6626;
  wire [63:0] T_6627;
  wire [63:0] T_6628;
  wire [4:0] T_6629;
  wire [4:0] GEN_137;
  wire [1:0] supportedModes_0;
  wire [1:0] supportedModes_1;
  wire [1:0] supportedModes_2;
  wire  T_6687_debug;
  wire [1:0] T_6687_prv;
  wire  T_6687_sd;
  wire [30:0] T_6687_zero3;
  wire  T_6687_sd_rv32;
  wire [1:0] T_6687_zero2;
  wire [4:0] T_6687_vm;
  wire [4:0] T_6687_zero1;
  wire  T_6687_pum;
  wire  T_6687_mprv;
  wire [1:0] T_6687_xs;
  wire [1:0] T_6687_fs;
  wire [1:0] T_6687_mpp;
  wire [1:0] T_6687_hpp;
  wire  T_6687_spp;
  wire  T_6687_mpie;
  wire  T_6687_hpie;
  wire  T_6687_spie;
  wire  T_6687_upie;
  wire  T_6687_mie;
  wire  T_6687_hie;
  wire  T_6687_sie;
  wire  T_6687_uie;
  wire [66:0] T_6712;
  wire  T_6713;
  wire  T_6714;
  wire  T_6715;
  wire  T_6716;
  wire  T_6717;
  wire  T_6718;
  wire  T_6719;
  wire  T_6720;
  wire  T_6721;
  wire [1:0] T_6722;
  wire [1:0] T_6723;
  wire [1:0] T_6724;
  wire [1:0] T_6725;
  wire  T_6726;
  wire  T_6727;
  wire [4:0] T_6728;
  wire [4:0] T_6729;
  wire [1:0] T_6730;
  wire  T_6731;
  wire [30:0] T_6732;
  wire  T_6733;
  wire [1:0] T_6734;
  wire  T_6735;
  wire  T_6736;
  wire  T_6737;
  wire  T_6738;
  wire  T_6741;
  wire  T_6742;
  wire [1:0] GEN_138;
  wire [4:0] GEN_717;
  wire  T_6744;
  wire [4:0] GEN_139;
  wire [4:0] GEN_718;
  wire  T_6747;
  wire [4:0] GEN_140;
  wire  T_6750;
  wire [1:0] GEN_720;
  wire [2:0] T_6752;
  wire [1:0] T_6753;
  wire  GEN_165;
  wire  GEN_166;
  wire  GEN_167;
  wire [1:0] GEN_168;
  wire  GEN_169;
  wire [1:0] GEN_170;
  wire  GEN_171;
  wire  GEN_172;
  wire [4:0] GEN_173;
  wire [1:0] GEN_174;
  wire  T_6782_rocc;
  wire  T_6782_meip;
  wire  T_6782_heip;
  wire  T_6782_seip;
  wire  T_6782_ueip;
  wire  T_6782_mtip;
  wire  T_6782_htip;
  wire  T_6782_stip;
  wire  T_6782_utip;
  wire  T_6782_msip;
  wire  T_6782_hsip;
  wire  T_6782_ssip;
  wire  T_6782_usip;
  wire  T_6796;
  wire  T_6797;
  wire  T_6798;
  wire  T_6799;
  wire  T_6800;
  wire  T_6801;
  wire  T_6802;
  wire  T_6803;
  wire  T_6804;
  wire  T_6805;
  wire  T_6806;
  wire  T_6807;
  wire  T_6808;
  wire  GEN_188;
  wire  GEN_189;
  wire [63:0] GEN_721;
  wire [63:0] T_6809;
  wire [63:0] GEN_190;
  wire [63:0] T_6810;
  wire [63:0] T_6812;
  wire [63:0] T_6813;
  wire [63:0] GEN_191;
  wire [63:0] GEN_192;
  wire [61:0] T_6814;
  wire [63:0] GEN_723;
  wire [63:0] T_6815;
  wire [63:0] GEN_193;
  wire [63:0] T_6817;
  wire [63:0] GEN_194;
  wire [39:0] T_6818;
  wire [39:0] GEN_195;
  wire [63:0] GEN_196;
  wire [63:0] GEN_197;
  wire [58:0] T_6819;
  wire [63:0] GEN_198;
  wire [63:0] GEN_199;
  wire [1:0] T_6856_xdebugver;
  wire  T_6856_ndreset;
  wire  T_6856_fullreset;
  wire [11:0] T_6856_hwbpcount;
  wire  T_6856_ebreakm;
  wire  T_6856_ebreakh;
  wire  T_6856_ebreaks;
  wire  T_6856_ebreaku;
  wire  T_6856_zero2;
  wire  T_6856_stopcycle;
  wire  T_6856_stoptime;
  wire [2:0] T_6856_cause;
  wire  T_6856_debugint;
  wire  T_6856_zero1;
  wire  T_6856_halt;
  wire  T_6856_step;
  wire [1:0] T_6856_prv;
  wire [1:0] T_6874;
  wire [2:0] T_6879;
  wire  T_6884;
  wire  T_6885;
  wire  T_6886;
  wire [11:0] T_6887;
  wire  T_6888;
  wire  T_6889;
  wire [1:0] T_6890;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire [1:0] GEN_221;
  wire [63:0] GEN_222;
  wire [63:0] GEN_223;
  wire  T_6943_debug;
  wire [1:0] T_6943_prv;
  wire  T_6943_sd;
  wire [30:0] T_6943_zero3;
  wire  T_6943_sd_rv32;
  wire [1:0] T_6943_zero2;
  wire [4:0] T_6943_vm;
  wire [4:0] T_6943_zero1;
  wire  T_6943_pum;
  wire  T_6943_mprv;
  wire [1:0] T_6943_xs;
  wire [1:0] T_6943_fs;
  wire [1:0] T_6943_mpp;
  wire [1:0] T_6943_hpp;
  wire  T_6943_spp;
  wire  T_6943_mpie;
  wire  T_6943_hpie;
  wire  T_6943_spie;
  wire  T_6943_upie;
  wire  T_6943_mie;
  wire  T_6943_hie;
  wire  T_6943_sie;
  wire  T_6943_uie;
  wire [66:0] T_6968;
  wire  T_6969;
  wire  T_6970;
  wire  T_6971;
  wire  T_6972;
  wire  T_6973;
  wire  T_6974;
  wire  T_6975;
  wire  T_6976;
  wire  T_6977;
  wire [1:0] T_6978;
  wire [1:0] T_6979;
  wire [1:0] T_6980;
  wire [1:0] T_6981;
  wire  T_6982;
  wire  T_6983;
  wire [4:0] T_6984;
  wire [4:0] T_6985;
  wire [1:0] T_6986;
  wire  T_6987;
  wire [30:0] T_6988;
  wire  T_6989;
  wire [1:0] T_6990;
  wire  T_6991;
  wire  T_6993;
  wire [1:0] GEN_726;
  wire [2:0] T_6995;
  wire [1:0] T_6996;
  wire  GEN_248;
  wire  GEN_249;
  wire [1:0] GEN_250;
  wire  GEN_251;
  wire [1:0] GEN_252;
  wire  T_7025_rocc;
  wire  T_7025_meip;
  wire  T_7025_heip;
  wire  T_7025_seip;
  wire  T_7025_ueip;
  wire  T_7025_mtip;
  wire  T_7025_htip;
  wire  T_7025_stip;
  wire  T_7025_utip;
  wire  T_7025_msip;
  wire  T_7025_hsip;
  wire  T_7025_ssip;
  wire  T_7025_usip;
  wire  GEN_266;
  wire [63:0] T_7053;
  wire [63:0] T_7054;
  wire [63:0] T_7055;
  wire [63:0] GEN_267;
  wire [63:0] GEN_268;
  wire [63:0] GEN_269;
  wire [63:0] GEN_270;
  wire [63:0] GEN_271;
  wire [63:0] GEN_272;
  wire [39:0] GEN_273;
  wire [63:0] GEN_729;
  wire [63:0] T_7063;
  wire [63:0] GEN_274;
  wire [63:0] GEN_730;
  wire [63:0] T_7064;
  wire [63:0] GEN_275;
  wire  T_7073_tdrmode;
  wire [61:0] T_7073_reserved;
  wire  T_7073_tdrindex;
  wire [61:0] T_7078;
  wire  T_7079;
  wire  GEN_276;
  wire  T_7080;
  wire [3:0] T_7107_tdrtype;
  wire [4:0] T_7107_bpamaskmax;
  wire [35:0] T_7107_reserved;
  wire [7:0] T_7107_bpaction;
  wire [3:0] T_7107_bpmatch;
  wire  T_7107_m;
  wire  T_7107_h;
  wire  T_7107_s;
  wire  T_7107_u;
  wire  T_7107_r;
  wire  T_7107_w;
  wire  T_7107_x;
  wire [3:0] T_7127;
  wire [7:0] T_7128;
  wire [35:0] T_7129;
  wire [4:0] T_7130;
  wire [3:0] T_7131;
  wire [3:0] GEN_13;
  wire [4:0] GEN_14;
  wire [35:0] GEN_15;
  wire [7:0] GEN_16;
  wire [3:0] GEN_17;
  wire [3:0] GEN_285;
  wire  GEN_18;
  wire  GEN_287;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_291;
  wire  GEN_21;
  wire  GEN_293;
  wire  GEN_22;
  wire  GEN_295;
  wire  GEN_23;
  wire  GEN_297;
  wire  GEN_24;
  wire  GEN_299;
  wire [3:0] GEN_731;
  wire [3:0] T_7161;
  wire [3:0] GEN_25;
  wire [3:0] GEN_301;
  wire [3:0] GEN_328;
  wire  GEN_331;
  wire  GEN_337;
  wire  GEN_340;
  wire  GEN_343;
  wire  GEN_346;
  wire  GEN_349;
  wire [38:0] GEN_26;
  wire [38:0] GEN_352;
  wire [38:0] GEN_355;
  wire [3:0] GEN_382;
  wire  GEN_385;
  wire  GEN_391;
  wire  GEN_394;
  wire  GEN_397;
  wire  GEN_400;
  wire  GEN_403;
  wire [38:0] GEN_407;
  wire  GEN_433;
  wire  GEN_434;
  wire  GEN_435;
  wire [1:0] GEN_436;
  wire  GEN_437;
  wire [1:0] GEN_438;
  wire  GEN_439;
  wire  GEN_440;
  wire [4:0] GEN_441;
  wire [1:0] GEN_442;
  wire  GEN_456;
  wire  GEN_457;
  wire [63:0] GEN_458;
  wire [63:0] GEN_459;
  wire [63:0] GEN_460;
  wire [63:0] GEN_461;
  wire [63:0] GEN_462;
  wire [39:0] GEN_463;
  wire [63:0] GEN_464;
  wire [63:0] GEN_465;
  wire  GEN_483;
  wire  GEN_484;
  wire  GEN_485;
  wire  GEN_486;
  wire [1:0] GEN_487;
  wire [63:0] GEN_488;
  wire [63:0] GEN_489;
  wire [63:0] GEN_527;
  wire [63:0] GEN_528;
  wire [63:0] GEN_529;
  wire [63:0] GEN_530;
  wire [63:0] GEN_531;
  wire [39:0] GEN_532;
  wire [63:0] GEN_533;
  wire [63:0] GEN_534;
  wire  GEN_538;
  wire [3:0] GEN_564;
  wire  GEN_567;
  wire  GEN_573;
  wire  GEN_576;
  wire  GEN_579;
  wire  GEN_582;
  wire  GEN_585;
  wire [38:0] GEN_589;
  wire  GEN_591;
  wire  GEN_592;
  wire  GEN_593;
  wire [3:0] T_7226_control_tdrtype;
  wire [4:0] T_7226_control_bpamaskmax;
  wire [35:0] T_7226_control_reserved;
  wire [7:0] T_7226_control_bpaction;
  wire [3:0] T_7226_control_bpmatch;
  wire  T_7226_control_m;
  wire  T_7226_control_h;
  wire  T_7226_control_s;
  wire  T_7226_control_u;
  wire  T_7226_control_r;
  wire  T_7226_control_w;
  wire  T_7226_control_x;
  wire [38:0] T_7226_address;
  wire [102:0] T_7242;
  wire [38:0] T_7243;
  wire  T_7244;
  wire  T_7245;
  wire  T_7246;
  wire  T_7247;
  wire  T_7248;
  wire  T_7249;
  wire  T_7250;
  wire [3:0] T_7251;
  wire [7:0] T_7252;
  wire [35:0] T_7253;
  wire [4:0] T_7254;
  wire [3:0] T_7255;
  reg [1:0] GEN_61;
  reg [31:0] GEN_416;
  reg  GEN_141;
  reg [31:0] GEN_417;
  reg [6:0] GEN_142;
  reg [31:0] GEN_418;
  reg [4:0] GEN_143;
  reg [31:0] GEN_419;
  reg [4:0] GEN_144;
  reg [31:0] GEN_420;
  reg  GEN_145;
  reg [31:0] GEN_421;
  reg  GEN_146;
  reg [31:0] GEN_422;
  reg  GEN_147;
  reg [31:0] GEN_423;
  reg [4:0] GEN_148;
  reg [31:0] GEN_424;
  reg [6:0] GEN_149;
  reg [31:0] GEN_425;
  reg [63:0] GEN_150;
  reg [63:0] GEN_426;
  reg [63:0] GEN_151;
  reg [63:0] GEN_427;
  reg  GEN_152;
  reg [31:0] GEN_428;
  reg  GEN_153;
  reg [31:0] GEN_429;
  reg  GEN_154;
  reg [31:0] GEN_430;
  reg  GEN_155;
  reg [31:0] GEN_431;
  reg [39:0] GEN_156;
  reg [63:0] GEN_432;
  reg [8:0] GEN_157;
  reg [31:0] GEN_443;
  reg [4:0] GEN_158;
  reg [31:0] GEN_444;
  reg [2:0] GEN_159;
  reg [31:0] GEN_445;
  reg [63:0] GEN_160;
  reg [63:0] GEN_446;
  reg  GEN_161;
  reg [31:0] GEN_447;
  reg  GEN_162;
  reg [31:0] GEN_448;
  reg [63:0] GEN_163;
  reg [63:0] GEN_449;
  reg [63:0] GEN_164;
  reg [63:0] GEN_450;
  reg  GEN_175;
  reg [31:0] GEN_451;
  reg  GEN_176;
  reg [31:0] GEN_452;
  reg  GEN_177;
  reg [31:0] GEN_453;
  reg  GEN_178;
  reg [31:0] GEN_454;
  reg  GEN_179;
  reg [31:0] GEN_455;
  reg  GEN_180;
  reg [31:0] GEN_466;
  reg  GEN_181;
  reg [31:0] GEN_467;
  reg [1:0] GEN_182;
  reg [31:0] GEN_468;
  reg  GEN_183;
  reg [31:0] GEN_469;
  reg [30:0] GEN_184;
  reg [31:0] GEN_470;
  reg  GEN_185;
  reg [31:0] GEN_471;
  reg [1:0] GEN_186;
  reg [31:0] GEN_472;
  reg [4:0] GEN_187;
  reg [31:0] GEN_473;
  reg [4:0] GEN_200;
  reg [31:0] GEN_474;
  reg  GEN_201;
  reg [31:0] GEN_475;
  reg  GEN_202;
  reg [31:0] GEN_476;
  reg [1:0] GEN_203;
  reg [31:0] GEN_477;
  reg [1:0] GEN_204;
  reg [31:0] GEN_478;
  reg [1:0] GEN_205;
  reg [31:0] GEN_479;
  reg [1:0] GEN_206;
  reg [31:0] GEN_480;
  reg  GEN_207;
  reg [31:0] GEN_481;
  reg  GEN_208;
  reg [31:0] GEN_482;
  reg  GEN_209;
  reg [31:0] GEN_490;
  reg  GEN_210;
  reg [31:0] GEN_491;
  reg  GEN_211;
  reg [31:0] GEN_492;
  reg  GEN_212;
  reg [31:0] GEN_493;
  reg  GEN_213;
  reg [31:0] GEN_494;
  reg  GEN_214;
  reg [31:0] GEN_495;
  reg  GEN_215;
  reg [31:0] GEN_496;
  reg  GEN_216;
  reg [31:0] GEN_497;
  reg  GEN_224;
  reg [31:0] GEN_498;
  reg [2:0] GEN_225;
  reg [31:0] GEN_499;
  reg [1:0] GEN_226;
  reg [31:0] GEN_500;
  reg [2:0] GEN_227;
  reg [31:0] GEN_501;
  reg  GEN_228;
  reg [31:0] GEN_502;
  reg [3:0] GEN_229;
  reg [31:0] GEN_503;
  reg [63:0] GEN_230;
  reg [63:0] GEN_504;
  reg  GEN_231;
  reg [31:0] GEN_505;
  reg  GEN_232;
  reg [31:0] GEN_506;
  reg [64:0] GEN_233;
  reg [95:0] GEN_507;
  reg [4:0] GEN_234;
  reg [31:0] GEN_508;
  reg  GEN_235;
  reg [31:0] GEN_509;
  reg  GEN_236;
  reg [31:0] GEN_510;
  assign io_rw_rdata = T_6628;
  assign io_csr_stall = reg_wfi;
  assign io_csr_xcpt = csr_xcpt;
  assign io_eret = insn_ret;
  assign io_prv = GEN_61;
  assign io_status_debug = reg_debug;
  assign io_status_prv = reg_mstatus_prv;
  assign io_status_sd = T_6433;
  assign io_status_zero3 = reg_mstatus_zero3;
  assign io_status_sd_rv32 = reg_mstatus_sd_rv32;
  assign io_status_zero2 = reg_mstatus_zero2;
  assign io_status_vm = reg_mstatus_vm;
  assign io_status_zero1 = reg_mstatus_zero1;
  assign io_status_pum = reg_mstatus_pum;
  assign io_status_mprv = reg_mstatus_mprv;
  assign io_status_xs = reg_mstatus_xs;
  assign io_status_fs = reg_mstatus_fs;
  assign io_status_mpp = reg_mstatus_mpp;
  assign io_status_hpp = reg_mstatus_hpp;
  assign io_status_spp = reg_mstatus_spp;
  assign io_status_mpie = reg_mstatus_mpie;
  assign io_status_hpie = reg_mstatus_hpie;
  assign io_status_spie = reg_mstatus_spie;
  assign io_status_upie = reg_mstatus_upie;
  assign io_status_mie = reg_mstatus_mie;
  assign io_status_hie = reg_mstatus_hie;
  assign io_status_sie = reg_mstatus_sie;
  assign io_status_uie = reg_mstatus_uie;
  assign io_ptbr = {{12'd0}, reg_sptbr};
  assign io_evec = T_6426;
  assign io_fatc = insn_sfence_vm;
  assign io_time = reg_cycle;
  assign io_fcsr_rm = reg_frm;
  assign io_rocc_cmd_valid = GEN_141;
  assign io_rocc_cmd_bits_inst_funct = GEN_142;
  assign io_rocc_cmd_bits_inst_rs2 = GEN_143;
  assign io_rocc_cmd_bits_inst_rs1 = GEN_144;
  assign io_rocc_cmd_bits_inst_xd = GEN_145;
  assign io_rocc_cmd_bits_inst_xs1 = GEN_146;
  assign io_rocc_cmd_bits_inst_xs2 = GEN_147;
  assign io_rocc_cmd_bits_inst_rd = GEN_148;
  assign io_rocc_cmd_bits_inst_opcode = GEN_149;
  assign io_rocc_cmd_bits_rs1 = GEN_150;
  assign io_rocc_cmd_bits_rs2 = GEN_151;
  assign io_rocc_resp_ready = GEN_152;
  assign io_rocc_mem_req_ready = GEN_153;
  assign io_rocc_mem_s2_nack = GEN_154;
  assign io_rocc_mem_resp_valid = GEN_155;
  assign io_rocc_mem_resp_bits_addr = GEN_156;
  assign io_rocc_mem_resp_bits_tag = GEN_157;
  assign io_rocc_mem_resp_bits_cmd = GEN_158;
  assign io_rocc_mem_resp_bits_typ = GEN_159;
  assign io_rocc_mem_resp_bits_data = GEN_160;
  assign io_rocc_mem_resp_bits_replay = GEN_161;
  assign io_rocc_mem_resp_bits_has_data = GEN_162;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_163;
  assign io_rocc_mem_resp_bits_store_data = GEN_164;
  assign io_rocc_mem_replay_next = GEN_175;
  assign io_rocc_mem_xcpt_ma_ld = GEN_176;
  assign io_rocc_mem_xcpt_ma_st = GEN_177;
  assign io_rocc_mem_xcpt_pf_ld = GEN_178;
  assign io_rocc_mem_xcpt_pf_st = GEN_179;
  assign io_rocc_mem_ordered = GEN_180;
  assign io_rocc_status_debug = GEN_181;
  assign io_rocc_status_prv = GEN_182;
  assign io_rocc_status_sd = GEN_183;
  assign io_rocc_status_zero3 = GEN_184;
  assign io_rocc_status_sd_rv32 = GEN_185;
  assign io_rocc_status_zero2 = GEN_186;
  assign io_rocc_status_vm = GEN_187;
  assign io_rocc_status_zero1 = GEN_200;
  assign io_rocc_status_pum = GEN_201;
  assign io_rocc_status_mprv = GEN_202;
  assign io_rocc_status_xs = GEN_203;
  assign io_rocc_status_fs = GEN_204;
  assign io_rocc_status_mpp = GEN_205;
  assign io_rocc_status_hpp = GEN_206;
  assign io_rocc_status_spp = GEN_207;
  assign io_rocc_status_mpie = GEN_208;
  assign io_rocc_status_hpie = GEN_209;
  assign io_rocc_status_spie = GEN_210;
  assign io_rocc_status_upie = GEN_211;
  assign io_rocc_status_mie = GEN_212;
  assign io_rocc_status_hie = GEN_213;
  assign io_rocc_status_sie = GEN_214;
  assign io_rocc_status_uie = GEN_215;
  assign io_rocc_autl_acquire_ready = GEN_216;
  assign io_rocc_autl_grant_valid = GEN_224;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_225;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_226;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_227;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_228;
  assign io_rocc_autl_grant_bits_g_type = GEN_229;
  assign io_rocc_autl_grant_bits_data = GEN_230;
  assign io_rocc_fpu_req_ready = GEN_231;
  assign io_rocc_fpu_resp_valid = GEN_232;
  assign io_rocc_fpu_resp_bits_data = GEN_233;
  assign io_rocc_fpu_resp_bits_exc = GEN_234;
  assign io_rocc_exception = GEN_235;
  assign io_rocc_csr_waddr = io_rw_addr;
  assign io_rocc_csr_wdata = wdata;
  assign io_rocc_csr_wen = wen;
  assign io_rocc_host_id = GEN_236;
  assign io_interrupt = GEN_63;
  assign io_interrupt_cause = GEN_64;
  assign io_bp_0_control_tdrtype = reg_bp_0_control_tdrtype;
  assign io_bp_0_control_bpamaskmax = reg_bp_0_control_bpamaskmax;
  assign io_bp_0_control_reserved = reg_bp_0_control_reserved;
  assign io_bp_0_control_bpaction = reg_bp_0_control_bpaction;
  assign io_bp_0_control_bpmatch = reg_bp_0_control_bpmatch;
  assign io_bp_0_control_m = reg_bp_0_control_m;
  assign io_bp_0_control_h = reg_bp_0_control_h;
  assign io_bp_0_control_s = reg_bp_0_control_s;
  assign io_bp_0_control_u = reg_bp_0_control_u;
  assign io_bp_0_control_r = reg_bp_0_control_r;
  assign io_bp_0_control_w = reg_bp_0_control_w;
  assign io_bp_0_control_x = reg_bp_0_control_x;
  assign io_bp_0_address = reg_bp_0_address;
  assign T_4951_debug = T_4999;
  assign T_4951_prv = T_4998;
  assign T_4951_sd = T_4997;
  assign T_4951_zero3 = T_4996;
  assign T_4951_sd_rv32 = T_4995;
  assign T_4951_zero2 = T_4994;
  assign T_4951_vm = T_4993;
  assign T_4951_zero1 = T_4992;
  assign T_4951_pum = T_4991;
  assign T_4951_mprv = T_4990;
  assign T_4951_xs = T_4989;
  assign T_4951_fs = T_4988;
  assign T_4951_mpp = T_4987;
  assign T_4951_hpp = T_4986;
  assign T_4951_spp = T_4985;
  assign T_4951_mpie = T_4984;
  assign T_4951_hpie = T_4983;
  assign T_4951_spie = T_4982;
  assign T_4951_upie = T_4981;
  assign T_4951_mie = T_4980;
  assign T_4951_hie = T_4979;
  assign T_4951_sie = T_4978;
  assign T_4951_uie = T_4977;
  assign T_4976 = {{66'd0}, 1'h0};
  assign T_4977 = T_4976[0];
  assign T_4978 = T_4976[1];
  assign T_4979 = T_4976[2];
  assign T_4980 = T_4976[3];
  assign T_4981 = T_4976[4];
  assign T_4982 = T_4976[5];
  assign T_4983 = T_4976[6];
  assign T_4984 = T_4976[7];
  assign T_4985 = T_4976[8];
  assign T_4986 = T_4976[10:9];
  assign T_4987 = T_4976[12:11];
  assign T_4988 = T_4976[14:13];
  assign T_4989 = T_4976[16:15];
  assign T_4990 = T_4976[17];
  assign T_4991 = T_4976[18];
  assign T_4992 = T_4976[23:19];
  assign T_4993 = T_4976[28:24];
  assign T_4994 = T_4976[30:29];
  assign T_4995 = T_4976[31];
  assign T_4996 = T_4976[62:32];
  assign T_4997 = T_4976[63];
  assign T_4998 = T_4976[65:64];
  assign T_4999 = T_4976[66];
  assign reset_mstatus_debug = T_4951_debug;
  assign reset_mstatus_prv = 2'h3;
  assign reset_mstatus_sd = T_4951_sd;
  assign reset_mstatus_zero3 = T_4951_zero3;
  assign reset_mstatus_sd_rv32 = T_4951_sd_rv32;
  assign reset_mstatus_zero2 = T_4951_zero2;
  assign reset_mstatus_vm = T_4951_vm;
  assign reset_mstatus_zero1 = T_4951_zero1;
  assign reset_mstatus_pum = T_4951_pum;
  assign reset_mstatus_mprv = T_4951_mprv;
  assign reset_mstatus_xs = T_4951_xs;
  assign reset_mstatus_fs = T_4951_fs;
  assign reset_mstatus_mpp = 2'h3;
  assign reset_mstatus_hpp = T_4951_hpp;
  assign reset_mstatus_spp = T_4951_spp;
  assign reset_mstatus_mpie = T_4951_mpie;
  assign reset_mstatus_hpie = T_4951_hpie;
  assign reset_mstatus_spie = T_4951_spie;
  assign reset_mstatus_upie = T_4951_upie;
  assign reset_mstatus_mie = T_4951_mie;
  assign reset_mstatus_hie = T_4951_hie;
  assign reset_mstatus_sie = T_4951_sie;
  assign reset_mstatus_uie = T_4951_uie;
  assign T_5085_xdebugver = T_5121;
  assign T_5085_ndreset = T_5120;
  assign T_5085_fullreset = T_5119;
  assign T_5085_hwbpcount = T_5118;
  assign T_5085_ebreakm = T_5117;
  assign T_5085_ebreakh = T_5116;
  assign T_5085_ebreaks = T_5115;
  assign T_5085_ebreaku = T_5114;
  assign T_5085_zero2 = T_5113;
  assign T_5085_stopcycle = T_5112;
  assign T_5085_stoptime = T_5111;
  assign T_5085_cause = T_5110;
  assign T_5085_debugint = T_5109;
  assign T_5085_zero1 = T_5108;
  assign T_5085_halt = T_5107;
  assign T_5085_step = T_5106;
  assign T_5085_prv = T_5105;
  assign T_5104 = {{31'd0}, 1'h0};
  assign T_5105 = T_5104[1:0];
  assign T_5106 = T_5104[2];
  assign T_5107 = T_5104[3];
  assign T_5108 = T_5104[4];
  assign T_5109 = T_5104[5];
  assign T_5110 = T_5104[8:6];
  assign T_5111 = T_5104[9];
  assign T_5112 = T_5104[10];
  assign T_5113 = T_5104[11];
  assign T_5114 = T_5104[12];
  assign T_5115 = T_5104[13];
  assign T_5116 = T_5104[14];
  assign T_5117 = T_5104[15];
  assign T_5118 = T_5104[27:16];
  assign T_5119 = T_5104[28];
  assign T_5120 = T_5104[29];
  assign T_5121 = T_5104[31:30];
  assign reset_dcsr_xdebugver = {{1'd0}, 1'h1};
  assign reset_dcsr_ndreset = T_5085_ndreset;
  assign reset_dcsr_fullreset = T_5085_fullreset;
  assign reset_dcsr_hwbpcount = T_5085_hwbpcount;
  assign reset_dcsr_ebreakm = T_5085_ebreakm;
  assign reset_dcsr_ebreakh = T_5085_ebreakh;
  assign reset_dcsr_ebreaks = T_5085_ebreaks;
  assign reset_dcsr_ebreaku = T_5085_ebreaku;
  assign reset_dcsr_zero2 = T_5085_zero2;
  assign reset_dcsr_stopcycle = T_5085_stopcycle;
  assign reset_dcsr_stoptime = T_5085_stoptime;
  assign reset_dcsr_cause = T_5085_cause;
  assign reset_dcsr_debugint = T_5085_debugint;
  assign reset_dcsr_zero1 = T_5085_zero1;
  assign reset_dcsr_halt = T_5085_halt;
  assign reset_dcsr_step = T_5085_step;
  assign reset_dcsr_prv = 2'h3;
  assign T_5187_rocc = T_5215;
  assign T_5187_meip = T_5214;
  assign T_5187_heip = T_5213;
  assign T_5187_seip = T_5212;
  assign T_5187_ueip = T_5211;
  assign T_5187_mtip = T_5210;
  assign T_5187_htip = T_5209;
  assign T_5187_stip = T_5208;
  assign T_5187_utip = T_5207;
  assign T_5187_msip = T_5206;
  assign T_5187_hsip = T_5205;
  assign T_5187_ssip = T_5204;
  assign T_5187_usip = T_5203;
  assign T_5202 = {{12'd0}, 1'h0};
  assign T_5203 = T_5202[0];
  assign T_5204 = T_5202[1];
  assign T_5205 = T_5202[2];
  assign T_5206 = T_5202[3];
  assign T_5207 = T_5202[4];
  assign T_5208 = T_5202[5];
  assign T_5209 = T_5202[6];
  assign T_5210 = T_5202[7];
  assign T_5211 = T_5202[8];
  assign T_5212 = T_5202[9];
  assign T_5213 = T_5202[10];
  assign T_5214 = T_5202[11];
  assign T_5215 = T_5202[12];
  assign T_5216_rocc = 1'h0;
  assign T_5216_meip = 1'h1;
  assign T_5216_heip = T_5187_heip;
  assign T_5216_seip = 1'h1;
  assign T_5216_ueip = T_5187_ueip;
  assign T_5216_mtip = 1'h1;
  assign T_5216_htip = T_5187_htip;
  assign T_5216_stip = 1'h1;
  assign T_5216_utip = T_5187_utip;
  assign T_5216_msip = 1'h1;
  assign T_5216_hsip = T_5187_hsip;
  assign T_5216_ssip = 1'h1;
  assign T_5216_usip = T_5187_usip;
  assign T_5237_rocc = T_5216_rocc;
  assign T_5237_meip = 1'h0;
  assign T_5237_heip = T_5216_heip;
  assign T_5237_seip = T_5216_seip;
  assign T_5237_ueip = T_5216_ueip;
  assign T_5237_mtip = 1'h0;
  assign T_5237_htip = T_5216_htip;
  assign T_5237_stip = T_5216_stip;
  assign T_5237_utip = T_5216_utip;
  assign T_5237_msip = 1'h0;
  assign T_5237_hsip = T_5216_hsip;
  assign T_5237_ssip = T_5216_ssip;
  assign T_5237_usip = T_5216_usip;
  assign T_5254 = {T_5216_hsip,T_5216_ssip};
  assign T_5255 = {T_5254,T_5216_usip};
  assign T_5256 = {T_5216_stip,T_5216_utip};
  assign T_5257 = {T_5256,T_5216_msip};
  assign T_5258 = {T_5257,T_5255};
  assign T_5259 = {T_5216_ueip,T_5216_mtip};
  assign T_5260 = {T_5259,T_5216_htip};
  assign T_5261 = {T_5216_heip,T_5216_seip};
  assign T_5262 = {T_5216_rocc,T_5216_meip};
  assign T_5263 = {T_5262,T_5261};
  assign T_5264 = {T_5263,T_5260};
  assign supported_interrupts = {T_5264,T_5258};
  assign T_5265 = {T_5237_hsip,T_5237_ssip};
  assign T_5266 = {T_5265,T_5237_usip};
  assign T_5267 = {T_5237_stip,T_5237_utip};
  assign T_5268 = {T_5267,T_5237_msip};
  assign T_5269 = {T_5268,T_5266};
  assign T_5270 = {T_5237_ueip,T_5237_mtip};
  assign T_5271 = {T_5270,T_5237_htip};
  assign T_5272 = {T_5237_heip,T_5237_seip};
  assign T_5273 = {T_5237_rocc,T_5237_meip};
  assign T_5274 = {T_5273,T_5272};
  assign T_5275 = {T_5274,T_5271};
  assign delegable_interrupts = {T_5275,T_5269};
  assign GEN_597 = {{1'd0}, T_5476};
  assign T_5480 = GEN_597 + 7'h1;
  assign T_5481 = T_5480[6:0];
  assign T_5482 = T_5481[5:0];
  assign GEN_27 = io_uarch_counters_0 ? T_5482 : T_5476;
  assign T_5485 = T_5481[6];
  assign T_5486 = io_uarch_counters_0 & T_5485;
  assign GEN_598 = {{57'd0}, 1'h1};
  assign T_5488 = T_5484 + GEN_598;
  assign T_5489 = T_5488[57:0];
  assign GEN_28 = T_5486 ? T_5489 : T_5484;
  assign GEN_599 = {{1'd0}, T_5492};
  assign T_5496 = GEN_599 + 7'h1;
  assign T_5497 = T_5496[6:0];
  assign T_5498 = T_5497[5:0];
  assign GEN_29 = io_uarch_counters_1 ? T_5498 : T_5492;
  assign T_5501 = T_5497[6];
  assign T_5502 = io_uarch_counters_1 & T_5501;
  assign T_5504 = T_5500 + GEN_598;
  assign T_5505 = T_5504[57:0];
  assign GEN_30 = T_5502 ? T_5505 : T_5500;
  assign GEN_601 = {{1'd0}, T_5508};
  assign T_5512 = GEN_601 + 7'h1;
  assign T_5513 = T_5512[6:0];
  assign T_5514 = T_5513[5:0];
  assign GEN_31 = io_uarch_counters_2 ? T_5514 : T_5508;
  assign T_5517 = T_5513[6];
  assign T_5518 = io_uarch_counters_2 & T_5517;
  assign T_5520 = T_5516 + GEN_598;
  assign T_5521 = T_5520[57:0];
  assign GEN_32 = T_5518 ? T_5521 : T_5516;
  assign GEN_603 = {{1'd0}, T_5524};
  assign T_5528 = GEN_603 + 7'h1;
  assign T_5529 = T_5528[6:0];
  assign T_5530 = T_5529[5:0];
  assign GEN_33 = io_uarch_counters_3 ? T_5530 : T_5524;
  assign T_5533 = T_5529[6];
  assign T_5534 = io_uarch_counters_3 & T_5533;
  assign T_5536 = T_5532 + GEN_598;
  assign T_5537 = T_5536[57:0];
  assign GEN_34 = T_5534 ? T_5537 : T_5532;
  assign GEN_605 = {{1'd0}, T_5540};
  assign T_5544 = GEN_605 + 7'h1;
  assign T_5545 = T_5544[6:0];
  assign T_5546 = T_5545[5:0];
  assign GEN_35 = io_uarch_counters_4 ? T_5546 : T_5540;
  assign T_5549 = T_5545[6];
  assign T_5550 = io_uarch_counters_4 & T_5549;
  assign T_5552 = T_5548 + GEN_598;
  assign T_5553 = T_5552[57:0];
  assign GEN_36 = T_5550 ? T_5553 : T_5548;
  assign GEN_607 = {{1'd0}, T_5556};
  assign T_5560 = GEN_607 + 7'h1;
  assign T_5561 = T_5560[6:0];
  assign T_5562 = T_5561[5:0];
  assign GEN_37 = io_uarch_counters_5 ? T_5562 : T_5556;
  assign T_5565 = T_5561[6];
  assign T_5566 = io_uarch_counters_5 & T_5565;
  assign T_5568 = T_5564 + GEN_598;
  assign T_5569 = T_5568[57:0];
  assign GEN_38 = T_5566 ? T_5569 : T_5564;
  assign GEN_609 = {{1'd0}, T_5572};
  assign T_5576 = GEN_609 + 7'h1;
  assign T_5577 = T_5576[6:0];
  assign T_5578 = T_5577[5:0];
  assign GEN_39 = io_uarch_counters_6 ? T_5578 : T_5572;
  assign T_5581 = T_5577[6];
  assign T_5582 = io_uarch_counters_6 & T_5581;
  assign T_5584 = T_5580 + GEN_598;
  assign T_5585 = T_5584[57:0];
  assign GEN_40 = T_5582 ? T_5585 : T_5580;
  assign GEN_611 = {{1'd0}, T_5588};
  assign T_5592 = GEN_611 + 7'h1;
  assign T_5593 = T_5592[6:0];
  assign T_5594 = T_5593[5:0];
  assign GEN_41 = io_uarch_counters_7 ? T_5594 : T_5588;
  assign T_5597 = T_5593[6];
  assign T_5598 = io_uarch_counters_7 & T_5597;
  assign T_5600 = T_5596 + GEN_598;
  assign T_5601 = T_5600[57:0];
  assign GEN_42 = T_5598 ? T_5601 : T_5596;
  assign GEN_613 = {{1'd0}, T_5604};
  assign T_5608 = GEN_613 + 7'h1;
  assign T_5609 = T_5608[6:0];
  assign T_5610 = T_5609[5:0];
  assign GEN_43 = io_uarch_counters_8 ? T_5610 : T_5604;
  assign T_5613 = T_5609[6];
  assign T_5614 = io_uarch_counters_8 & T_5613;
  assign T_5616 = T_5612 + GEN_598;
  assign T_5617 = T_5616[57:0];
  assign GEN_44 = T_5614 ? T_5617 : T_5612;
  assign GEN_615 = {{1'd0}, T_5620};
  assign T_5624 = GEN_615 + 7'h1;
  assign T_5625 = T_5624[6:0];
  assign T_5626 = T_5625[5:0];
  assign GEN_45 = io_uarch_counters_9 ? T_5626 : T_5620;
  assign T_5629 = T_5625[6];
  assign T_5630 = io_uarch_counters_9 & T_5629;
  assign T_5632 = T_5628 + GEN_598;
  assign T_5633 = T_5632[57:0];
  assign GEN_46 = T_5630 ? T_5633 : T_5628;
  assign GEN_617 = {{1'd0}, T_5636};
  assign T_5640 = GEN_617 + 7'h1;
  assign T_5641 = T_5640[6:0];
  assign T_5642 = T_5641[5:0];
  assign GEN_47 = io_uarch_counters_10 ? T_5642 : T_5636;
  assign T_5645 = T_5641[6];
  assign T_5646 = io_uarch_counters_10 & T_5645;
  assign T_5648 = T_5644 + GEN_598;
  assign T_5649 = T_5648[57:0];
  assign GEN_48 = T_5646 ? T_5649 : T_5644;
  assign GEN_619 = {{1'd0}, T_5652};
  assign T_5656 = GEN_619 + 7'h1;
  assign T_5657 = T_5656[6:0];
  assign T_5658 = T_5657[5:0];
  assign GEN_49 = io_uarch_counters_11 ? T_5658 : T_5652;
  assign T_5661 = T_5657[6];
  assign T_5662 = io_uarch_counters_11 & T_5661;
  assign T_5664 = T_5660 + GEN_598;
  assign T_5665 = T_5664[57:0];
  assign GEN_50 = T_5662 ? T_5665 : T_5660;
  assign GEN_621 = {{1'd0}, T_5668};
  assign T_5672 = GEN_621 + 7'h1;
  assign T_5673 = T_5672[6:0];
  assign T_5674 = T_5673[5:0];
  assign GEN_51 = io_uarch_counters_12 ? T_5674 : T_5668;
  assign T_5677 = T_5673[6];
  assign T_5678 = io_uarch_counters_12 & T_5677;
  assign T_5680 = T_5676 + GEN_598;
  assign T_5681 = T_5680[57:0];
  assign GEN_52 = T_5678 ? T_5681 : T_5676;
  assign GEN_623 = {{1'd0}, T_5684};
  assign T_5688 = GEN_623 + 7'h1;
  assign T_5689 = T_5688[6:0];
  assign T_5690 = T_5689[5:0];
  assign GEN_53 = io_uarch_counters_13 ? T_5690 : T_5684;
  assign T_5693 = T_5689[6];
  assign T_5694 = io_uarch_counters_13 & T_5693;
  assign T_5696 = T_5692 + GEN_598;
  assign T_5697 = T_5696[57:0];
  assign GEN_54 = T_5694 ? T_5697 : T_5692;
  assign GEN_625 = {{1'd0}, T_5700};
  assign T_5704 = GEN_625 + 7'h1;
  assign T_5705 = T_5704[6:0];
  assign T_5706 = T_5705[5:0];
  assign GEN_55 = io_uarch_counters_14 ? T_5706 : T_5700;
  assign T_5709 = T_5705[6];
  assign T_5710 = io_uarch_counters_14 & T_5709;
  assign T_5712 = T_5708 + GEN_598;
  assign T_5713 = T_5712[57:0];
  assign GEN_56 = T_5710 ? T_5713 : T_5708;
  assign GEN_627 = {{1'd0}, T_5716};
  assign T_5720 = GEN_627 + 7'h1;
  assign T_5721 = T_5720[6:0];
  assign T_5722 = T_5721[5:0];
  assign GEN_57 = io_uarch_counters_15 ? T_5722 : T_5716;
  assign T_5725 = T_5721[6];
  assign T_5726 = io_uarch_counters_15 & T_5725;
  assign T_5728 = T_5724 + GEN_598;
  assign T_5729 = T_5728[57:0];
  assign GEN_58 = T_5726 ? T_5729 : T_5724;
  assign GEN_629 = {{1'd0}, T_5734};
  assign T_5738 = GEN_629 + 7'h1;
  assign T_5739 = T_5738[6:0];
  assign T_5740 = T_5739[5:0];
  assign GEN_59 = io_retire ? T_5740 : T_5734;
  assign T_5743 = T_5739[6];
  assign T_5744 = io_retire & T_5743;
  assign T_5746 = T_5742 + GEN_598;
  assign T_5747 = T_5746[57:0];
  assign GEN_60 = T_5744 ? T_5747 : T_5742;
  assign T_5748 = {T_5742,T_5734};
  assign GEN_631 = {{1'd0}, T_5751};
  assign T_5755 = GEN_631 + 7'h1;
  assign T_5756 = T_5755[6:0];
  assign T_5757 = T_5756[5:0];
  assign T_5760 = T_5756[6];
  assign T_5763 = T_5759 + GEN_598;
  assign T_5764 = T_5763[57:0];
  assign GEN_62 = T_5760 ? T_5764 : T_5759;
  assign reg_cycle = {T_5759,T_5751};
  assign mip_rocc = io_rocc_interrupt;
  assign mip_meip = reg_mip_meip;
  assign mip_heip = reg_mip_heip;
  assign mip_seip = reg_mip_seip;
  assign mip_ueip = reg_mip_ueip;
  assign mip_mtip = reg_mip_mtip;
  assign mip_htip = reg_mip_htip;
  assign mip_stip = reg_mip_stip;
  assign mip_utip = reg_mip_utip;
  assign mip_msip = reg_mip_msip;
  assign mip_hsip = reg_mip_hsip;
  assign mip_ssip = reg_mip_ssip;
  assign mip_usip = reg_mip_usip;
  assign T_5778 = {mip_hsip,mip_ssip};
  assign T_5779 = {T_5778,mip_usip};
  assign T_5780 = {mip_stip,mip_utip};
  assign T_5781 = {T_5780,mip_msip};
  assign T_5782 = {T_5781,T_5779};
  assign T_5783 = {mip_ueip,mip_mtip};
  assign T_5784 = {T_5783,mip_htip};
  assign T_5785 = {mip_heip,mip_seip};
  assign T_5786 = {mip_rocc,mip_meip};
  assign T_5787 = {T_5786,T_5785};
  assign T_5788 = {T_5787,T_5784};
  assign T_5789 = {T_5788,T_5782};
  assign read_mip = T_5789 & supported_interrupts;
  assign GEN_633 = {{51'd0}, read_mip};
  assign pending_interrupts = GEN_633 & reg_mie;
  assign T_5791 = reg_debug == 1'h0;
  assign T_5793 = reg_mstatus_prv < 2'h3;
  assign T_5795 = reg_mstatus_prv == 2'h3;
  assign T_5796 = T_5795 & reg_mstatus_mie;
  assign T_5797 = T_5793 | T_5796;
  assign T_5798 = T_5791 & T_5797;
  assign T_5799 = ~ reg_mideleg;
  assign T_5800 = pending_interrupts & T_5799;
  assign m_interrupts = T_5798 ? T_5800 : {{63'd0}, 1'h0};
  assign GEN_634 = {{1'd0}, 1'h1};
  assign T_5805 = reg_mstatus_prv < GEN_634;
  assign T_5807 = reg_mstatus_prv == GEN_634;
  assign T_5808 = T_5807 & reg_mstatus_sie;
  assign T_5809 = T_5805 | T_5808;
  assign T_5810 = T_5791 & T_5809;
  assign T_5811 = pending_interrupts & reg_mideleg;
  assign s_interrupts = T_5810 ? T_5811 : {{63'd0}, 1'h0};
  assign all_interrupts = m_interrupts | s_interrupts;
  assign T_5814 = all_interrupts[0];
  assign T_5815 = all_interrupts[1];
  assign T_5816 = all_interrupts[2];
  assign T_5817 = all_interrupts[3];
  assign T_5818 = all_interrupts[4];
  assign T_5819 = all_interrupts[5];
  assign T_5820 = all_interrupts[6];
  assign T_5821 = all_interrupts[7];
  assign T_5822 = all_interrupts[8];
  assign T_5823 = all_interrupts[9];
  assign T_5824 = all_interrupts[10];
  assign T_5825 = all_interrupts[11];
  assign T_5826 = all_interrupts[12];
  assign T_5827 = all_interrupts[13];
  assign T_5828 = all_interrupts[14];
  assign T_5829 = all_interrupts[15];
  assign T_5830 = all_interrupts[16];
  assign T_5831 = all_interrupts[17];
  assign T_5832 = all_interrupts[18];
  assign T_5833 = all_interrupts[19];
  assign T_5834 = all_interrupts[20];
  assign T_5835 = all_interrupts[21];
  assign T_5836 = all_interrupts[22];
  assign T_5837 = all_interrupts[23];
  assign T_5838 = all_interrupts[24];
  assign T_5839 = all_interrupts[25];
  assign T_5840 = all_interrupts[26];
  assign T_5841 = all_interrupts[27];
  assign T_5842 = all_interrupts[28];
  assign T_5843 = all_interrupts[29];
  assign T_5844 = all_interrupts[30];
  assign T_5845 = all_interrupts[31];
  assign T_5846 = all_interrupts[32];
  assign T_5847 = all_interrupts[33];
  assign T_5848 = all_interrupts[34];
  assign T_5849 = all_interrupts[35];
  assign T_5850 = all_interrupts[36];
  assign T_5851 = all_interrupts[37];
  assign T_5852 = all_interrupts[38];
  assign T_5853 = all_interrupts[39];
  assign T_5854 = all_interrupts[40];
  assign T_5855 = all_interrupts[41];
  assign T_5856 = all_interrupts[42];
  assign T_5857 = all_interrupts[43];
  assign T_5858 = all_interrupts[44];
  assign T_5859 = all_interrupts[45];
  assign T_5860 = all_interrupts[46];
  assign T_5861 = all_interrupts[47];
  assign T_5862 = all_interrupts[48];
  assign T_5863 = all_interrupts[49];
  assign T_5864 = all_interrupts[50];
  assign T_5865 = all_interrupts[51];
  assign T_5866 = all_interrupts[52];
  assign T_5867 = all_interrupts[53];
  assign T_5868 = all_interrupts[54];
  assign T_5869 = all_interrupts[55];
  assign T_5870 = all_interrupts[56];
  assign T_5871 = all_interrupts[57];
  assign T_5872 = all_interrupts[58];
  assign T_5873 = all_interrupts[59];
  assign T_5874 = all_interrupts[60];
  assign T_5875 = all_interrupts[61];
  assign T_5876 = all_interrupts[62];
  assign T_5942 = T_5876 ? 6'h3e : 6'h3f;
  assign T_5943 = T_5875 ? 6'h3d : T_5942;
  assign T_5944 = T_5874 ? 6'h3c : T_5943;
  assign T_5945 = T_5873 ? 6'h3b : T_5944;
  assign T_5946 = T_5872 ? 6'h3a : T_5945;
  assign T_5947 = T_5871 ? 6'h39 : T_5946;
  assign T_5948 = T_5870 ? 6'h38 : T_5947;
  assign T_5949 = T_5869 ? 6'h37 : T_5948;
  assign T_5950 = T_5868 ? 6'h36 : T_5949;
  assign T_5951 = T_5867 ? 6'h35 : T_5950;
  assign T_5952 = T_5866 ? 6'h34 : T_5951;
  assign T_5953 = T_5865 ? 6'h33 : T_5952;
  assign T_5954 = T_5864 ? 6'h32 : T_5953;
  assign T_5955 = T_5863 ? 6'h31 : T_5954;
  assign T_5956 = T_5862 ? 6'h30 : T_5955;
  assign T_5957 = T_5861 ? 6'h2f : T_5956;
  assign T_5958 = T_5860 ? 6'h2e : T_5957;
  assign T_5959 = T_5859 ? 6'h2d : T_5958;
  assign T_5960 = T_5858 ? 6'h2c : T_5959;
  assign T_5961 = T_5857 ? 6'h2b : T_5960;
  assign T_5962 = T_5856 ? 6'h2a : T_5961;
  assign T_5963 = T_5855 ? 6'h29 : T_5962;
  assign T_5964 = T_5854 ? 6'h28 : T_5963;
  assign T_5965 = T_5853 ? 6'h27 : T_5964;
  assign T_5966 = T_5852 ? 6'h26 : T_5965;
  assign T_5967 = T_5851 ? 6'h25 : T_5966;
  assign T_5968 = T_5850 ? 6'h24 : T_5967;
  assign T_5969 = T_5849 ? 6'h23 : T_5968;
  assign T_5970 = T_5848 ? 6'h22 : T_5969;
  assign T_5971 = T_5847 ? 6'h21 : T_5970;
  assign T_5972 = T_5846 ? 6'h20 : T_5971;
  assign T_5973 = T_5845 ? {{1'd0}, 5'h1f} : T_5972;
  assign T_5974 = T_5844 ? {{1'd0}, 5'h1e} : T_5973;
  assign T_5975 = T_5843 ? {{1'd0}, 5'h1d} : T_5974;
  assign T_5976 = T_5842 ? {{1'd0}, 5'h1c} : T_5975;
  assign T_5977 = T_5841 ? {{1'd0}, 5'h1b} : T_5976;
  assign T_5978 = T_5840 ? {{1'd0}, 5'h1a} : T_5977;
  assign T_5979 = T_5839 ? {{1'd0}, 5'h19} : T_5978;
  assign T_5980 = T_5838 ? {{1'd0}, 5'h18} : T_5979;
  assign T_5981 = T_5837 ? {{1'd0}, 5'h17} : T_5980;
  assign T_5982 = T_5836 ? {{1'd0}, 5'h16} : T_5981;
  assign T_5983 = T_5835 ? {{1'd0}, 5'h15} : T_5982;
  assign T_5984 = T_5834 ? {{1'd0}, 5'h14} : T_5983;
  assign T_5985 = T_5833 ? {{1'd0}, 5'h13} : T_5984;
  assign T_5986 = T_5832 ? {{1'd0}, 5'h12} : T_5985;
  assign T_5987 = T_5831 ? {{1'd0}, 5'h11} : T_5986;
  assign T_5988 = T_5830 ? {{1'd0}, 5'h10} : T_5987;
  assign T_5989 = T_5829 ? {{2'd0}, 4'hf} : T_5988;
  assign T_5990 = T_5828 ? {{2'd0}, 4'he} : T_5989;
  assign T_5991 = T_5827 ? {{2'd0}, 4'hd} : T_5990;
  assign T_5992 = T_5826 ? {{2'd0}, 4'hc} : T_5991;
  assign T_5993 = T_5825 ? {{2'd0}, 4'hb} : T_5992;
  assign T_5994 = T_5824 ? {{2'd0}, 4'ha} : T_5993;
  assign T_5995 = T_5823 ? {{2'd0}, 4'h9} : T_5994;
  assign T_5996 = T_5822 ? {{2'd0}, 4'h8} : T_5995;
  assign T_5997 = T_5821 ? {{3'd0}, 3'h7} : T_5996;
  assign T_5998 = T_5820 ? {{3'd0}, 3'h6} : T_5997;
  assign T_5999 = T_5819 ? {{3'd0}, 3'h5} : T_5998;
  assign T_6000 = T_5818 ? {{3'd0}, 3'h4} : T_5999;
  assign T_6001 = T_5817 ? {{4'd0}, 2'h3} : T_6000;
  assign T_6002 = T_5816 ? {{4'd0}, 2'h2} : T_6001;
  assign T_6003 = T_5815 ? {{5'd0}, 1'h1} : T_6002;
  assign T_6004 = T_5814 ? {{5'd0}, 1'h0} : T_6003;
  assign GEN_636 = {{58'd0}, T_6004};
  assign T_6005 = 64'h8000000000000000 + GEN_636;
  assign interruptCause = T_6005[63:0];
  assign GEN_637 = {{63'd0}, 1'h0};
  assign T_6007 = all_interrupts != GEN_637;
  assign T_6012 = reg_dcsr_debugint & T_5791;
  assign GEN_63 = T_6012 ? 1'h1 : T_6007;
  assign GEN_64 = T_6012 ? 64'h800000000000000d : interruptCause;
  assign system_insn = io_rw_cmd == 3'h4;
  assign T_6015 = io_rw_cmd != 3'h0;
  assign T_6017 = system_insn == 1'h0;
  assign cpu_ren = T_6015 & T_6017;
  assign T_6018 = {io_status_sie,io_status_uie};
  assign T_6019 = {io_status_upie,io_status_mie};
  assign T_6020 = {T_6019,io_status_hie};
  assign T_6021 = {T_6020,T_6018};
  assign T_6022 = {io_status_mpie,io_status_hpie};
  assign T_6023 = {T_6022,io_status_spie};
  assign T_6024 = {io_status_mpp,io_status_hpp};
  assign T_6025 = {T_6024,io_status_spp};
  assign T_6026 = {T_6025,T_6023};
  assign T_6027 = {T_6026,T_6021};
  assign T_6028 = {io_status_mprv,io_status_xs};
  assign T_6029 = {T_6028,io_status_fs};
  assign T_6030 = {io_status_vm,io_status_zero1};
  assign T_6031 = {T_6030,io_status_pum};
  assign T_6032 = {T_6031,T_6029};
  assign T_6033 = {io_status_zero3,io_status_sd_rv32};
  assign T_6034 = {T_6033,io_status_zero2};
  assign T_6035 = {io_status_debug,io_status_prv};
  assign T_6036 = {T_6035,io_status_sd};
  assign T_6037 = {T_6036,T_6034};
  assign T_6038 = {T_6037,T_6032};
  assign T_6039 = {T_6038,T_6027};
  assign read_mstatus = T_6039[63:0];
  assign T_6040 = {reg_tdrselect_tdrmode,reg_tdrselect_reserved};
  assign T_6041 = {T_6040,reg_tdrselect_tdrindex};
  assign GEN_0 = GEN_65;
  assign GEN_65 = reg_tdrselect_tdrindex ? reg_bp_1_control_r : reg_bp_0_control_r;
  assign GEN_1 = GEN_66;
  assign GEN_66 = reg_tdrselect_tdrindex ? reg_bp_1_control_w : reg_bp_0_control_w;
  assign T_6056 = {GEN_0,GEN_1};
  assign GEN_2 = GEN_67;
  assign GEN_67 = reg_tdrselect_tdrindex ? reg_bp_1_control_x : reg_bp_0_control_x;
  assign T_6057 = {T_6056,GEN_2};
  assign GEN_3 = GEN_68;
  assign GEN_68 = reg_tdrselect_tdrindex ? reg_bp_1_control_h : reg_bp_0_control_h;
  assign GEN_4 = GEN_69;
  assign GEN_69 = reg_tdrselect_tdrindex ? reg_bp_1_control_s : reg_bp_0_control_s;
  assign T_6058 = {GEN_3,GEN_4};
  assign GEN_5 = GEN_70;
  assign GEN_70 = reg_tdrselect_tdrindex ? reg_bp_1_control_u : reg_bp_0_control_u;
  assign T_6059 = {T_6058,GEN_5};
  assign T_6060 = {T_6059,T_6057};
  assign GEN_6 = GEN_71;
  assign GEN_71 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpaction : reg_bp_0_control_bpaction;
  assign GEN_7 = GEN_72;
  assign GEN_72 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpmatch : reg_bp_0_control_bpmatch;
  assign T_6061 = {GEN_6,GEN_7};
  assign GEN_8 = GEN_73;
  assign GEN_73 = reg_tdrselect_tdrindex ? reg_bp_1_control_m : reg_bp_0_control_m;
  assign T_6062 = {T_6061,GEN_8};
  assign GEN_9 = GEN_74;
  assign GEN_74 = reg_tdrselect_tdrindex ? reg_bp_1_control_tdrtype : reg_bp_0_control_tdrtype;
  assign GEN_10 = GEN_75;
  assign GEN_75 = reg_tdrselect_tdrindex ? reg_bp_1_control_bpamaskmax : reg_bp_0_control_bpamaskmax;
  assign T_6063 = {GEN_9,GEN_10};
  assign GEN_11 = GEN_76;
  assign GEN_76 = reg_tdrselect_tdrindex ? reg_bp_1_control_reserved : reg_bp_0_control_reserved;
  assign T_6064 = {T_6063,GEN_11};
  assign T_6065 = {T_6064,T_6062};
  assign T_6066 = {T_6065,T_6060};
  assign T_6089 = reg_mepc[39];
  assign GEN_638 = {{23'd0}, T_6089};
  assign T_6091 = 24'h0 - GEN_638;
  assign T_6092 = T_6091[23:0];
  assign T_6093 = {T_6092,reg_mepc};
  assign T_6094 = reg_mbadaddr[39];
  assign GEN_639 = {{23'd0}, T_6094};
  assign T_6096 = 24'h0 - GEN_639;
  assign T_6097 = T_6096[23:0];
  assign T_6098 = {T_6097,reg_mbadaddr};
  assign T_6099 = {reg_dcsr_step,reg_dcsr_prv};
  assign T_6100 = {reg_dcsr_zero1,reg_dcsr_halt};
  assign T_6101 = {T_6100,T_6099};
  assign T_6102 = {reg_dcsr_cause,reg_dcsr_debugint};
  assign T_6103 = {reg_dcsr_stopcycle,reg_dcsr_stoptime};
  assign T_6104 = {T_6103,T_6102};
  assign T_6105 = {T_6104,T_6101};
  assign T_6106 = {reg_dcsr_ebreaku,reg_dcsr_zero2};
  assign T_6107 = {reg_dcsr_ebreakh,reg_dcsr_ebreaks};
  assign T_6108 = {T_6107,T_6106};
  assign T_6109 = {reg_dcsr_hwbpcount,reg_dcsr_ebreakm};
  assign T_6110 = {reg_dcsr_xdebugver,reg_dcsr_ndreset};
  assign T_6111 = {T_6110,reg_dcsr_fullreset};
  assign T_6112 = {T_6111,T_6109};
  assign T_6113 = {T_6112,T_6108};
  assign T_6114 = {T_6113,T_6105};
  assign T_6115 = {reg_frm,reg_fflags};
  assign T_6116 = reg_mie & reg_mideleg;
  assign T_6117 = GEN_633 & reg_mideleg;
  assign T_6118_debug = io_status_debug;
  assign T_6118_prv = io_status_prv;
  assign T_6118_sd = io_status_sd;
  assign T_6118_zero3 = io_status_zero3;
  assign T_6118_sd_rv32 = io_status_sd_rv32;
  assign T_6118_zero2 = io_status_zero2;
  assign T_6118_vm = {{4'd0}, 1'h0};
  assign T_6118_zero1 = io_status_zero1;
  assign T_6118_pum = io_status_pum;
  assign T_6118_mprv = 1'h0;
  assign T_6118_xs = io_status_xs;
  assign T_6118_fs = io_status_fs;
  assign T_6118_mpp = {{1'd0}, 1'h0};
  assign T_6118_hpp = {{1'd0}, 1'h0};
  assign T_6118_spp = io_status_spp;
  assign T_6118_mpie = 1'h0;
  assign T_6118_hpie = 1'h0;
  assign T_6118_spie = io_status_spie;
  assign T_6118_upie = io_status_upie;
  assign T_6118_mie = 1'h0;
  assign T_6118_hie = 1'h0;
  assign T_6118_sie = io_status_sie;
  assign T_6118_uie = io_status_uie;
  assign T_6150 = {T_6118_sie,T_6118_uie};
  assign T_6151 = {T_6118_upie,T_6118_mie};
  assign T_6152 = {T_6151,T_6118_hie};
  assign T_6153 = {T_6152,T_6150};
  assign T_6154 = {T_6118_mpie,T_6118_hpie};
  assign T_6155 = {T_6154,T_6118_spie};
  assign T_6156 = {T_6118_mpp,T_6118_hpp};
  assign T_6157 = {T_6156,T_6118_spp};
  assign T_6158 = {T_6157,T_6155};
  assign T_6159 = {T_6158,T_6153};
  assign T_6160 = {T_6118_mprv,T_6118_xs};
  assign T_6161 = {T_6160,T_6118_fs};
  assign T_6162 = {T_6118_vm,T_6118_zero1};
  assign T_6163 = {T_6162,T_6118_pum};
  assign T_6164 = {T_6163,T_6161};
  assign T_6165 = {T_6118_zero3,T_6118_sd_rv32};
  assign T_6166 = {T_6165,T_6118_zero2};
  assign T_6167 = {T_6118_debug,T_6118_prv};
  assign T_6168 = {T_6167,T_6118_sd};
  assign T_6169 = {T_6168,T_6166};
  assign T_6170 = {T_6169,T_6164};
  assign T_6171 = {T_6170,T_6159};
  assign T_6172 = T_6171[63:0];
  assign T_6173 = reg_sbadaddr[39];
  assign GEN_641 = {{23'd0}, T_6173};
  assign T_6175 = 24'h0 - GEN_641;
  assign T_6176 = T_6175[23:0];
  assign T_6177 = {T_6176,reg_sbadaddr};
  assign T_6179 = reg_sepc[39];
  assign GEN_642 = {{23'd0}, T_6179};
  assign T_6181 = 24'h0 - GEN_642;
  assign T_6182 = T_6181[23:0];
  assign T_6183 = {T_6182,reg_sepc};
  assign T_6184 = reg_stvec[38];
  assign GEN_643 = {{24'd0}, T_6184};
  assign T_6186 = 25'h0 - GEN_643;
  assign T_6187 = T_6186[24:0];
  assign T_6188 = {T_6187,reg_stvec};
  assign GEN_644 = {{1'd0}, 11'h7a0};
  assign T_6194 = io_rw_addr == GEN_644;
  assign GEN_645 = {{1'd0}, 11'h7a1};
  assign T_6196 = io_rw_addr == GEN_645;
  assign GEN_646 = {{1'd0}, 11'h7a2};
  assign T_6198 = io_rw_addr == GEN_646;
  assign T_6200 = io_rw_addr == 12'hf13;
  assign T_6202 = io_rw_addr == 12'hf12;
  assign T_6204 = io_rw_addr == 12'hf11;
  assign T_6206 = io_rw_addr == 12'hf00;
  assign T_6208 = io_rw_addr == 12'hf02;
  assign GEN_647 = {{2'd0}, 10'h310};
  assign T_6210 = io_rw_addr == GEN_647;
  assign GEN_648 = {{1'd0}, 11'h701};
  assign T_6212 = io_rw_addr == GEN_648;
  assign GEN_649 = {{1'd0}, 11'h700};
  assign T_6214 = io_rw_addr == GEN_649;
  assign GEN_650 = {{1'd0}, 11'h702};
  assign T_6216 = io_rw_addr == GEN_650;
  assign T_6218 = io_rw_addr == 12'hf10;
  assign GEN_651 = {{2'd0}, 10'h300};
  assign T_6220 = io_rw_addr == GEN_651;
  assign GEN_652 = {{2'd0}, 10'h305};
  assign T_6222 = io_rw_addr == GEN_652;
  assign GEN_653 = {{2'd0}, 10'h344};
  assign T_6224 = io_rw_addr == GEN_653;
  assign GEN_654 = {{2'd0}, 10'h304};
  assign T_6226 = io_rw_addr == GEN_654;
  assign GEN_655 = {{2'd0}, 10'h303};
  assign T_6228 = io_rw_addr == GEN_655;
  assign GEN_656 = {{2'd0}, 10'h302};
  assign T_6230 = io_rw_addr == GEN_656;
  assign GEN_657 = {{2'd0}, 10'h340};
  assign T_6232 = io_rw_addr == GEN_657;
  assign GEN_658 = {{2'd0}, 10'h341};
  assign T_6234 = io_rw_addr == GEN_658;
  assign GEN_659 = {{2'd0}, 10'h343};
  assign T_6236 = io_rw_addr == GEN_659;
  assign GEN_660 = {{2'd0}, 10'h342};
  assign T_6238 = io_rw_addr == GEN_660;
  assign T_6240 = io_rw_addr == 12'hf14;
  assign GEN_661 = {{1'd0}, 11'h7b0};
  assign T_6242 = io_rw_addr == GEN_661;
  assign GEN_662 = {{1'd0}, 11'h7b1};
  assign T_6244 = io_rw_addr == GEN_662;
  assign GEN_663 = {{1'd0}, 11'h7b2};
  assign T_6246 = io_rw_addr == GEN_663;
  assign GEN_664 = {{11'd0}, 1'h1};
  assign T_6248 = io_rw_addr == GEN_664;
  assign GEN_665 = {{10'd0}, 2'h2};
  assign T_6250 = io_rw_addr == GEN_665;
  assign GEN_666 = {{10'd0}, 2'h3};
  assign T_6252 = io_rw_addr == GEN_666;
  assign GEN_667 = {{3'd0}, 9'h100};
  assign T_6254 = io_rw_addr == GEN_667;
  assign GEN_668 = {{3'd0}, 9'h144};
  assign T_6256 = io_rw_addr == GEN_668;
  assign GEN_669 = {{3'd0}, 9'h104};
  assign T_6258 = io_rw_addr == GEN_669;
  assign GEN_670 = {{3'd0}, 9'h140};
  assign T_6260 = io_rw_addr == GEN_670;
  assign GEN_671 = {{3'd0}, 9'h142};
  assign T_6262 = io_rw_addr == GEN_671;
  assign GEN_672 = {{3'd0}, 9'h143};
  assign T_6264 = io_rw_addr == GEN_672;
  assign GEN_673 = {{3'd0}, 9'h180};
  assign T_6266 = io_rw_addr == GEN_673;
  assign GEN_674 = {{3'd0}, 9'h181};
  assign T_6268 = io_rw_addr == GEN_674;
  assign GEN_675 = {{3'd0}, 9'h141};
  assign T_6270 = io_rw_addr == GEN_675;
  assign GEN_676 = {{3'd0}, 9'h105};
  assign T_6272 = io_rw_addr == GEN_676;
  assign GEN_677 = {{2'd0}, 10'h311};
  assign T_6274 = io_rw_addr == GEN_677;
  assign GEN_678 = {{1'd0}, 11'h705};
  assign T_6276 = io_rw_addr == GEN_678;
  assign GEN_679 = {{1'd0}, 11'h704};
  assign T_6278 = io_rw_addr == GEN_679;
  assign GEN_680 = {{1'd0}, 11'h706};
  assign T_6280 = io_rw_addr == GEN_680;
  assign T_6281 = T_6194 | T_6196;
  assign T_6282 = T_6281 | T_6198;
  assign T_6283 = T_6282 | T_6200;
  assign T_6284 = T_6283 | T_6202;
  assign T_6285 = T_6284 | T_6204;
  assign T_6286 = T_6285 | T_6206;
  assign T_6287 = T_6286 | T_6208;
  assign T_6288 = T_6287 | T_6210;
  assign T_6289 = T_6288 | T_6212;
  assign T_6290 = T_6289 | T_6214;
  assign T_6291 = T_6290 | T_6216;
  assign T_6292 = T_6291 | T_6218;
  assign T_6293 = T_6292 | T_6220;
  assign T_6294 = T_6293 | T_6222;
  assign T_6295 = T_6294 | T_6224;
  assign T_6296 = T_6295 | T_6226;
  assign T_6297 = T_6296 | T_6228;
  assign T_6298 = T_6297 | T_6230;
  assign T_6299 = T_6298 | T_6232;
  assign T_6300 = T_6299 | T_6234;
  assign T_6301 = T_6300 | T_6236;
  assign T_6302 = T_6301 | T_6238;
  assign T_6303 = T_6302 | T_6240;
  assign T_6304 = T_6303 | T_6242;
  assign T_6305 = T_6304 | T_6244;
  assign T_6306 = T_6305 | T_6246;
  assign T_6307 = T_6306 | T_6248;
  assign T_6308 = T_6307 | T_6250;
  assign T_6309 = T_6308 | T_6252;
  assign T_6310 = T_6309 | T_6254;
  assign T_6311 = T_6310 | T_6256;
  assign T_6312 = T_6311 | T_6258;
  assign T_6313 = T_6312 | T_6260;
  assign T_6314 = T_6313 | T_6262;
  assign T_6315 = T_6314 | T_6264;
  assign T_6316 = T_6315 | T_6266;
  assign T_6317 = T_6316 | T_6268;
  assign T_6318 = T_6317 | T_6270;
  assign T_6319 = T_6318 | T_6272;
  assign T_6320 = T_6319 | T_6274;
  assign T_6321 = T_6320 | T_6276;
  assign T_6322 = T_6321 | T_6278;
  assign addr_valid = T_6322 | T_6280;
  assign T_6323 = T_6248 | T_6250;
  assign fp_csr = T_6323 | T_6252;
  assign T_6325 = io_rw_addr[5];
  assign T_6326 = io_rw_addr[6:5];
  assign T_6327 = ~ T_6326;
  assign GEN_681 = {{1'd0}, 1'h0};
  assign T_6329 = T_6327 == GEN_681;
  assign T_6330 = io_rw_addr[9:8];
  assign csr_addr_priv = {T_6329,T_6330};
  assign T_6331 = {reg_debug,reg_mstatus_prv};
  assign priv_sufficient = T_6331 >= csr_addr_priv;
  assign T_6332 = io_rw_addr[11:10];
  assign T_6333 = ~ T_6332;
  assign read_only = T_6333 == GEN_681;
  assign T_6335 = io_rw_cmd != 3'h5;
  assign T_6336 = cpu_ren & T_6335;
  assign cpu_wen = T_6336 & priv_sufficient;
  assign T_6338 = read_only == 1'h0;
  assign wen = cpu_wen & T_6338;
  assign T_6339 = io_rw_cmd == 3'h2;
  assign T_6340 = io_rw_cmd == 3'h3;
  assign T_6341 = T_6339 | T_6340;
  assign T_6343 = T_6341 ? io_rw_rdata : {{63'd0}, 1'h0};
  assign T_6344 = io_rw_cmd != 3'h3;
  assign T_6346 = T_6344 ? io_rw_wdata : {{63'd0}, 1'h0};
  assign T_6347 = T_6343 | T_6346;
  assign T_6350 = T_6340 ? io_rw_wdata : {{63'd0}, 1'h0};
  assign T_6351 = ~ T_6350;
  assign wdata = T_6347 & T_6351;
  assign do_system_insn = priv_sufficient & system_insn;
  assign T_6353 = io_rw_addr[2:0];
  assign GEN_683 = {{7'd0}, 1'h1};
  assign opcode = GEN_683 << T_6353;
  assign T_6354 = opcode[0];
  assign insn_call = do_system_insn & T_6354;
  assign T_6355 = opcode[1];
  assign insn_break = do_system_insn & T_6355;
  assign T_6356 = opcode[2];
  assign insn_ret = do_system_insn & T_6356;
  assign T_6357 = opcode[4];
  assign insn_sfence_vm = do_system_insn & T_6357;
  assign T_6358 = opcode[5];
  assign insn_wfi = do_system_insn & T_6358;
  assign T_6359 = cpu_wen & read_only;
  assign T_6361 = priv_sufficient == 1'h0;
  assign T_6363 = addr_valid == 1'h0;
  assign T_6364 = T_6361 | T_6363;
  assign T_6366 = io_status_fs != GEN_681;
  assign T_6368 = T_6366 == 1'h0;
  assign T_6369 = fp_csr & T_6368;
  assign T_6370 = T_6364 | T_6369;
  assign T_6371 = cpu_ren & T_6370;
  assign T_6372 = T_6359 | T_6371;
  assign T_6375 = system_insn & T_6361;
  assign T_6376 = T_6372 | T_6375;
  assign T_6377 = T_6376 | insn_call;
  assign csr_xcpt = T_6377 | insn_break;
  assign GEN_77 = insn_wfi ? 1'h1 : reg_wfi;
  assign GEN_685 = {{12'd0}, 1'h0};
  assign T_6380 = read_mip != GEN_685;
  assign GEN_78 = T_6380 ? 1'h0 : GEN_77;
  assign T_6383 = csr_xcpt == 1'h0;
  assign GEN_686 = {{2'd0}, reg_mstatus_prv};
  assign T_6385 = GEN_686 + 4'h8;
  assign T_6386 = T_6385[3:0];
  assign T_6389 = insn_break ? 2'h3 : 2'h2;
  assign T_6390 = insn_call ? T_6386 : {{2'd0}, T_6389};
  assign cause = T_6383 ? io_cause : {{60'd0}, T_6390};
  assign cause_lsbs = cause[5:0];
  assign T_6391 = cause[63];
  assign GEN_687 = {{2'd0}, 4'hd};
  assign T_6393 = cause_lsbs == GEN_687;
  assign causeIsDebugInt = T_6391 & T_6393;
  assign GEN_688 = {{62'd0}, 2'h3};
  assign T_6395 = cause == GEN_688;
  assign T_6396 = {reg_dcsr_ebreaks,reg_dcsr_ebreaku};
  assign T_6397 = {reg_dcsr_ebreakm,reg_dcsr_ebreakh};
  assign T_6398 = {T_6397,T_6396};
  assign T_6399 = T_6398 >> reg_mstatus_prv;
  assign T_6400 = T_6399[0];
  assign causeIsDebugBreak = T_6395 & T_6400;
  assign T_6402 = causeIsDebugInt | causeIsDebugBreak;
  assign T_6403 = T_6402 | reg_debug;
  assign T_6409 = reg_mideleg >> cause_lsbs;
  assign T_6410 = T_6409[0];
  assign T_6411 = reg_medeleg >> cause_lsbs;
  assign T_6412 = T_6411[0];
  assign T_6413 = T_6391 ? T_6410 : T_6412;
  assign delegate = T_5793 & T_6413;
  assign debugTVec = reg_debug ? 12'h808 : 12'h800;
  assign T_6417 = {T_6184,reg_stvec};
  assign T_6418 = delegate ? T_6417 : {{8'd0}, reg_mtvec};
  assign tvec = T_6403 ? {{28'd0}, debugTVec} : T_6418;
  assign T_6420 = csr_addr_priv[1];
  assign T_6422 = T_6420 == 1'h0;
  assign T_6424 = T_6422 ? reg_sepc : reg_mepc;
  assign epc = T_6325 ? reg_dpc : T_6424;
  assign T_6425 = io_exception | csr_xcpt;
  assign T_6426 = T_6425 ? tvec : epc;
  assign T_6427 = ~ io_status_fs;
  assign T_6429 = T_6427 == GEN_681;
  assign T_6430 = ~ io_status_xs;
  assign T_6432 = T_6430 == GEN_681;
  assign T_6433 = T_6429 | T_6432;
  assign T_6435 = ~ io_pc;
  assign GEN_691 = {{38'd0}, 2'h3};
  assign T_6437 = T_6435 | GEN_691;
  assign T_6438 = ~ T_6437;
  assign T_6439 = read_mstatus >> reg_mstatus_prv;
  assign T_6440 = T_6439[0];
  assign T_6444 = causeIsDebugInt ? 2'h3 : {{1'd0}, 1'h1};
  assign GEN_79 = T_6403 ? 1'h1 : reg_debug;
  assign GEN_80 = T_6403 ? T_6438 : reg_dpc;
  assign GEN_81 = T_6403 ? {{1'd0}, T_6444} : reg_dcsr_cause;
  assign GEN_82 = T_6403 ? reg_mstatus_prv : reg_dcsr_prv;
  assign T_6446 = T_6403 == 1'h0;
  assign T_6447 = T_6446 & delegate;
  assign GEN_83 = T_6447 ? T_6438 : reg_sepc;
  assign GEN_84 = T_6447 ? cause : reg_scause;
  assign GEN_85 = T_6447 ? io_badaddr : reg_sbadaddr;
  assign GEN_86 = T_6447 ? T_6440 : reg_mstatus_spie;
  assign GEN_87 = T_6447 ? reg_mstatus_prv : {{1'd0}, reg_mstatus_spp};
  assign GEN_88 = T_6447 ? 1'h0 : reg_mstatus_sie;
  assign GEN_89 = T_6447 ? {{1'd0}, 1'h1} : reg_mstatus_prv;
  assign T_6453 = delegate == 1'h0;
  assign T_6454 = T_6446 & T_6453;
  assign GEN_90 = T_6454 ? T_6438 : reg_mepc;
  assign GEN_91 = T_6454 ? cause : reg_mcause;
  assign GEN_92 = T_6454 ? io_badaddr : reg_mbadaddr;
  assign GEN_93 = T_6454 ? T_6440 : reg_mstatus_mpie;
  assign GEN_94 = T_6454 ? reg_mstatus_prv : reg_mstatus_mpp;
  assign GEN_95 = T_6454 ? 1'h0 : reg_mstatus_mie;
  assign GEN_96 = T_6454 ? 2'h3 : GEN_89;
  assign GEN_97 = T_6425 ? GEN_79 : reg_debug;
  assign GEN_98 = T_6425 ? GEN_80 : reg_dpc;
  assign GEN_99 = T_6425 ? GEN_81 : reg_dcsr_cause;
  assign GEN_100 = T_6425 ? GEN_82 : reg_dcsr_prv;
  assign GEN_101 = T_6425 ? GEN_83 : reg_sepc;
  assign GEN_102 = T_6425 ? GEN_84 : reg_scause;
  assign GEN_103 = T_6425 ? GEN_85 : reg_sbadaddr;
  assign GEN_104 = T_6425 ? GEN_86 : reg_mstatus_spie;
  assign GEN_105 = T_6425 ? GEN_87 : {{1'd0}, reg_mstatus_spp};
  assign GEN_106 = T_6425 ? GEN_88 : reg_mstatus_sie;
  assign GEN_107 = T_6425 ? GEN_96 : reg_mstatus_prv;
  assign GEN_108 = T_6425 ? GEN_90 : reg_mepc;
  assign GEN_109 = T_6425 ? GEN_91 : reg_mcause;
  assign GEN_110 = T_6425 ? GEN_92 : reg_mbadaddr;
  assign GEN_111 = T_6425 ? GEN_93 : reg_mstatus_mpie;
  assign GEN_112 = T_6425 ? GEN_94 : reg_mstatus_mpp;
  assign GEN_113 = T_6425 ? GEN_95 : reg_mstatus_mie;
  assign GEN_114 = reg_mstatus_spp ? reg_mstatus_spie : GEN_106;
  assign GEN_115 = T_6422 ? GEN_114 : GEN_106;
  assign GEN_116 = T_6422 ? 1'h0 : GEN_104;
  assign GEN_117 = T_6422 ? {{1'd0}, 1'h0} : GEN_105;
  assign GEN_118 = T_6422 ? {{1'd0}, reg_mstatus_spp} : GEN_107;
  assign T_6466 = T_6422 == 1'h0;
  assign T_6467 = T_6466 & T_6325;
  assign GEN_119 = T_6467 ? reg_dcsr_prv : GEN_118;
  assign GEN_120 = T_6467 ? 1'h0 : GEN_97;
  assign T_6472 = T_6325 == 1'h0;
  assign T_6473 = T_6466 & T_6472;
  assign T_6474 = reg_mstatus_mpp[1];
  assign GEN_121 = T_6474 ? reg_mstatus_mpie : GEN_113;
  assign T_6476 = reg_mstatus_mpp[0];
  assign T_6479 = T_6474 == 1'h0;
  assign T_6480 = T_6479 & T_6476;
  assign GEN_122 = T_6480 ? reg_mstatus_mpie : GEN_115;
  assign GEN_123 = T_6473 ? GEN_121 : GEN_113;
  assign GEN_124 = T_6473 ? GEN_122 : GEN_115;
  assign GEN_125 = T_6473 ? 1'h0 : GEN_111;
  assign GEN_126 = T_6473 ? {{1'd0}, 1'h0} : GEN_112;
  assign GEN_127 = T_6473 ? reg_mstatus_mpp : GEN_119;
  assign GEN_128 = insn_ret ? GEN_124 : GEN_106;
  assign GEN_129 = insn_ret ? GEN_116 : GEN_104;
  assign GEN_130 = insn_ret ? GEN_117 : GEN_105;
  assign GEN_131 = insn_ret ? GEN_127 : GEN_107;
  assign GEN_132 = insn_ret ? GEN_120 : GEN_97;
  assign GEN_133 = insn_ret ? GEN_123 : GEN_113;
  assign GEN_134 = insn_ret ? GEN_125 : GEN_111;
  assign GEN_135 = insn_ret ? GEN_126 : GEN_112;
  assign T_6485 = {1'h0,csr_xcpt};
  assign GEN_692 = {{1'd0}, io_exception};
  assign T_6486 = GEN_692 + T_6485;
  assign T_6487 = T_6486[1:0];
  assign T_6488 = {1'h0,T_6487};
  assign GEN_693 = {{2'd0}, insn_ret};
  assign T_6489 = GEN_693 + T_6488;
  assign T_6490 = T_6489[2:0];
  assign GEN_694 = {{2'd0}, 1'h1};
  assign T_6492 = T_6490 <= GEN_694;
  assign T_6493 = T_6492 | reset;
  assign T_6495 = T_6493 == 1'h0;
  assign T_6497 = T_6194 ? T_6041 : {{63'd0}, 1'h0};
  assign T_6499 = T_6196 ? T_6066 : {{63'd0}, 1'h0};
  assign GEN_12 = GEN_136;
  assign GEN_136 = reg_tdrselect_tdrindex ? reg_bp_1_address : reg_bp_0_address;
  assign T_6501 = T_6198 ? GEN_12 : {{38'd0}, 1'h0};
  assign T_6509 = T_6206 ? reg_cycle : {{63'd0}, 1'h0};
  assign T_6511 = T_6208 ? T_5748 : {{63'd0}, 1'h0};
  assign T_6521 = T_6218 ? 64'h8000000000041129 : {{63'd0}, 1'h0};
  assign T_6523 = T_6220 ? read_mstatus : {{63'd0}, 1'h0};
  assign T_6525 = T_6222 ? reg_mtvec : {{31'd0}, 1'h0};
  assign T_6527 = T_6224 ? read_mip : {{12'd0}, 1'h0};
  assign T_6529 = T_6226 ? reg_mie : {{63'd0}, 1'h0};
  assign T_6531 = T_6228 ? reg_mideleg : {{63'd0}, 1'h0};
  assign T_6533 = T_6230 ? reg_medeleg : {{63'd0}, 1'h0};
  assign T_6535 = T_6232 ? reg_mscratch : {{63'd0}, 1'h0};
  assign T_6537 = T_6234 ? T_6093 : {{63'd0}, 1'h0};
  assign T_6539 = T_6236 ? T_6098 : {{63'd0}, 1'h0};
  assign T_6541 = T_6238 ? reg_mcause : {{63'd0}, 1'h0};
  assign T_6543 = T_6240 ? io_prci_id : 1'h0;
  assign T_6545 = T_6242 ? T_6114 : {{31'd0}, 1'h0};
  assign T_6547 = T_6244 ? reg_dpc : {{39'd0}, 1'h0};
  assign T_6549 = T_6246 ? reg_dscratch : {{63'd0}, 1'h0};
  assign T_6551 = T_6248 ? reg_fflags : {{4'd0}, 1'h0};
  assign T_6553 = T_6250 ? reg_frm : {{2'd0}, 1'h0};
  assign T_6555 = T_6252 ? T_6115 : {{7'd0}, 1'h0};
  assign T_6557 = T_6254 ? T_6172 : {{63'd0}, 1'h0};
  assign T_6559 = T_6256 ? T_6117 : {{63'd0}, 1'h0};
  assign T_6561 = T_6258 ? T_6116 : {{63'd0}, 1'h0};
  assign T_6563 = T_6260 ? reg_sscratch : {{63'd0}, 1'h0};
  assign T_6565 = T_6262 ? reg_scause : {{63'd0}, 1'h0};
  assign T_6567 = T_6264 ? T_6177 : {{63'd0}, 1'h0};
  assign T_6569 = T_6266 ? reg_sptbr : {{19'd0}, 1'h0};
  assign T_6573 = T_6270 ? T_6183 : {{63'd0}, 1'h0};
  assign T_6575 = T_6272 ? T_6188 : {{63'd0}, 1'h0};
  assign T_6585 = T_6497 | T_6499;
  assign GEN_695 = {{25'd0}, T_6501};
  assign T_6586 = T_6585 | GEN_695;
  assign T_6587 = T_6586 | GEN_637;
  assign T_6588 = T_6587 | GEN_637;
  assign T_6589 = T_6588 | GEN_637;
  assign T_6590 = T_6589 | T_6509;
  assign T_6591 = T_6590 | T_6511;
  assign T_6592 = T_6591 | GEN_637;
  assign T_6593 = T_6592 | GEN_637;
  assign T_6594 = T_6593 | GEN_637;
  assign T_6595 = T_6594 | GEN_637;
  assign T_6596 = T_6595 | T_6521;
  assign T_6597 = T_6596 | T_6523;
  assign GEN_703 = {{32'd0}, T_6525};
  assign T_6598 = T_6597 | GEN_703;
  assign GEN_704 = {{51'd0}, T_6527};
  assign T_6599 = T_6598 | GEN_704;
  assign T_6600 = T_6599 | T_6529;
  assign T_6601 = T_6600 | T_6531;
  assign T_6602 = T_6601 | T_6533;
  assign T_6603 = T_6602 | T_6535;
  assign T_6604 = T_6603 | T_6537;
  assign T_6605 = T_6604 | T_6539;
  assign T_6606 = T_6605 | T_6541;
  assign GEN_705 = {{63'd0}, T_6543};
  assign T_6607 = T_6606 | GEN_705;
  assign GEN_706 = {{32'd0}, T_6545};
  assign T_6608 = T_6607 | GEN_706;
  assign GEN_707 = {{24'd0}, T_6547};
  assign T_6609 = T_6608 | GEN_707;
  assign T_6610 = T_6609 | T_6549;
  assign GEN_708 = {{59'd0}, T_6551};
  assign T_6611 = T_6610 | GEN_708;
  assign GEN_709 = {{61'd0}, T_6553};
  assign T_6612 = T_6611 | GEN_709;
  assign GEN_710 = {{56'd0}, T_6555};
  assign T_6613 = T_6612 | GEN_710;
  assign T_6614 = T_6613 | T_6557;
  assign T_6615 = T_6614 | T_6559;
  assign T_6616 = T_6615 | T_6561;
  assign T_6617 = T_6616 | T_6563;
  assign T_6618 = T_6617 | T_6565;
  assign T_6619 = T_6618 | T_6567;
  assign GEN_711 = {{44'd0}, T_6569};
  assign T_6620 = T_6619 | GEN_711;
  assign T_6621 = T_6620 | GEN_637;
  assign T_6622 = T_6621 | T_6573;
  assign T_6623 = T_6622 | T_6575;
  assign T_6624 = T_6623 | GEN_637;
  assign T_6625 = T_6624 | GEN_637;
  assign T_6626 = T_6625 | GEN_637;
  assign T_6627 = T_6626 | GEN_637;
  assign T_6628 = T_6627;
  assign T_6629 = reg_fflags | io_fcsr_flags_bits;
  assign GEN_137 = io_fcsr_flags_valid ? T_6629 : reg_fflags;
  assign supportedModes_0 = 2'h3;
  assign supportedModes_1 = {{1'd0}, 1'h0};
  assign supportedModes_2 = {{1'd0}, 1'h1};
  assign T_6687_debug = T_6735;
  assign T_6687_prv = T_6734;
  assign T_6687_sd = T_6733;
  assign T_6687_zero3 = T_6732;
  assign T_6687_sd_rv32 = T_6731;
  assign T_6687_zero2 = T_6730;
  assign T_6687_vm = T_6729;
  assign T_6687_zero1 = T_6728;
  assign T_6687_pum = T_6727;
  assign T_6687_mprv = T_6726;
  assign T_6687_xs = T_6725;
  assign T_6687_fs = T_6724;
  assign T_6687_mpp = T_6723;
  assign T_6687_hpp = T_6722;
  assign T_6687_spp = T_6721;
  assign T_6687_mpie = T_6720;
  assign T_6687_hpie = T_6719;
  assign T_6687_spie = T_6718;
  assign T_6687_upie = T_6717;
  assign T_6687_mie = T_6716;
  assign T_6687_hie = T_6715;
  assign T_6687_sie = T_6714;
  assign T_6687_uie = T_6713;
  assign T_6712 = {{3'd0}, wdata};
  assign T_6713 = T_6712[0];
  assign T_6714 = T_6712[1];
  assign T_6715 = T_6712[2];
  assign T_6716 = T_6712[3];
  assign T_6717 = T_6712[4];
  assign T_6718 = T_6712[5];
  assign T_6719 = T_6712[6];
  assign T_6720 = T_6712[7];
  assign T_6721 = T_6712[8];
  assign T_6722 = T_6712[10:9];
  assign T_6723 = T_6712[12:11];
  assign T_6724 = T_6712[14:13];
  assign T_6725 = T_6712[16:15];
  assign T_6726 = T_6712[17];
  assign T_6727 = T_6712[18];
  assign T_6728 = T_6712[23:19];
  assign T_6729 = T_6712[28:24];
  assign T_6730 = T_6712[30:29];
  assign T_6731 = T_6712[31];
  assign T_6732 = T_6712[62:32];
  assign T_6733 = T_6712[63];
  assign T_6734 = T_6712[65:64];
  assign T_6735 = T_6712[66];
  assign T_6736 = supportedModes_0 == T_6687_mpp;
  assign T_6737 = supportedModes_1 == T_6687_mpp;
  assign T_6738 = supportedModes_2 == T_6687_mpp;
  assign T_6741 = T_6736 | T_6737;
  assign T_6742 = T_6741 | T_6738;
  assign GEN_138 = T_6742 ? T_6687_mpp : GEN_135;
  assign GEN_717 = {{4'd0}, 1'h0};
  assign T_6744 = T_6687_vm == GEN_717;
  assign GEN_139 = T_6744 ? {{4'd0}, 1'h0} : reg_mstatus_vm;
  assign GEN_718 = {{1'd0}, 4'h9};
  assign T_6747 = T_6687_vm == GEN_718;
  assign GEN_140 = T_6747 ? {{1'd0}, 4'h9} : GEN_139;
  assign T_6750 = T_6687_fs != GEN_681;
  assign GEN_720 = {{1'd0}, T_6750};
  assign T_6752 = 2'h0 - GEN_720;
  assign T_6753 = T_6752[1:0];
  assign GEN_165 = T_6220 ? T_6687_mie : GEN_133;
  assign GEN_166 = T_6220 ? T_6687_mpie : GEN_134;
  assign GEN_167 = T_6220 ? T_6687_mprv : reg_mstatus_mprv;
  assign GEN_168 = T_6220 ? GEN_138 : GEN_135;
  assign GEN_169 = T_6220 ? T_6687_pum : reg_mstatus_pum;
  assign GEN_170 = T_6220 ? {{1'd0}, T_6687_spp} : GEN_130;
  assign GEN_171 = T_6220 ? T_6687_spie : GEN_129;
  assign GEN_172 = T_6220 ? T_6687_sie : GEN_128;
  assign GEN_173 = T_6220 ? GEN_140 : reg_mstatus_vm;
  assign GEN_174 = T_6220 ? T_6753 : reg_mstatus_fs;
  assign T_6782_rocc = T_6808;
  assign T_6782_meip = T_6807;
  assign T_6782_heip = T_6806;
  assign T_6782_seip = T_6805;
  assign T_6782_ueip = T_6804;
  assign T_6782_mtip = T_6803;
  assign T_6782_htip = T_6802;
  assign T_6782_stip = T_6801;
  assign T_6782_utip = T_6800;
  assign T_6782_msip = T_6799;
  assign T_6782_hsip = T_6798;
  assign T_6782_ssip = T_6797;
  assign T_6782_usip = T_6796;
  assign T_6796 = wdata[0];
  assign T_6797 = wdata[1];
  assign T_6798 = wdata[2];
  assign T_6799 = wdata[3];
  assign T_6800 = wdata[4];
  assign T_6801 = wdata[5];
  assign T_6802 = wdata[6];
  assign T_6803 = wdata[7];
  assign T_6804 = wdata[8];
  assign T_6805 = wdata[9];
  assign T_6806 = wdata[10];
  assign T_6807 = wdata[11];
  assign T_6808 = wdata[12];
  assign GEN_188 = T_6224 ? T_6782_ssip : reg_mip_ssip;
  assign GEN_189 = T_6224 ? T_6782_stip : reg_mip_stip;
  assign GEN_721 = {{51'd0}, supported_interrupts};
  assign T_6809 = wdata & GEN_721;
  assign GEN_190 = T_6226 ? T_6809 : reg_mie;
  assign T_6810 = ~ wdata;
  assign T_6812 = T_6810 | GEN_688;
  assign T_6813 = ~ T_6812;
  assign GEN_191 = T_6234 ? T_6813 : {{24'd0}, GEN_108};
  assign GEN_192 = T_6232 ? wdata : reg_mscratch;
  assign T_6814 = wdata[63:2];
  assign GEN_723 = {{2'd0}, T_6814};
  assign T_6815 = GEN_723 << 2;
  assign GEN_193 = T_6222 ? T_6815 : {{32'd0}, reg_mtvec};
  assign T_6817 = wdata & 64'h800000000000001f;
  assign GEN_194 = T_6238 ? T_6817 : GEN_109;
  assign T_6818 = wdata[39:0];
  assign GEN_195 = T_6236 ? T_6818 : GEN_110;
  assign GEN_196 = T_6248 ? wdata : {{59'd0}, GEN_137};
  assign GEN_197 = T_6250 ? wdata : {{61'd0}, reg_frm};
  assign T_6819 = wdata[63:5];
  assign GEN_198 = T_6252 ? wdata : GEN_196;
  assign GEN_199 = T_6252 ? {{5'd0}, T_6819} : GEN_197;
  assign T_6856_xdebugver = T_6890;
  assign T_6856_ndreset = T_6889;
  assign T_6856_fullreset = T_6888;
  assign T_6856_hwbpcount = T_6887;
  assign T_6856_ebreakm = T_6886;
  assign T_6856_ebreakh = T_6885;
  assign T_6856_ebreaks = T_6884;
  assign T_6856_ebreaku = T_6808;
  assign T_6856_zero2 = T_6807;
  assign T_6856_stopcycle = T_6806;
  assign T_6856_stoptime = T_6805;
  assign T_6856_cause = T_6879;
  assign T_6856_debugint = T_6801;
  assign T_6856_zero1 = T_6800;
  assign T_6856_halt = T_6799;
  assign T_6856_step = T_6798;
  assign T_6856_prv = T_6874;
  assign T_6874 = wdata[1:0];
  assign T_6879 = wdata[8:6];
  assign T_6884 = wdata[13];
  assign T_6885 = wdata[14];
  assign T_6886 = wdata[15];
  assign T_6887 = wdata[27:16];
  assign T_6888 = wdata[28];
  assign T_6889 = wdata[29];
  assign T_6890 = wdata[31:30];
  assign GEN_217 = T_6242 ? T_6856_halt : reg_dcsr_halt;
  assign GEN_218 = T_6242 ? T_6856_ebreakm : reg_dcsr_ebreakm;
  assign GEN_219 = T_6242 ? T_6856_ebreaks : reg_dcsr_ebreaks;
  assign GEN_220 = T_6242 ? T_6856_ebreaku : reg_dcsr_ebreaku;
  assign GEN_221 = T_6242 ? T_6856_prv : GEN_100;
  assign GEN_222 = T_6244 ? T_6813 : {{24'd0}, GEN_98};
  assign GEN_223 = T_6246 ? wdata : reg_dscratch;
  assign T_6943_debug = T_6991;
  assign T_6943_prv = T_6990;
  assign T_6943_sd = T_6989;
  assign T_6943_zero3 = T_6988;
  assign T_6943_sd_rv32 = T_6987;
  assign T_6943_zero2 = T_6986;
  assign T_6943_vm = T_6985;
  assign T_6943_zero1 = T_6984;
  assign T_6943_pum = T_6983;
  assign T_6943_mprv = T_6982;
  assign T_6943_xs = T_6981;
  assign T_6943_fs = T_6980;
  assign T_6943_mpp = T_6979;
  assign T_6943_hpp = T_6978;
  assign T_6943_spp = T_6977;
  assign T_6943_mpie = T_6976;
  assign T_6943_hpie = T_6975;
  assign T_6943_spie = T_6974;
  assign T_6943_upie = T_6973;
  assign T_6943_mie = T_6972;
  assign T_6943_hie = T_6971;
  assign T_6943_sie = T_6970;
  assign T_6943_uie = T_6969;
  assign T_6968 = {{3'd0}, wdata};
  assign T_6969 = T_6968[0];
  assign T_6970 = T_6968[1];
  assign T_6971 = T_6968[2];
  assign T_6972 = T_6968[3];
  assign T_6973 = T_6968[4];
  assign T_6974 = T_6968[5];
  assign T_6975 = T_6968[6];
  assign T_6976 = T_6968[7];
  assign T_6977 = T_6968[8];
  assign T_6978 = T_6968[10:9];
  assign T_6979 = T_6968[12:11];
  assign T_6980 = T_6968[14:13];
  assign T_6981 = T_6968[16:15];
  assign T_6982 = T_6968[17];
  assign T_6983 = T_6968[18];
  assign T_6984 = T_6968[23:19];
  assign T_6985 = T_6968[28:24];
  assign T_6986 = T_6968[30:29];
  assign T_6987 = T_6968[31];
  assign T_6988 = T_6968[62:32];
  assign T_6989 = T_6968[63];
  assign T_6990 = T_6968[65:64];
  assign T_6991 = T_6968[66];
  assign T_6993 = T_6943_fs != GEN_681;
  assign GEN_726 = {{1'd0}, T_6993};
  assign T_6995 = 2'h0 - GEN_726;
  assign T_6996 = T_6995[1:0];
  assign GEN_248 = T_6254 ? T_6943_sie : GEN_172;
  assign GEN_249 = T_6254 ? T_6943_spie : GEN_171;
  assign GEN_250 = T_6254 ? {{1'd0}, T_6943_spp} : GEN_170;
  assign GEN_251 = T_6254 ? T_6943_pum : GEN_169;
  assign GEN_252 = T_6254 ? T_6996 : GEN_174;
  assign T_7025_rocc = T_6808;
  assign T_7025_meip = T_6807;
  assign T_7025_heip = T_6806;
  assign T_7025_seip = T_6805;
  assign T_7025_ueip = T_6804;
  assign T_7025_mtip = T_6803;
  assign T_7025_htip = T_6802;
  assign T_7025_stip = T_6801;
  assign T_7025_utip = T_6800;
  assign T_7025_msip = T_6799;
  assign T_7025_hsip = T_6798;
  assign T_7025_ssip = T_6797;
  assign T_7025_usip = T_6796;
  assign GEN_266 = T_6256 ? T_7025_ssip : GEN_188;
  assign T_7053 = reg_mie & T_5799;
  assign T_7054 = wdata & reg_mideleg;
  assign T_7055 = T_7053 | T_7054;
  assign GEN_267 = T_6258 ? T_7055 : GEN_190;
  assign GEN_268 = T_6260 ? wdata : reg_sscratch;
  assign GEN_269 = T_6266 ? wdata : {{44'd0}, reg_sptbr};
  assign GEN_270 = T_6270 ? T_6815 : {{24'd0}, GEN_101};
  assign GEN_271 = T_6272 ? T_6815 : {{25'd0}, reg_stvec};
  assign GEN_272 = T_6262 ? T_6817 : GEN_102;
  assign GEN_273 = T_6264 ? T_6818 : GEN_103;
  assign GEN_729 = {{51'd0}, delegable_interrupts};
  assign T_7063 = wdata & GEN_729;
  assign GEN_274 = T_6228 ? T_7063 : reg_mideleg;
  assign GEN_730 = {{55'd0}, 9'h1ab};
  assign T_7064 = wdata & GEN_730;
  assign GEN_275 = T_6230 ? T_7064 : reg_medeleg;
  assign T_7073_tdrmode = T_7079;
  assign T_7073_reserved = T_7078;
  assign T_7073_tdrindex = T_6796;
  assign T_7078 = wdata[62:1];
  assign T_7079 = wdata[63];
  assign GEN_276 = T_6194 ? T_7073_tdrindex : reg_tdrselect_tdrindex;
  assign T_7080 = reg_tdrselect_tdrmode | reg_debug;
  assign T_7107_tdrtype = T_7131;
  assign T_7107_bpamaskmax = T_7130;
  assign T_7107_reserved = T_7129;
  assign T_7107_bpaction = T_7128;
  assign T_7107_bpmatch = T_7127;
  assign T_7107_m = T_6802;
  assign T_7107_h = T_6801;
  assign T_7107_s = T_6800;
  assign T_7107_u = T_6799;
  assign T_7107_r = T_6798;
  assign T_7107_w = T_6797;
  assign T_7107_x = T_6796;
  assign T_7127 = wdata[10:7];
  assign T_7128 = wdata[18:11];
  assign T_7129 = wdata[54:19];
  assign T_7130 = wdata[59:55];
  assign T_7131 = wdata[63:60];
  assign GEN_13 = T_7107_tdrtype;
  assign GEN_14 = T_7107_bpamaskmax;
  assign GEN_15 = T_7107_reserved;
  assign GEN_16 = T_7107_bpaction;
  assign GEN_17 = T_7107_bpmatch;
  assign GEN_285 = 1'h0 == reg_tdrselect_tdrindex ? GEN_17 : reg_bp_0_control_bpmatch;
  assign GEN_18 = T_7107_m;
  assign GEN_287 = 1'h0 == reg_tdrselect_tdrindex ? GEN_18 : reg_bp_0_control_m;
  assign GEN_19 = T_7107_h;
  assign GEN_20 = T_7107_s;
  assign GEN_291 = 1'h0 == reg_tdrselect_tdrindex ? GEN_20 : reg_bp_0_control_s;
  assign GEN_21 = T_7107_u;
  assign GEN_293 = 1'h0 == reg_tdrselect_tdrindex ? GEN_21 : reg_bp_0_control_u;
  assign GEN_22 = T_7107_r;
  assign GEN_295 = 1'h0 == reg_tdrselect_tdrindex ? GEN_22 : reg_bp_0_control_r;
  assign GEN_23 = T_7107_w;
  assign GEN_297 = 1'h0 == reg_tdrselect_tdrindex ? GEN_23 : reg_bp_0_control_w;
  assign GEN_24 = T_7107_x;
  assign GEN_299 = 1'h0 == reg_tdrselect_tdrindex ? GEN_24 : reg_bp_0_control_x;
  assign GEN_731 = {{2'd0}, 2'h2};
  assign T_7161 = T_7107_bpmatch & GEN_731;
  assign GEN_25 = T_7161;
  assign GEN_301 = 1'h0 == reg_tdrselect_tdrindex ? GEN_25 : GEN_285;
  assign GEN_328 = T_6196 ? GEN_301 : reg_bp_0_control_bpmatch;
  assign GEN_331 = T_6196 ? GEN_287 : reg_bp_0_control_m;
  assign GEN_337 = T_6196 ? GEN_291 : reg_bp_0_control_s;
  assign GEN_340 = T_6196 ? GEN_293 : reg_bp_0_control_u;
  assign GEN_343 = T_6196 ? GEN_295 : reg_bp_0_control_r;
  assign GEN_346 = T_6196 ? GEN_297 : reg_bp_0_control_w;
  assign GEN_349 = T_6196 ? GEN_299 : reg_bp_0_control_x;
  assign GEN_26 = wdata[38:0];
  assign GEN_352 = 1'h0 == reg_tdrselect_tdrindex ? GEN_26 : reg_bp_0_address;
  assign GEN_355 = T_6198 ? GEN_352 : reg_bp_0_address;
  assign GEN_382 = T_7080 ? GEN_328 : reg_bp_0_control_bpmatch;
  assign GEN_385 = T_7080 ? GEN_331 : reg_bp_0_control_m;
  assign GEN_391 = T_7080 ? GEN_337 : reg_bp_0_control_s;
  assign GEN_394 = T_7080 ? GEN_340 : reg_bp_0_control_u;
  assign GEN_397 = T_7080 ? GEN_343 : reg_bp_0_control_r;
  assign GEN_400 = T_7080 ? GEN_346 : reg_bp_0_control_w;
  assign GEN_403 = T_7080 ? GEN_349 : reg_bp_0_control_x;
  assign GEN_407 = T_7080 ? GEN_355 : reg_bp_0_address;
  assign GEN_433 = wen ? GEN_165 : GEN_133;
  assign GEN_434 = wen ? GEN_166 : GEN_134;
  assign GEN_435 = wen ? GEN_167 : reg_mstatus_mprv;
  assign GEN_436 = wen ? GEN_168 : GEN_135;
  assign GEN_437 = wen ? GEN_251 : reg_mstatus_pum;
  assign GEN_438 = wen ? GEN_250 : GEN_130;
  assign GEN_439 = wen ? GEN_249 : GEN_129;
  assign GEN_440 = wen ? GEN_248 : GEN_128;
  assign GEN_441 = wen ? GEN_173 : reg_mstatus_vm;
  assign GEN_442 = wen ? GEN_252 : reg_mstatus_fs;
  assign GEN_456 = wen ? GEN_266 : reg_mip_ssip;
  assign GEN_457 = wen ? GEN_189 : reg_mip_stip;
  assign GEN_458 = wen ? GEN_267 : reg_mie;
  assign GEN_459 = wen ? GEN_191 : {{24'd0}, GEN_108};
  assign GEN_460 = wen ? GEN_192 : reg_mscratch;
  assign GEN_461 = wen ? GEN_193 : {{32'd0}, reg_mtvec};
  assign GEN_462 = wen ? GEN_194 : GEN_109;
  assign GEN_463 = wen ? GEN_195 : GEN_110;
  assign GEN_464 = wen ? GEN_198 : {{59'd0}, GEN_137};
  assign GEN_465 = wen ? GEN_199 : {{61'd0}, reg_frm};
  assign GEN_483 = wen ? GEN_217 : reg_dcsr_halt;
  assign GEN_484 = wen ? GEN_218 : reg_dcsr_ebreakm;
  assign GEN_485 = wen ? GEN_219 : reg_dcsr_ebreaks;
  assign GEN_486 = wen ? GEN_220 : reg_dcsr_ebreaku;
  assign GEN_487 = wen ? GEN_221 : GEN_100;
  assign GEN_488 = wen ? GEN_222 : {{24'd0}, GEN_98};
  assign GEN_489 = wen ? GEN_223 : reg_dscratch;
  assign GEN_527 = wen ? GEN_268 : reg_sscratch;
  assign GEN_528 = wen ? GEN_269 : {{44'd0}, reg_sptbr};
  assign GEN_529 = wen ? GEN_270 : {{24'd0}, GEN_101};
  assign GEN_530 = wen ? GEN_271 : {{25'd0}, reg_stvec};
  assign GEN_531 = wen ? GEN_272 : GEN_102;
  assign GEN_532 = wen ? GEN_273 : GEN_103;
  assign GEN_533 = wen ? GEN_274 : reg_mideleg;
  assign GEN_534 = wen ? GEN_275 : reg_medeleg;
  assign GEN_538 = wen ? GEN_276 : reg_tdrselect_tdrindex;
  assign GEN_564 = wen ? GEN_382 : reg_bp_0_control_bpmatch;
  assign GEN_567 = wen ? GEN_385 : reg_bp_0_control_m;
  assign GEN_573 = wen ? GEN_391 : reg_bp_0_control_s;
  assign GEN_576 = wen ? GEN_394 : reg_bp_0_control_u;
  assign GEN_579 = wen ? GEN_397 : reg_bp_0_control_r;
  assign GEN_582 = wen ? GEN_400 : reg_bp_0_control_w;
  assign GEN_585 = wen ? GEN_403 : reg_bp_0_control_x;
  assign GEN_589 = wen ? GEN_407 : reg_bp_0_address;
  assign GEN_591 = reset ? 1'h0 : GEN_579;
  assign GEN_592 = reset ? 1'h0 : GEN_582;
  assign GEN_593 = reset ? 1'h0 : GEN_585;
  assign T_7226_control_tdrtype = T_7255;
  assign T_7226_control_bpamaskmax = T_7254;
  assign T_7226_control_reserved = T_7253;
  assign T_7226_control_bpaction = T_7252;
  assign T_7226_control_bpmatch = T_7251;
  assign T_7226_control_m = T_7250;
  assign T_7226_control_h = T_7249;
  assign T_7226_control_s = T_7248;
  assign T_7226_control_u = T_7247;
  assign T_7226_control_r = T_7246;
  assign T_7226_control_w = T_7245;
  assign T_7226_control_x = T_7244;
  assign T_7226_address = T_7243;
  assign T_7242 = {{102'd0}, 1'h0};
  assign T_7243 = T_7242[38:0];
  assign T_7244 = T_7242[39];
  assign T_7245 = T_7242[40];
  assign T_7246 = T_7242[41];
  assign T_7247 = T_7242[42];
  assign T_7248 = T_7242[43];
  assign T_7249 = T_7242[44];
  assign T_7250 = T_7242[45];
  assign T_7251 = T_7242[49:46];
  assign T_7252 = T_7242[57:50];
  assign T_7253 = T_7242[93:58];
  assign T_7254 = T_7242[98:94];
  assign T_7255 = T_7242[102:99];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_237 = {1{$random}};
  reg_mstatus_debug = GEN_237[0:0];
  GEN_238 = {1{$random}};
  reg_mstatus_prv = GEN_238[1:0];
  GEN_239 = {1{$random}};
  reg_mstatus_sd = GEN_239[0:0];
  GEN_240 = {1{$random}};
  reg_mstatus_zero3 = GEN_240[30:0];
  GEN_241 = {1{$random}};
  reg_mstatus_sd_rv32 = GEN_241[0:0];
  GEN_242 = {1{$random}};
  reg_mstatus_zero2 = GEN_242[1:0];
  GEN_243 = {1{$random}};
  reg_mstatus_vm = GEN_243[4:0];
  GEN_244 = {1{$random}};
  reg_mstatus_zero1 = GEN_244[4:0];
  GEN_245 = {1{$random}};
  reg_mstatus_pum = GEN_245[0:0];
  GEN_246 = {1{$random}};
  reg_mstatus_mprv = GEN_246[0:0];
  GEN_247 = {1{$random}};
  reg_mstatus_xs = GEN_247[1:0];
  GEN_253 = {1{$random}};
  reg_mstatus_fs = GEN_253[1:0];
  GEN_254 = {1{$random}};
  reg_mstatus_mpp = GEN_254[1:0];
  GEN_255 = {1{$random}};
  reg_mstatus_hpp = GEN_255[1:0];
  GEN_256 = {1{$random}};
  reg_mstatus_spp = GEN_256[0:0];
  GEN_257 = {1{$random}};
  reg_mstatus_mpie = GEN_257[0:0];
  GEN_258 = {1{$random}};
  reg_mstatus_hpie = GEN_258[0:0];
  GEN_259 = {1{$random}};
  reg_mstatus_spie = GEN_259[0:0];
  GEN_260 = {1{$random}};
  reg_mstatus_upie = GEN_260[0:0];
  GEN_261 = {1{$random}};
  reg_mstatus_mie = GEN_261[0:0];
  GEN_262 = {1{$random}};
  reg_mstatus_hie = GEN_262[0:0];
  GEN_263 = {1{$random}};
  reg_mstatus_sie = GEN_263[0:0];
  GEN_264 = {1{$random}};
  reg_mstatus_uie = GEN_264[0:0];
  GEN_265 = {1{$random}};
  reg_dcsr_xdebugver = GEN_265[1:0];
  GEN_277 = {1{$random}};
  reg_dcsr_ndreset = GEN_277[0:0];
  GEN_278 = {1{$random}};
  reg_dcsr_fullreset = GEN_278[0:0];
  GEN_279 = {1{$random}};
  reg_dcsr_hwbpcount = GEN_279[11:0];
  GEN_280 = {1{$random}};
  reg_dcsr_ebreakm = GEN_280[0:0];
  GEN_281 = {1{$random}};
  reg_dcsr_ebreakh = GEN_281[0:0];
  GEN_282 = {1{$random}};
  reg_dcsr_ebreaks = GEN_282[0:0];
  GEN_283 = {1{$random}};
  reg_dcsr_ebreaku = GEN_283[0:0];
  GEN_284 = {1{$random}};
  reg_dcsr_zero2 = GEN_284[0:0];
  GEN_286 = {1{$random}};
  reg_dcsr_stopcycle = GEN_286[0:0];
  GEN_288 = {1{$random}};
  reg_dcsr_stoptime = GEN_288[0:0];
  GEN_289 = {1{$random}};
  reg_dcsr_cause = GEN_289[2:0];
  GEN_290 = {1{$random}};
  reg_dcsr_debugint = GEN_290[0:0];
  GEN_292 = {1{$random}};
  reg_dcsr_zero1 = GEN_292[0:0];
  GEN_294 = {1{$random}};
  reg_dcsr_halt = GEN_294[0:0];
  GEN_296 = {1{$random}};
  reg_dcsr_step = GEN_296[0:0];
  GEN_298 = {1{$random}};
  reg_dcsr_prv = GEN_298[1:0];
  GEN_300 = {1{$random}};
  reg_debug = GEN_300[0:0];
  GEN_302 = {2{$random}};
  reg_dpc = GEN_302[39:0];
  GEN_303 = {2{$random}};
  reg_dscratch = GEN_303[63:0];
  GEN_304 = {1{$random}};
  reg_tdrselect_tdrmode = GEN_304[0:0];
  GEN_305 = {2{$random}};
  reg_tdrselect_reserved = GEN_305[61:0];
  GEN_306 = {1{$random}};
  reg_tdrselect_tdrindex = GEN_306[0:0];
  GEN_307 = {1{$random}};
  reg_bp_0_control_tdrtype = GEN_307[3:0];
  GEN_308 = {1{$random}};
  reg_bp_0_control_bpamaskmax = GEN_308[4:0];
  GEN_309 = {2{$random}};
  reg_bp_0_control_reserved = GEN_309[35:0];
  GEN_310 = {1{$random}};
  reg_bp_0_control_bpaction = GEN_310[7:0];
  GEN_311 = {1{$random}};
  reg_bp_0_control_bpmatch = GEN_311[3:0];
  GEN_312 = {1{$random}};
  reg_bp_0_control_m = GEN_312[0:0];
  GEN_313 = {1{$random}};
  reg_bp_0_control_h = GEN_313[0:0];
  GEN_314 = {1{$random}};
  reg_bp_0_control_s = GEN_314[0:0];
  GEN_315 = {1{$random}};
  reg_bp_0_control_u = GEN_315[0:0];
  GEN_316 = {1{$random}};
  reg_bp_0_control_r = GEN_316[0:0];
  GEN_317 = {1{$random}};
  reg_bp_0_control_w = GEN_317[0:0];
  GEN_318 = {1{$random}};
  reg_bp_0_control_x = GEN_318[0:0];
  GEN_319 = {2{$random}};
  reg_bp_0_address = GEN_319[38:0];
  GEN_320 = {1{$random}};
  reg_bp_1_control_tdrtype = GEN_320[3:0];
  GEN_321 = {1{$random}};
  reg_bp_1_control_bpamaskmax = GEN_321[4:0];
  GEN_322 = {2{$random}};
  reg_bp_1_control_reserved = GEN_322[35:0];
  GEN_323 = {1{$random}};
  reg_bp_1_control_bpaction = GEN_323[7:0];
  GEN_324 = {1{$random}};
  reg_bp_1_control_bpmatch = GEN_324[3:0];
  GEN_325 = {1{$random}};
  reg_bp_1_control_m = GEN_325[0:0];
  GEN_326 = {1{$random}};
  reg_bp_1_control_h = GEN_326[0:0];
  GEN_327 = {1{$random}};
  reg_bp_1_control_s = GEN_327[0:0];
  GEN_329 = {1{$random}};
  reg_bp_1_control_u = GEN_329[0:0];
  GEN_330 = {1{$random}};
  reg_bp_1_control_r = GEN_330[0:0];
  GEN_332 = {1{$random}};
  reg_bp_1_control_w = GEN_332[0:0];
  GEN_333 = {1{$random}};
  reg_bp_1_control_x = GEN_333[0:0];
  GEN_334 = {2{$random}};
  reg_bp_1_address = GEN_334[38:0];
  GEN_335 = {2{$random}};
  reg_mie = GEN_335[63:0];
  GEN_336 = {2{$random}};
  reg_mideleg = GEN_336[63:0];
  GEN_338 = {2{$random}};
  reg_medeleg = GEN_338[63:0];
  GEN_339 = {1{$random}};
  reg_mip_rocc = GEN_339[0:0];
  GEN_341 = {1{$random}};
  reg_mip_meip = GEN_341[0:0];
  GEN_342 = {1{$random}};
  reg_mip_heip = GEN_342[0:0];
  GEN_344 = {1{$random}};
  reg_mip_seip = GEN_344[0:0];
  GEN_345 = {1{$random}};
  reg_mip_ueip = GEN_345[0:0];
  GEN_347 = {1{$random}};
  reg_mip_mtip = GEN_347[0:0];
  GEN_348 = {1{$random}};
  reg_mip_htip = GEN_348[0:0];
  GEN_350 = {1{$random}};
  reg_mip_stip = GEN_350[0:0];
  GEN_351 = {1{$random}};
  reg_mip_utip = GEN_351[0:0];
  GEN_353 = {1{$random}};
  reg_mip_msip = GEN_353[0:0];
  GEN_354 = {1{$random}};
  reg_mip_hsip = GEN_354[0:0];
  GEN_356 = {1{$random}};
  reg_mip_ssip = GEN_356[0:0];
  GEN_357 = {1{$random}};
  reg_mip_usip = GEN_357[0:0];
  GEN_358 = {2{$random}};
  reg_mepc = GEN_358[39:0];
  GEN_359 = {2{$random}};
  reg_mcause = GEN_359[63:0];
  GEN_360 = {2{$random}};
  reg_mbadaddr = GEN_360[39:0];
  GEN_361 = {2{$random}};
  reg_mscratch = GEN_361[63:0];
  GEN_362 = {1{$random}};
  reg_mtvec = GEN_362[31:0];
  GEN_363 = {2{$random}};
  reg_sepc = GEN_363[39:0];
  GEN_364 = {2{$random}};
  reg_scause = GEN_364[63:0];
  GEN_365 = {2{$random}};
  reg_sbadaddr = GEN_365[39:0];
  GEN_366 = {2{$random}};
  reg_sscratch = GEN_366[63:0];
  GEN_367 = {2{$random}};
  reg_stvec = GEN_367[38:0];
  GEN_368 = {1{$random}};
  reg_sptbr = GEN_368[19:0];
  GEN_369 = {1{$random}};
  reg_wfi = GEN_369[0:0];
  GEN_370 = {1{$random}};
  T_5476 = GEN_370[5:0];
  GEN_371 = {2{$random}};
  T_5484 = GEN_371[57:0];
  GEN_372 = {1{$random}};
  T_5492 = GEN_372[5:0];
  GEN_373 = {2{$random}};
  T_5500 = GEN_373[57:0];
  GEN_374 = {1{$random}};
  T_5508 = GEN_374[5:0];
  GEN_375 = {2{$random}};
  T_5516 = GEN_375[57:0];
  GEN_376 = {1{$random}};
  T_5524 = GEN_376[5:0];
  GEN_377 = {2{$random}};
  T_5532 = GEN_377[57:0];
  GEN_378 = {1{$random}};
  T_5540 = GEN_378[5:0];
  GEN_379 = {2{$random}};
  T_5548 = GEN_379[57:0];
  GEN_380 = {1{$random}};
  T_5556 = GEN_380[5:0];
  GEN_381 = {2{$random}};
  T_5564 = GEN_381[57:0];
  GEN_383 = {1{$random}};
  T_5572 = GEN_383[5:0];
  GEN_384 = {2{$random}};
  T_5580 = GEN_384[57:0];
  GEN_386 = {1{$random}};
  T_5588 = GEN_386[5:0];
  GEN_387 = {2{$random}};
  T_5596 = GEN_387[57:0];
  GEN_388 = {1{$random}};
  T_5604 = GEN_388[5:0];
  GEN_389 = {2{$random}};
  T_5612 = GEN_389[57:0];
  GEN_390 = {1{$random}};
  T_5620 = GEN_390[5:0];
  GEN_392 = {2{$random}};
  T_5628 = GEN_392[57:0];
  GEN_393 = {1{$random}};
  T_5636 = GEN_393[5:0];
  GEN_395 = {2{$random}};
  T_5644 = GEN_395[57:0];
  GEN_396 = {1{$random}};
  T_5652 = GEN_396[5:0];
  GEN_398 = {2{$random}};
  T_5660 = GEN_398[57:0];
  GEN_399 = {1{$random}};
  T_5668 = GEN_399[5:0];
  GEN_401 = {2{$random}};
  T_5676 = GEN_401[57:0];
  GEN_402 = {1{$random}};
  T_5684 = GEN_402[5:0];
  GEN_404 = {2{$random}};
  T_5692 = GEN_404[57:0];
  GEN_405 = {1{$random}};
  T_5700 = GEN_405[5:0];
  GEN_406 = {2{$random}};
  T_5708 = GEN_406[57:0];
  GEN_408 = {1{$random}};
  T_5716 = GEN_408[5:0];
  GEN_409 = {2{$random}};
  T_5724 = GEN_409[57:0];
  GEN_410 = {1{$random}};
  reg_fflags = GEN_410[4:0];
  GEN_411 = {1{$random}};
  reg_frm = GEN_411[2:0];
  GEN_412 = {1{$random}};
  T_5734 = GEN_412[5:0];
  GEN_413 = {2{$random}};
  T_5742 = GEN_413[57:0];
  GEN_414 = {1{$random}};
  T_5751 = GEN_414[5:0];
  GEN_415 = {2{$random}};
  T_5759 = GEN_415[57:0];
  GEN_416 = {1{$random}};
  GEN_61 = GEN_416[1:0];
  GEN_417 = {1{$random}};
  GEN_141 = GEN_417[0:0];
  GEN_418 = {1{$random}};
  GEN_142 = GEN_418[6:0];
  GEN_419 = {1{$random}};
  GEN_143 = GEN_419[4:0];
  GEN_420 = {1{$random}};
  GEN_144 = GEN_420[4:0];
  GEN_421 = {1{$random}};
  GEN_145 = GEN_421[0:0];
  GEN_422 = {1{$random}};
  GEN_146 = GEN_422[0:0];
  GEN_423 = {1{$random}};
  GEN_147 = GEN_423[0:0];
  GEN_424 = {1{$random}};
  GEN_148 = GEN_424[4:0];
  GEN_425 = {1{$random}};
  GEN_149 = GEN_425[6:0];
  GEN_426 = {2{$random}};
  GEN_150 = GEN_426[63:0];
  GEN_427 = {2{$random}};
  GEN_151 = GEN_427[63:0];
  GEN_428 = {1{$random}};
  GEN_152 = GEN_428[0:0];
  GEN_429 = {1{$random}};
  GEN_153 = GEN_429[0:0];
  GEN_430 = {1{$random}};
  GEN_154 = GEN_430[0:0];
  GEN_431 = {1{$random}};
  GEN_155 = GEN_431[0:0];
  GEN_432 = {2{$random}};
  GEN_156 = GEN_432[39:0];
  GEN_443 = {1{$random}};
  GEN_157 = GEN_443[8:0];
  GEN_444 = {1{$random}};
  GEN_158 = GEN_444[4:0];
  GEN_445 = {1{$random}};
  GEN_159 = GEN_445[2:0];
  GEN_446 = {2{$random}};
  GEN_160 = GEN_446[63:0];
  GEN_447 = {1{$random}};
  GEN_161 = GEN_447[0:0];
  GEN_448 = {1{$random}};
  GEN_162 = GEN_448[0:0];
  GEN_449 = {2{$random}};
  GEN_163 = GEN_449[63:0];
  GEN_450 = {2{$random}};
  GEN_164 = GEN_450[63:0];
  GEN_451 = {1{$random}};
  GEN_175 = GEN_451[0:0];
  GEN_452 = {1{$random}};
  GEN_176 = GEN_452[0:0];
  GEN_453 = {1{$random}};
  GEN_177 = GEN_453[0:0];
  GEN_454 = {1{$random}};
  GEN_178 = GEN_454[0:0];
  GEN_455 = {1{$random}};
  GEN_179 = GEN_455[0:0];
  GEN_466 = {1{$random}};
  GEN_180 = GEN_466[0:0];
  GEN_467 = {1{$random}};
  GEN_181 = GEN_467[0:0];
  GEN_468 = {1{$random}};
  GEN_182 = GEN_468[1:0];
  GEN_469 = {1{$random}};
  GEN_183 = GEN_469[0:0];
  GEN_470 = {1{$random}};
  GEN_184 = GEN_470[30:0];
  GEN_471 = {1{$random}};
  GEN_185 = GEN_471[0:0];
  GEN_472 = {1{$random}};
  GEN_186 = GEN_472[1:0];
  GEN_473 = {1{$random}};
  GEN_187 = GEN_473[4:0];
  GEN_474 = {1{$random}};
  GEN_200 = GEN_474[4:0];
  GEN_475 = {1{$random}};
  GEN_201 = GEN_475[0:0];
  GEN_476 = {1{$random}};
  GEN_202 = GEN_476[0:0];
  GEN_477 = {1{$random}};
  GEN_203 = GEN_477[1:0];
  GEN_478 = {1{$random}};
  GEN_204 = GEN_478[1:0];
  GEN_479 = {1{$random}};
  GEN_205 = GEN_479[1:0];
  GEN_480 = {1{$random}};
  GEN_206 = GEN_480[1:0];
  GEN_481 = {1{$random}};
  GEN_207 = GEN_481[0:0];
  GEN_482 = {1{$random}};
  GEN_208 = GEN_482[0:0];
  GEN_490 = {1{$random}};
  GEN_209 = GEN_490[0:0];
  GEN_491 = {1{$random}};
  GEN_210 = GEN_491[0:0];
  GEN_492 = {1{$random}};
  GEN_211 = GEN_492[0:0];
  GEN_493 = {1{$random}};
  GEN_212 = GEN_493[0:0];
  GEN_494 = {1{$random}};
  GEN_213 = GEN_494[0:0];
  GEN_495 = {1{$random}};
  GEN_214 = GEN_495[0:0];
  GEN_496 = {1{$random}};
  GEN_215 = GEN_496[0:0];
  GEN_497 = {1{$random}};
  GEN_216 = GEN_497[0:0];
  GEN_498 = {1{$random}};
  GEN_224 = GEN_498[0:0];
  GEN_499 = {1{$random}};
  GEN_225 = GEN_499[2:0];
  GEN_500 = {1{$random}};
  GEN_226 = GEN_500[1:0];
  GEN_501 = {1{$random}};
  GEN_227 = GEN_501[2:0];
  GEN_502 = {1{$random}};
  GEN_228 = GEN_502[0:0];
  GEN_503 = {1{$random}};
  GEN_229 = GEN_503[3:0];
  GEN_504 = {2{$random}};
  GEN_230 = GEN_504[63:0];
  GEN_505 = {1{$random}};
  GEN_231 = GEN_505[0:0];
  GEN_506 = {1{$random}};
  GEN_232 = GEN_506[0:0];
  GEN_507 = {3{$random}};
  GEN_233 = GEN_507[64:0];
  GEN_508 = {1{$random}};
  GEN_234 = GEN_508[4:0];
  GEN_509 = {1{$random}};
  GEN_235 = GEN_509[0:0];
  GEN_510 = {1{$random}};
  GEN_236 = GEN_510[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      reg_mstatus_debug <= reset_mstatus_debug;
    end
    if(reset) begin
      reg_mstatus_prv <= reset_mstatus_prv;
    end else begin
      reg_mstatus_prv <= GEN_131;
    end
    if(reset) begin
      reg_mstatus_sd <= reset_mstatus_sd;
    end
    if(reset) begin
      reg_mstatus_zero3 <= reset_mstatus_zero3;
    end
    if(reset) begin
      reg_mstatus_sd_rv32 <= reset_mstatus_sd_rv32;
    end
    if(reset) begin
      reg_mstatus_zero2 <= reset_mstatus_zero2;
    end
    if(reset) begin
      reg_mstatus_vm <= reset_mstatus_vm;
    end else begin
      reg_mstatus_vm <= GEN_441;
    end
    if(reset) begin
      reg_mstatus_zero1 <= reset_mstatus_zero1;
    end
    if(reset) begin
      reg_mstatus_pum <= reset_mstatus_pum;
    end else begin
      reg_mstatus_pum <= GEN_437;
    end
    if(reset) begin
      reg_mstatus_mprv <= reset_mstatus_mprv;
    end else begin
      reg_mstatus_mprv <= GEN_435;
    end
    if(reset) begin
      reg_mstatus_xs <= reset_mstatus_xs;
    end
    if(reset) begin
      reg_mstatus_fs <= reset_mstatus_fs;
    end else begin
      reg_mstatus_fs <= GEN_442;
    end
    if(reset) begin
      reg_mstatus_mpp <= reset_mstatus_mpp;
    end else begin
      reg_mstatus_mpp <= GEN_436;
    end
    if(reset) begin
      reg_mstatus_hpp <= reset_mstatus_hpp;
    end
    if(reset) begin
      reg_mstatus_spp <= reset_mstatus_spp;
    end else begin
      reg_mstatus_spp <= GEN_438[0];
    end
    if(reset) begin
      reg_mstatus_mpie <= reset_mstatus_mpie;
    end else begin
      reg_mstatus_mpie <= GEN_434;
    end
    if(reset) begin
      reg_mstatus_hpie <= reset_mstatus_hpie;
    end
    if(reset) begin
      reg_mstatus_spie <= reset_mstatus_spie;
    end else begin
      reg_mstatus_spie <= GEN_439;
    end
    if(reset) begin
      reg_mstatus_upie <= reset_mstatus_upie;
    end
    if(reset) begin
      reg_mstatus_mie <= reset_mstatus_mie;
    end else begin
      reg_mstatus_mie <= GEN_433;
    end
    if(reset) begin
      reg_mstatus_hie <= reset_mstatus_hie;
    end
    if(reset) begin
      reg_mstatus_sie <= reset_mstatus_sie;
    end else begin
      reg_mstatus_sie <= GEN_440;
    end
    if(reset) begin
      reg_mstatus_uie <= reset_mstatus_uie;
    end
    if(reset) begin
      reg_dcsr_xdebugver <= reset_dcsr_xdebugver;
    end
    if(reset) begin
      reg_dcsr_ndreset <= reset_dcsr_ndreset;
    end
    if(reset) begin
      reg_dcsr_fullreset <= reset_dcsr_fullreset;
    end
    if(reset) begin
      reg_dcsr_hwbpcount <= reset_dcsr_hwbpcount;
    end else begin
      reg_dcsr_hwbpcount <= {{11'd0}, 1'h1};
    end
    if(reset) begin
      reg_dcsr_ebreakm <= reset_dcsr_ebreakm;
    end else begin
      reg_dcsr_ebreakm <= GEN_484;
    end
    if(reset) begin
      reg_dcsr_ebreakh <= reset_dcsr_ebreakh;
    end
    if(reset) begin
      reg_dcsr_ebreaks <= reset_dcsr_ebreaks;
    end else begin
      reg_dcsr_ebreaks <= GEN_485;
    end
    if(reset) begin
      reg_dcsr_ebreaku <= reset_dcsr_ebreaku;
    end else begin
      reg_dcsr_ebreaku <= GEN_486;
    end
    if(reset) begin
      reg_dcsr_zero2 <= reset_dcsr_zero2;
    end
    if(reset) begin
      reg_dcsr_stopcycle <= reset_dcsr_stopcycle;
    end
    if(reset) begin
      reg_dcsr_stoptime <= reset_dcsr_stoptime;
    end
    if(reset) begin
      reg_dcsr_cause <= reset_dcsr_cause;
    end else begin
      reg_dcsr_cause <= GEN_99;
    end
    if(reset) begin
      reg_dcsr_debugint <= reset_dcsr_debugint;
    end else begin
      reg_dcsr_debugint <= io_prci_interrupts_debug;
    end
    if(reset) begin
      reg_dcsr_zero1 <= reset_dcsr_zero1;
    end
    if(reset) begin
      reg_dcsr_halt <= reset_dcsr_halt;
    end else begin
      reg_dcsr_halt <= GEN_483;
    end
    if(reset) begin
      reg_dcsr_step <= reset_dcsr_step;
    end
    if(reset) begin
      reg_dcsr_prv <= reset_dcsr_prv;
    end else begin
      reg_dcsr_prv <= GEN_487;
    end
    if(reset) begin
      reg_debug <= 1'h0;
    end else begin
      reg_debug <= GEN_132;
    end
    if(1'h0) begin
    end else begin
      reg_dpc <= GEN_488[39:0];
    end
    if(1'h0) begin
    end else begin
      reg_dscratch <= GEN_489;
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_tdrmode <= 1'h1;
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_reserved <= {{61'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      reg_tdrselect_tdrindex <= GEN_538;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_tdrtype <= {{3'd0}, 1'h1};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpamaskmax <= {{2'd0}, 3'h4};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_reserved <= {{35'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpaction <= {{7'd0}, 1'h0};
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_bpmatch <= GEN_564;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_m <= GEN_567;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_h <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_s <= GEN_573;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_u <= GEN_576;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_r <= GEN_591;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_w <= GEN_592;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_control_x <= GEN_593;
    end
    if(1'h0) begin
    end else begin
      reg_bp_0_address <= GEN_589;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_tdrtype <= T_7226_control_tdrtype;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpamaskmax <= T_7226_control_bpamaskmax;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_reserved <= T_7226_control_reserved;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpaction <= T_7226_control_bpaction;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_bpmatch <= T_7226_control_bpmatch;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_m <= T_7226_control_m;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_h <= T_7226_control_h;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_s <= T_7226_control_s;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_u <= T_7226_control_u;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_r <= T_7226_control_r;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_w <= T_7226_control_w;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_control_x <= T_7226_control_x;
    end
    if(1'h0) begin
    end else begin
      reg_bp_1_address <= T_7226_address;
    end
    if(reset) begin
      reg_mie <= 64'h0;
    end else begin
      reg_mie <= GEN_458;
    end
    if(reset) begin
      reg_mideleg <= 64'h0;
    end else begin
      reg_mideleg <= GEN_533;
    end
    if(reset) begin
      reg_medeleg <= 64'h0;
    end else begin
      reg_medeleg <= GEN_534;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_meip <= io_prci_interrupts_meip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_seip <= io_prci_interrupts_seip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_mtip <= io_prci_interrupts_mtip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_stip <= GEN_457;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_msip <= io_prci_interrupts_msip;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mip_ssip <= GEN_456;
    end
    if(1'h0) begin
    end
    if(1'h0) begin
    end else begin
      reg_mepc <= GEN_459[39:0];
    end
    if(1'h0) begin
    end else begin
      reg_mcause <= GEN_462;
    end
    if(1'h0) begin
    end else begin
      reg_mbadaddr <= GEN_463;
    end
    if(1'h0) begin
    end else begin
      reg_mscratch <= GEN_460;
    end
    if(reset) begin
      reg_mtvec <= 32'h1010;
    end else begin
      reg_mtvec <= GEN_461[31:0];
    end
    if(1'h0) begin
    end else begin
      reg_sepc <= GEN_529[39:0];
    end
    if(1'h0) begin
    end else begin
      reg_scause <= GEN_531;
    end
    if(1'h0) begin
    end else begin
      reg_sbadaddr <= GEN_532;
    end
    if(1'h0) begin
    end else begin
      reg_sscratch <= GEN_527;
    end
    if(1'h0) begin
    end else begin
      reg_stvec <= GEN_530[38:0];
    end
    if(1'h0) begin
    end else begin
      reg_sptbr <= GEN_528[19:0];
    end
    if(reset) begin
      reg_wfi <= 1'h0;
    end else begin
      reg_wfi <= GEN_78;
    end
    if(reset) begin
      T_5476 <= 6'h0;
    end else begin
      T_5476 <= GEN_27;
    end
    if(reset) begin
      T_5484 <= 58'h0;
    end else begin
      T_5484 <= GEN_28;
    end
    if(reset) begin
      T_5492 <= 6'h0;
    end else begin
      T_5492 <= GEN_29;
    end
    if(reset) begin
      T_5500 <= 58'h0;
    end else begin
      T_5500 <= GEN_30;
    end
    if(reset) begin
      T_5508 <= 6'h0;
    end else begin
      T_5508 <= GEN_31;
    end
    if(reset) begin
      T_5516 <= 58'h0;
    end else begin
      T_5516 <= GEN_32;
    end
    if(reset) begin
      T_5524 <= 6'h0;
    end else begin
      T_5524 <= GEN_33;
    end
    if(reset) begin
      T_5532 <= 58'h0;
    end else begin
      T_5532 <= GEN_34;
    end
    if(reset) begin
      T_5540 <= 6'h0;
    end else begin
      T_5540 <= GEN_35;
    end
    if(reset) begin
      T_5548 <= 58'h0;
    end else begin
      T_5548 <= GEN_36;
    end
    if(reset) begin
      T_5556 <= 6'h0;
    end else begin
      T_5556 <= GEN_37;
    end
    if(reset) begin
      T_5564 <= 58'h0;
    end else begin
      T_5564 <= GEN_38;
    end
    if(reset) begin
      T_5572 <= 6'h0;
    end else begin
      T_5572 <= GEN_39;
    end
    if(reset) begin
      T_5580 <= 58'h0;
    end else begin
      T_5580 <= GEN_40;
    end
    if(reset) begin
      T_5588 <= 6'h0;
    end else begin
      T_5588 <= GEN_41;
    end
    if(reset) begin
      T_5596 <= 58'h0;
    end else begin
      T_5596 <= GEN_42;
    end
    if(reset) begin
      T_5604 <= 6'h0;
    end else begin
      T_5604 <= GEN_43;
    end
    if(reset) begin
      T_5612 <= 58'h0;
    end else begin
      T_5612 <= GEN_44;
    end
    if(reset) begin
      T_5620 <= 6'h0;
    end else begin
      T_5620 <= GEN_45;
    end
    if(reset) begin
      T_5628 <= 58'h0;
    end else begin
      T_5628 <= GEN_46;
    end
    if(reset) begin
      T_5636 <= 6'h0;
    end else begin
      T_5636 <= GEN_47;
    end
    if(reset) begin
      T_5644 <= 58'h0;
    end else begin
      T_5644 <= GEN_48;
    end
    if(reset) begin
      T_5652 <= 6'h0;
    end else begin
      T_5652 <= GEN_49;
    end
    if(reset) begin
      T_5660 <= 58'h0;
    end else begin
      T_5660 <= GEN_50;
    end
    if(reset) begin
      T_5668 <= 6'h0;
    end else begin
      T_5668 <= GEN_51;
    end
    if(reset) begin
      T_5676 <= 58'h0;
    end else begin
      T_5676 <= GEN_52;
    end
    if(reset) begin
      T_5684 <= 6'h0;
    end else begin
      T_5684 <= GEN_53;
    end
    if(reset) begin
      T_5692 <= 58'h0;
    end else begin
      T_5692 <= GEN_54;
    end
    if(reset) begin
      T_5700 <= 6'h0;
    end else begin
      T_5700 <= GEN_55;
    end
    if(reset) begin
      T_5708 <= 58'h0;
    end else begin
      T_5708 <= GEN_56;
    end
    if(reset) begin
      T_5716 <= 6'h0;
    end else begin
      T_5716 <= GEN_57;
    end
    if(reset) begin
      T_5724 <= 58'h0;
    end else begin
      T_5724 <= GEN_58;
    end
    if(1'h0) begin
    end else begin
      reg_fflags <= GEN_464[4:0];
    end
    if(1'h0) begin
    end else begin
      reg_frm <= GEN_465[2:0];
    end
    if(reset) begin
      T_5734 <= 6'h0;
    end else begin
      T_5734 <= GEN_59;
    end
    if(reset) begin
      T_5742 <= 58'h0;
    end else begin
      T_5742 <= GEN_60;
    end
    if(reset) begin
      T_5751 <= 6'h0;
    end else begin
      T_5751 <= T_5757;
    end
    if(reset) begin
      T_5759 <= 58'h0;
    end else begin
      T_5759 <= GEN_62;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6495) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at csr.scala:430 assert(PopCount(insn_ret :: io.exception :: csr_xcpt :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_6495) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module BreakpointUnit(
  input   clk,
  input   reset,
  input   io_status_debug,
  input  [1:0] io_status_prv,
  input   io_status_sd,
  input  [30:0] io_status_zero3,
  input   io_status_sd_rv32,
  input  [1:0] io_status_zero2,
  input  [4:0] io_status_vm,
  input  [4:0] io_status_zero1,
  input   io_status_pum,
  input   io_status_mprv,
  input  [1:0] io_status_xs,
  input  [1:0] io_status_fs,
  input  [1:0] io_status_mpp,
  input  [1:0] io_status_hpp,
  input   io_status_spp,
  input   io_status_mpie,
  input   io_status_hpie,
  input   io_status_spie,
  input   io_status_upie,
  input   io_status_mie,
  input   io_status_hie,
  input   io_status_sie,
  input   io_status_uie,
  input  [3:0] io_bp_0_control_tdrtype,
  input  [4:0] io_bp_0_control_bpamaskmax,
  input  [35:0] io_bp_0_control_reserved,
  input  [7:0] io_bp_0_control_bpaction,
  input  [3:0] io_bp_0_control_bpmatch,
  input   io_bp_0_control_m,
  input   io_bp_0_control_h,
  input   io_bp_0_control_s,
  input   io_bp_0_control_u,
  input   io_bp_0_control_r,
  input   io_bp_0_control_w,
  input   io_bp_0_control_x,
  input  [38:0] io_bp_0_address,
  input  [38:0] io_pc,
  input  [38:0] io_ea,
  output  io_xcpt_if,
  output  io_xcpt_ld,
  output  io_xcpt_st
);
  wire [1:0] T_176;
  wire [1:0] T_177;
  wire [3:0] T_178;
  wire [3:0] T_179;
  wire  T_180;
  wire [38:0] T_181;
  wire  T_182;
  wire  T_184;
  wire  T_185;
  wire [1:0] T_186;
  wire  T_187;
  wire  T_188;
  wire  T_189;
  wire [2:0] T_190;
  wire  T_191;
  wire  T_192;
  wire  T_193;
  wire [3:0] T_194;
  wire [38:0] GEN_6;
  wire [38:0] T_195;
  wire [38:0] T_196;
  wire [38:0] T_210;
  wire  T_211;
  wire  T_212;
  wire [38:0] T_214;
  wire [38:0] T_228;
  wire  T_244;
  wire  T_245;
  wire  T_278;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  assign io_xcpt_if = GEN_3;
  assign io_xcpt_ld = GEN_4;
  assign io_xcpt_st = GEN_5;
  assign T_176 = {io_bp_0_control_s,io_bp_0_control_u};
  assign T_177 = {io_bp_0_control_m,io_bp_0_control_h};
  assign T_178 = {T_177,T_176};
  assign T_179 = T_178 >> io_status_prv;
  assign T_180 = T_179[0];
  assign T_181 = ~ io_pc;
  assign T_182 = io_bp_0_control_bpmatch[1];
  assign T_184 = io_bp_0_address[0];
  assign T_185 = T_182 & T_184;
  assign T_186 = {T_185,T_182};
  assign T_187 = T_186[1];
  assign T_188 = io_bp_0_address[1];
  assign T_189 = T_187 & T_188;
  assign T_190 = {T_189,T_186};
  assign T_191 = T_190[2];
  assign T_192 = io_bp_0_address[2];
  assign T_193 = T_191 & T_192;
  assign T_194 = {T_193,T_190};
  assign GEN_6 = {{35'd0}, T_194};
  assign T_195 = T_181 | GEN_6;
  assign T_196 = ~ io_bp_0_address;
  assign T_210 = T_196 | GEN_6;
  assign T_211 = T_195 == T_210;
  assign T_212 = T_211 & io_bp_0_control_x;
  assign T_214 = ~ io_ea;
  assign T_228 = T_214 | GEN_6;
  assign T_244 = T_228 == T_210;
  assign T_245 = T_244 & io_bp_0_control_r;
  assign T_278 = T_244 & io_bp_0_control_w;
  assign GEN_3 = T_180 ? T_212 : 1'h0;
  assign GEN_4 = T_180 ? T_245 : 1'h0;
  assign GEN_5 = T_180 ? T_278 : 1'h0;
endmodule
module ALU(
  input   clk,
  input   reset,
  input   io_dw,
  input  [3:0] io_fn,
  input  [63:0] io_in2,
  input  [63:0] io_in1,
  output [63:0] io_out,
  output [63:0] io_adder_out,
  output  io_cmp_out
);
  wire  T_7;
  wire [63:0] T_8;
  wire [63:0] in2_inv;
  wire [63:0] in1_xor_in2;
  wire [64:0] T_9;
  wire [63:0] T_10;
  wire [63:0] GEN_1;
  wire [64:0] T_12;
  wire [63:0] T_13;
  wire  T_14;
  wire  T_17;
  wire [63:0] GEN_2;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire  T_29;
  wire  T_30;
  wire  T_32;
  wire  T_33;
  wire [31:0] GEN_3;
  wire [32:0] T_35;
  wire [31:0] T_36;
  wire [31:0] T_41;
  wire [31:0] T_42;
  wire  T_43;
  wire  T_48;
  wire [4:0] T_49;
  wire [5:0] shamt;
  wire [31:0] T_50;
  wire [63:0] shin_r;
  wire [3:0] GEN_4;
  wire  T_51;
  wire  T_52;
  wire  T_53;
  wire [31:0] T_58;
  wire [63:0] GEN_5;
  wire [63:0] T_59;
  wire [31:0] T_60;
  wire [63:0] GEN_6;
  wire [63:0] T_61;
  wire [63:0] T_63;
  wire [63:0] T_64;
  wire [47:0] T_68;
  wire [63:0] GEN_7;
  wire [63:0] T_69;
  wire [47:0] T_70;
  wire [63:0] GEN_8;
  wire [63:0] T_71;
  wire [63:0] T_73;
  wire [63:0] T_74;
  wire [55:0] T_78;
  wire [63:0] GEN_9;
  wire [63:0] T_79;
  wire [55:0] T_80;
  wire [63:0] GEN_10;
  wire [63:0] T_81;
  wire [63:0] T_83;
  wire [63:0] T_84;
  wire [59:0] T_88;
  wire [63:0] GEN_11;
  wire [63:0] T_89;
  wire [59:0] T_90;
  wire [63:0] GEN_12;
  wire [63:0] T_91;
  wire [63:0] T_93;
  wire [63:0] T_94;
  wire [61:0] T_98;
  wire [63:0] GEN_13;
  wire [63:0] T_99;
  wire [61:0] T_100;
  wire [63:0] GEN_14;
  wire [63:0] T_101;
  wire [63:0] T_103;
  wire [63:0] T_104;
  wire [62:0] T_108;
  wire [63:0] GEN_15;
  wire [63:0] T_109;
  wire [62:0] T_110;
  wire [63:0] GEN_16;
  wire [63:0] T_111;
  wire [63:0] T_113;
  wire [63:0] T_114;
  wire [63:0] shin;
  wire  T_116;
  wire  T_117;
  wire [64:0] T_118;
  wire [64:0] T_119;
  wire [64:0] T_120;
  wire [63:0] shout_r;
  wire [31:0] T_125;
  wire [63:0] GEN_17;
  wire [63:0] T_126;
  wire [31:0] T_127;
  wire [63:0] GEN_18;
  wire [63:0] T_128;
  wire [63:0] T_130;
  wire [63:0] T_131;
  wire [47:0] T_135;
  wire [63:0] GEN_19;
  wire [63:0] T_136;
  wire [47:0] T_137;
  wire [63:0] GEN_20;
  wire [63:0] T_138;
  wire [63:0] T_140;
  wire [63:0] T_141;
  wire [55:0] T_145;
  wire [63:0] GEN_21;
  wire [63:0] T_146;
  wire [55:0] T_147;
  wire [63:0] GEN_22;
  wire [63:0] T_148;
  wire [63:0] T_150;
  wire [63:0] T_151;
  wire [59:0] T_155;
  wire [63:0] GEN_23;
  wire [63:0] T_156;
  wire [59:0] T_157;
  wire [63:0] GEN_24;
  wire [63:0] T_158;
  wire [63:0] T_160;
  wire [63:0] T_161;
  wire [61:0] T_165;
  wire [63:0] GEN_25;
  wire [63:0] T_166;
  wire [61:0] T_167;
  wire [63:0] GEN_26;
  wire [63:0] T_168;
  wire [63:0] T_170;
  wire [63:0] T_171;
  wire [62:0] T_175;
  wire [63:0] GEN_27;
  wire [63:0] T_176;
  wire [62:0] T_177;
  wire [63:0] GEN_28;
  wire [63:0] T_178;
  wire [63:0] T_180;
  wire [63:0] shout_l;
  wire [63:0] T_185;
  wire [3:0] GEN_30;
  wire  T_186;
  wire [63:0] T_188;
  wire [63:0] shout;
  wire [3:0] GEN_31;
  wire  T_189;
  wire [3:0] GEN_32;
  wire  T_190;
  wire  T_191;
  wire [63:0] T_193;
  wire [3:0] GEN_34;
  wire  T_195;
  wire  T_196;
  wire [63:0] T_197;
  wire [63:0] T_199;
  wire [63:0] logic$;
  wire [3:0] GEN_35;
  wire  T_200;
  wire [3:0] GEN_36;
  wire  T_201;
  wire  T_202;
  wire  T_203;
  wire  T_204;
  wire  T_205;
  wire [63:0] GEN_37;
  wire [63:0] T_206;
  wire [63:0] shift_logic;
  wire [3:0] GEN_38;
  wire  T_207;
  wire  T_208;
  wire  T_209;
  wire [63:0] out;
  wire  T_213;
  wire  T_214;
  wire [31:0] GEN_39;
  wire [32:0] T_216;
  wire [31:0] T_217;
  wire [31:0] T_218;
  wire [63:0] T_219;
  wire [63:0] GEN_0;
  assign io_out = GEN_0;
  assign io_adder_out = T_13;
  assign io_cmp_out = T_30;
  assign T_7 = io_fn[3];
  assign T_8 = ~ io_in2;
  assign in2_inv = T_7 ? T_8 : io_in2;
  assign in1_xor_in2 = io_in1 ^ in2_inv;
  assign T_9 = io_in1 + in2_inv;
  assign T_10 = T_9[63:0];
  assign GEN_1 = {{63'd0}, T_7};
  assign T_12 = T_10 + GEN_1;
  assign T_13 = T_12[63:0];
  assign T_14 = io_fn[0];
  assign T_17 = T_7 == 1'h0;
  assign GEN_2 = {{63'd0}, 1'h0};
  assign T_19 = in1_xor_in2 == GEN_2;
  assign T_20 = io_in1[63];
  assign T_21 = io_in2[63];
  assign T_22 = T_20 == T_21;
  assign T_23 = io_adder_out[63];
  assign T_24 = io_fn[1];
  assign T_27 = T_24 ? T_21 : T_20;
  assign T_28 = T_22 ? T_23 : T_27;
  assign T_29 = T_17 ? T_19 : T_28;
  assign T_30 = T_14 ^ T_29;
  assign T_32 = io_in1[31];
  assign T_33 = T_7 & T_32;
  assign GEN_3 = {{31'd0}, T_33};
  assign T_35 = 32'h0 - GEN_3;
  assign T_36 = T_35[31:0];
  assign T_41 = io_in1[63:32];
  assign T_42 = io_dw ? T_41 : T_36;
  assign T_43 = io_in2[5];
  assign T_48 = T_43 & io_dw;
  assign T_49 = io_in2[4:0];
  assign shamt = {T_48,T_49};
  assign T_50 = io_in1[31:0];
  assign shin_r = {T_42,T_50};
  assign GEN_4 = {{1'd0}, 3'h5};
  assign T_51 = io_fn == GEN_4;
  assign T_52 = io_fn == 4'hb;
  assign T_53 = T_51 | T_52;
  assign T_58 = shin_r[63:32];
  assign GEN_5 = {{32'd0}, T_58};
  assign T_59 = GEN_5 & 64'hffffffff;
  assign T_60 = shin_r[31:0];
  assign GEN_6 = {{32'd0}, T_60};
  assign T_61 = GEN_6 << 32;
  assign T_63 = T_61 & 64'hffffffff00000000;
  assign T_64 = T_59 | T_63;
  assign T_68 = T_64[63:16];
  assign GEN_7 = {{16'd0}, T_68};
  assign T_69 = GEN_7 & 64'hffff0000ffff;
  assign T_70 = T_64[47:0];
  assign GEN_8 = {{16'd0}, T_70};
  assign T_71 = GEN_8 << 16;
  assign T_73 = T_71 & 64'hffff0000ffff0000;
  assign T_74 = T_69 | T_73;
  assign T_78 = T_74[63:8];
  assign GEN_9 = {{8'd0}, T_78};
  assign T_79 = GEN_9 & 64'hff00ff00ff00ff;
  assign T_80 = T_74[55:0];
  assign GEN_10 = {{8'd0}, T_80};
  assign T_81 = GEN_10 << 8;
  assign T_83 = T_81 & 64'hff00ff00ff00ff00;
  assign T_84 = T_79 | T_83;
  assign T_88 = T_84[63:4];
  assign GEN_11 = {{4'd0}, T_88};
  assign T_89 = GEN_11 & 64'hf0f0f0f0f0f0f0f;
  assign T_90 = T_84[59:0];
  assign GEN_12 = {{4'd0}, T_90};
  assign T_91 = GEN_12 << 4;
  assign T_93 = T_91 & 64'hf0f0f0f0f0f0f0f0;
  assign T_94 = T_89 | T_93;
  assign T_98 = T_94[63:2];
  assign GEN_13 = {{2'd0}, T_98};
  assign T_99 = GEN_13 & 64'h3333333333333333;
  assign T_100 = T_94[61:0];
  assign GEN_14 = {{2'd0}, T_100};
  assign T_101 = GEN_14 << 2;
  assign T_103 = T_101 & 64'hcccccccccccccccc;
  assign T_104 = T_99 | T_103;
  assign T_108 = T_104[63:1];
  assign GEN_15 = {{1'd0}, T_108};
  assign T_109 = GEN_15 & 64'h5555555555555555;
  assign T_110 = T_104[62:0];
  assign GEN_16 = {{1'd0}, T_110};
  assign T_111 = GEN_16 << 1;
  assign T_113 = T_111 & 64'haaaaaaaaaaaaaaaa;
  assign T_114 = T_109 | T_113;
  assign shin = T_53 ? shin_r : T_114;
  assign T_116 = shin[63];
  assign T_117 = T_7 & T_116;
  assign T_118 = {T_117,shin};
  assign T_119 = $signed(T_118);
  assign T_120 = $signed(T_119) >>> shamt;
  assign shout_r = T_120[63:0];
  assign T_125 = shout_r[63:32];
  assign GEN_17 = {{32'd0}, T_125};
  assign T_126 = GEN_17 & 64'hffffffff;
  assign T_127 = shout_r[31:0];
  assign GEN_18 = {{32'd0}, T_127};
  assign T_128 = GEN_18 << 32;
  assign T_130 = T_128 & 64'hffffffff00000000;
  assign T_131 = T_126 | T_130;
  assign T_135 = T_131[63:16];
  assign GEN_19 = {{16'd0}, T_135};
  assign T_136 = GEN_19 & 64'hffff0000ffff;
  assign T_137 = T_131[47:0];
  assign GEN_20 = {{16'd0}, T_137};
  assign T_138 = GEN_20 << 16;
  assign T_140 = T_138 & 64'hffff0000ffff0000;
  assign T_141 = T_136 | T_140;
  assign T_145 = T_141[63:8];
  assign GEN_21 = {{8'd0}, T_145};
  assign T_146 = GEN_21 & 64'hff00ff00ff00ff;
  assign T_147 = T_141[55:0];
  assign GEN_22 = {{8'd0}, T_147};
  assign T_148 = GEN_22 << 8;
  assign T_150 = T_148 & 64'hff00ff00ff00ff00;
  assign T_151 = T_146 | T_150;
  assign T_155 = T_151[63:4];
  assign GEN_23 = {{4'd0}, T_155};
  assign T_156 = GEN_23 & 64'hf0f0f0f0f0f0f0f;
  assign T_157 = T_151[59:0];
  assign GEN_24 = {{4'd0}, T_157};
  assign T_158 = GEN_24 << 4;
  assign T_160 = T_158 & 64'hf0f0f0f0f0f0f0f0;
  assign T_161 = T_156 | T_160;
  assign T_165 = T_161[63:2];
  assign GEN_25 = {{2'd0}, T_165};
  assign T_166 = GEN_25 & 64'h3333333333333333;
  assign T_167 = T_161[61:0];
  assign GEN_26 = {{2'd0}, T_167};
  assign T_168 = GEN_26 << 2;
  assign T_170 = T_168 & 64'hcccccccccccccccc;
  assign T_171 = T_166 | T_170;
  assign T_175 = T_171[63:1];
  assign GEN_27 = {{1'd0}, T_175};
  assign T_176 = GEN_27 & 64'h5555555555555555;
  assign T_177 = T_171[62:0];
  assign GEN_28 = {{1'd0}, T_177};
  assign T_178 = GEN_28 << 1;
  assign T_180 = T_178 & 64'haaaaaaaaaaaaaaaa;
  assign shout_l = T_176 | T_180;
  assign T_185 = T_53 ? shout_r : {{63'd0}, 1'h0};
  assign GEN_30 = {{3'd0}, 1'h1};
  assign T_186 = io_fn == GEN_30;
  assign T_188 = T_186 ? shout_l : {{63'd0}, 1'h0};
  assign shout = T_185 | T_188;
  assign GEN_31 = {{1'd0}, 3'h4};
  assign T_189 = io_fn == GEN_31;
  assign GEN_32 = {{1'd0}, 3'h6};
  assign T_190 = io_fn == GEN_32;
  assign T_191 = T_189 | T_190;
  assign T_193 = T_191 ? in1_xor_in2 : {{63'd0}, 1'h0};
  assign GEN_34 = {{1'd0}, 3'h7};
  assign T_195 = io_fn == GEN_34;
  assign T_196 = T_190 | T_195;
  assign T_197 = io_in1 & io_in2;
  assign T_199 = T_196 ? T_197 : {{63'd0}, 1'h0};
  assign logic$ = T_193 | T_199;
  assign GEN_35 = {{2'd0}, 2'h2};
  assign T_200 = io_fn == GEN_35;
  assign GEN_36 = {{2'd0}, 2'h3};
  assign T_201 = io_fn == GEN_36;
  assign T_202 = T_200 | T_201;
  assign T_203 = io_fn >= 4'hc;
  assign T_204 = T_202 | T_203;
  assign T_205 = T_204 & io_cmp_out;
  assign GEN_37 = {{63'd0}, T_205};
  assign T_206 = GEN_37 | logic$;
  assign shift_logic = T_206 | shout;
  assign GEN_38 = {{3'd0}, 1'h0};
  assign T_207 = io_fn == GEN_38;
  assign T_208 = io_fn == 4'ha;
  assign T_209 = T_207 | T_208;
  assign out = T_209 ? io_adder_out : shift_logic;
  assign T_213 = 1'h0 == io_dw;
  assign T_214 = out[31];
  assign GEN_39 = {{31'd0}, T_214};
  assign T_216 = 32'h0 - GEN_39;
  assign T_217 = T_216[31:0];
  assign T_218 = out[31:0];
  assign T_219 = {T_217,T_218};
  assign GEN_0 = T_213 ? T_219 : out;
endmodule
module MulDiv(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [3:0] io_req_bits_fn,
  input   io_req_bits_dw,
  input  [63:0] io_req_bits_in1,
  input  [63:0] io_req_bits_in2,
  input  [4:0] io_req_bits_tag,
  input   io_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [63:0] io_resp_bits_data,
  output [4:0] io_resp_bits_tag
);
  reg [2:0] state;
  reg [31:0] GEN_43;
  reg [3:0] req_fn;
  reg [31:0] GEN_44;
  reg  req_dw;
  reg [31:0] GEN_47;
  reg [63:0] req_in1;
  reg [63:0] GEN_48;
  reg [63:0] req_in2;
  reg [63:0] GEN_49;
  reg [4:0] req_tag;
  reg [31:0] GEN_52;
  reg [6:0] count;
  reg [31:0] GEN_54;
  reg  neg_out;
  reg [31:0] GEN_55;
  reg  isMul;
  reg [31:0] GEN_56;
  reg  isHi;
  reg [31:0] GEN_57;
  reg [64:0] divisor;
  reg [95:0] GEN_58;
  reg [129:0] remainder;
  reg [159:0] GEN_59;
  wire [3:0] T_62;
  wire  T_64;
  wire [3:0] T_66;
  wire  T_68;
  wire  T_71;
  wire [3:0] T_73;
  wire  T_75;
  wire [3:0] T_77;
  wire  T_79;
  wire  T_82;
  wire  T_83;
  wire [3:0] T_85;
  wire  T_87;
  wire [3:0] T_89;
  wire  T_91;
  wire  T_94;
  wire  T_95;
  wire  T_103;
  wire  T_105;
  wire  T_106;
  wire  T_107;
  wire  lhs_sign;
  wire [31:0] GEN_34;
  wire [32:0] T_109;
  wire [31:0] T_110;
  wire [31:0] T_111;
  wire [31:0] T_112;
  wire [31:0] T_113;
  wire [63:0] lhs_in;
  wire  T_120;
  wire  T_121;
  wire  T_122;
  wire  rhs_sign;
  wire [31:0] GEN_35;
  wire [32:0] T_124;
  wire [31:0] T_125;
  wire [31:0] T_126;
  wire [31:0] T_127;
  wire [31:0] T_128;
  wire [63:0] rhs_in;
  wire [64:0] T_129;
  wire [65:0] T_131;
  wire [64:0] subtractor;
  wire  less;
  wire [63:0] T_132;
  wire [63:0] GEN_36;
  wire [64:0] T_134;
  wire [63:0] negated_remainder;
  wire  T_135;
  wire  T_136;
  wire  T_137;
  wire [129:0] GEN_0;
  wire  T_138;
  wire  T_139;
  wire [64:0] GEN_1;
  wire [129:0] GEN_2;
  wire [64:0] GEN_3;
  wire [2:0] GEN_4;
  wire  T_140;
  wire [129:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_141;
  wire [63:0] T_142;
  wire [2:0] T_143;
  wire [129:0] GEN_7;
  wire [2:0] GEN_8;
  wire  T_144;
  wire  T_145;
  wire [64:0] T_146;
  wire [128:0] T_148;
  wire [63:0] T_149;
  wire [64:0] T_150;
  wire [64:0] T_151;
  wire [64:0] T_152;
  wire [7:0] T_153;
  wire [64:0] GEN_37;
  wire [72:0] T_154;
  wire [72:0] GEN_38;
  wire [73:0] T_155;
  wire [72:0] T_156;
  wire [72:0] T_157;
  wire [55:0] T_158;
  wire [72:0] T_159;
  wire [128:0] T_160;
  wire [6:0] GEN_39;
  wire [10:0] T_163;
  wire [5:0] T_164;
  wire [64:0] GEN_40;
  wire [64:0] T_165;
  wire [63:0] T_166;
  wire [6:0] GEN_41;
  wire  T_169;
  wire [6:0] GEN_42;
  wire  T_172;
  wire  T_173;
  wire  T_175;
  wire  T_176;
  wire [63:0] T_177;
  wire [63:0] T_178;
  wire  T_180;
  wire  T_181;
  wire [10:0] GEN_45;
  wire [11:0] T_185;
  wire [10:0] T_186;
  wire [5:0] T_187;
  wire [128:0] T_188;
  wire [64:0] T_189;
  wire [128:0] T_190;
  wire [63:0] T_191;
  wire [128:0] T_192;
  wire [64:0] T_193;
  wire [63:0] T_195;
  wire [65:0] T_196;
  wire [129:0] T_197;
  wire [6:0] GEN_46;
  wire [7:0] T_199;
  wire [6:0] T_200;
  wire  T_202;
  wire  T_203;
  wire [2:0] T_204;
  wire [2:0] GEN_9;
  wire [129:0] GEN_10;
  wire [6:0] GEN_11;
  wire [2:0] GEN_12;
  wire  T_207;
  wire  T_208;
  wire  T_210;
  wire [2:0] T_212;
  wire [2:0] GEN_13;
  wire [63:0] T_216;
  wire [63:0] T_217;
  wire [63:0] T_218;
  wire  T_221;
  wire [127:0] T_222;
  wire [128:0] T_223;
  wire [63:0] T_224;
  wire  T_225;
  wire  T_227;
  wire  T_229;
  wire  T_231;
  wire  T_233;
  wire  T_235;
  wire  T_237;
  wire  T_239;
  wire  T_241;
  wire  T_243;
  wire  T_245;
  wire  T_247;
  wire  T_249;
  wire  T_251;
  wire  T_253;
  wire  T_255;
  wire  T_257;
  wire  T_259;
  wire  T_261;
  wire  T_263;
  wire  T_265;
  wire  T_267;
  wire  T_269;
  wire  T_271;
  wire  T_273;
  wire  T_275;
  wire  T_277;
  wire  T_279;
  wire  T_281;
  wire  T_283;
  wire  T_285;
  wire  T_287;
  wire  T_289;
  wire  T_291;
  wire  T_293;
  wire  T_295;
  wire  T_297;
  wire  T_299;
  wire  T_301;
  wire  T_303;
  wire  T_305;
  wire  T_307;
  wire  T_309;
  wire  T_311;
  wire  T_313;
  wire  T_315;
  wire  T_317;
  wire  T_319;
  wire  T_321;
  wire  T_323;
  wire  T_325;
  wire  T_327;
  wire  T_329;
  wire  T_331;
  wire  T_333;
  wire  T_335;
  wire  T_337;
  wire  T_339;
  wire  T_341;
  wire  T_343;
  wire  T_345;
  wire  T_347;
  wire  T_349;
  wire [1:0] T_351;
  wire [1:0] T_352;
  wire [2:0] T_353;
  wire [2:0] T_354;
  wire [2:0] T_355;
  wire [2:0] T_356;
  wire [3:0] T_357;
  wire [3:0] T_358;
  wire [3:0] T_359;
  wire [3:0] T_360;
  wire [3:0] T_361;
  wire [3:0] T_362;
  wire [3:0] T_363;
  wire [3:0] T_364;
  wire [4:0] T_365;
  wire [4:0] T_366;
  wire [4:0] T_367;
  wire [4:0] T_368;
  wire [4:0] T_369;
  wire [4:0] T_370;
  wire [4:0] T_371;
  wire [4:0] T_372;
  wire [4:0] T_373;
  wire [4:0] T_374;
  wire [4:0] T_375;
  wire [4:0] T_376;
  wire [4:0] T_377;
  wire [4:0] T_378;
  wire [4:0] T_379;
  wire [4:0] T_380;
  wire [5:0] T_381;
  wire [5:0] T_382;
  wire [5:0] T_383;
  wire [5:0] T_384;
  wire [5:0] T_385;
  wire [5:0] T_386;
  wire [5:0] T_387;
  wire [5:0] T_388;
  wire [5:0] T_389;
  wire [5:0] T_390;
  wire [5:0] T_391;
  wire [5:0] T_392;
  wire [5:0] T_393;
  wire [5:0] T_394;
  wire [5:0] T_395;
  wire [5:0] T_396;
  wire [5:0] T_397;
  wire [5:0] T_398;
  wire [5:0] T_399;
  wire [5:0] T_400;
  wire [5:0] T_401;
  wire [5:0] T_402;
  wire [5:0] T_403;
  wire [5:0] T_404;
  wire [5:0] T_405;
  wire [5:0] T_406;
  wire [5:0] T_407;
  wire [5:0] T_408;
  wire [5:0] T_409;
  wire [5:0] T_410;
  wire [5:0] T_411;
  wire [5:0] T_412;
  wire  T_414;
  wire  T_416;
  wire  T_418;
  wire  T_420;
  wire  T_422;
  wire  T_424;
  wire  T_426;
  wire  T_428;
  wire  T_430;
  wire  T_432;
  wire  T_434;
  wire  T_436;
  wire  T_438;
  wire  T_440;
  wire  T_442;
  wire  T_444;
  wire  T_446;
  wire  T_448;
  wire  T_450;
  wire  T_452;
  wire  T_454;
  wire  T_456;
  wire  T_458;
  wire  T_460;
  wire  T_462;
  wire  T_464;
  wire  T_466;
  wire  T_468;
  wire  T_470;
  wire  T_472;
  wire  T_474;
  wire  T_476;
  wire  T_478;
  wire  T_480;
  wire  T_482;
  wire  T_484;
  wire  T_486;
  wire  T_488;
  wire  T_490;
  wire  T_492;
  wire  T_494;
  wire  T_496;
  wire  T_498;
  wire  T_500;
  wire  T_502;
  wire  T_504;
  wire  T_506;
  wire  T_508;
  wire  T_510;
  wire  T_512;
  wire  T_514;
  wire  T_516;
  wire  T_518;
  wire  T_520;
  wire  T_522;
  wire  T_524;
  wire  T_526;
  wire  T_528;
  wire  T_530;
  wire  T_532;
  wire  T_534;
  wire  T_536;
  wire  T_538;
  wire [1:0] T_540;
  wire [1:0] T_541;
  wire [2:0] T_542;
  wire [2:0] T_543;
  wire [2:0] T_544;
  wire [2:0] T_545;
  wire [3:0] T_546;
  wire [3:0] T_547;
  wire [3:0] T_548;
  wire [3:0] T_549;
  wire [3:0] T_550;
  wire [3:0] T_551;
  wire [3:0] T_552;
  wire [3:0] T_553;
  wire [4:0] T_554;
  wire [4:0] T_555;
  wire [4:0] T_556;
  wire [4:0] T_557;
  wire [4:0] T_558;
  wire [4:0] T_559;
  wire [4:0] T_560;
  wire [4:0] T_561;
  wire [4:0] T_562;
  wire [4:0] T_563;
  wire [4:0] T_564;
  wire [4:0] T_565;
  wire [4:0] T_566;
  wire [4:0] T_567;
  wire [4:0] T_568;
  wire [4:0] T_569;
  wire [5:0] T_570;
  wire [5:0] T_571;
  wire [5:0] T_572;
  wire [5:0] T_573;
  wire [5:0] T_574;
  wire [5:0] T_575;
  wire [5:0] T_576;
  wire [5:0] T_577;
  wire [5:0] T_578;
  wire [5:0] T_579;
  wire [5:0] T_580;
  wire [5:0] T_581;
  wire [5:0] T_582;
  wire [5:0] T_583;
  wire [5:0] T_584;
  wire [5:0] T_585;
  wire [5:0] T_586;
  wire [5:0] T_587;
  wire [5:0] T_588;
  wire [5:0] T_589;
  wire [5:0] T_590;
  wire [5:0] T_591;
  wire [5:0] T_592;
  wire [5:0] T_593;
  wire [5:0] T_594;
  wire [5:0] T_595;
  wire [5:0] T_596;
  wire [5:0] T_597;
  wire [5:0] T_598;
  wire [5:0] T_599;
  wire [5:0] T_600;
  wire [5:0] T_601;
  wire [6:0] T_603;
  wire [5:0] T_604;
  wire [6:0] T_605;
  wire [5:0] T_606;
  wire  T_607;
  wire  T_609;
  wire  T_610;
  wire [5:0] GEN_50;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire [5:0] T_619;
  wire [126:0] GEN_51;
  wire [126:0] T_621;
  wire [128:0] GEN_14;
  wire [6:0] GEN_15;
  wire  T_626;
  wire  T_629;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [6:0] GEN_18;
  wire [129:0] GEN_19;
  wire  GEN_20;
  wire  T_631;
  wire  T_632;
  wire [2:0] GEN_21;
  wire  T_633;
  wire  T_635;
  wire  T_636;
  wire  T_637;
  wire [2:0] T_638;
  wire  T_642;
  wire  T_643;
  wire  T_644;
  wire [64:0] T_645;
  wire [2:0] GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire [6:0] GEN_25;
  wire  GEN_26;
  wire [64:0] GEN_27;
  wire [129:0] GEN_28;
  wire [3:0] GEN_29;
  wire  GEN_30;
  wire [63:0] GEN_31;
  wire [63:0] GEN_32;
  wire [4:0] GEN_33;
  wire  T_650;
  wire  T_652;
  wire [31:0] GEN_53;
  wire [32:0] T_654;
  wire [31:0] T_655;
  wire [31:0] T_656;
  wire [63:0] T_657;
  wire [63:0] T_659;
  wire  T_660;
  wire  T_661;
  assign io_req_ready = T_661;
  assign io_resp_valid = T_660;
  assign io_resp_bits_data = T_659;
  assign io_resp_bits_tag = req_tag;
  assign T_62 = io_req_bits_fn & 4'h4;
  assign T_64 = T_62 == 4'h0;
  assign T_66 = io_req_bits_fn & 4'h8;
  assign T_68 = T_66 == 4'h8;
  assign T_71 = T_64 | T_68;
  assign T_73 = io_req_bits_fn & 4'h5;
  assign T_75 = T_73 == 4'h1;
  assign T_77 = io_req_bits_fn & 4'h2;
  assign T_79 = T_77 == 4'h2;
  assign T_82 = T_75 | T_79;
  assign T_83 = T_82 | T_68;
  assign T_85 = io_req_bits_fn & 4'h9;
  assign T_87 = T_85 == 4'h0;
  assign T_89 = io_req_bits_fn & 4'h3;
  assign T_91 = T_89 == 4'h0;
  assign T_94 = T_87 | T_64;
  assign T_95 = T_94 | T_91;
  assign T_103 = 1'h0 == io_req_bits_dw;
  assign T_105 = io_req_bits_in1[31];
  assign T_106 = io_req_bits_in1[63];
  assign T_107 = T_103 ? T_105 : T_106;
  assign lhs_sign = T_95 & T_107;
  assign GEN_34 = {{31'd0}, lhs_sign};
  assign T_109 = 32'h0 - GEN_34;
  assign T_110 = T_109[31:0];
  assign T_111 = io_req_bits_in1[63:32];
  assign T_112 = T_103 ? T_110 : T_111;
  assign T_113 = io_req_bits_in1[31:0];
  assign lhs_in = {T_112,T_113};
  assign T_120 = io_req_bits_in2[31];
  assign T_121 = io_req_bits_in2[63];
  assign T_122 = T_103 ? T_120 : T_121;
  assign rhs_sign = T_94 & T_122;
  assign GEN_35 = {{31'd0}, rhs_sign};
  assign T_124 = 32'h0 - GEN_35;
  assign T_125 = T_124[31:0];
  assign T_126 = io_req_bits_in2[63:32];
  assign T_127 = T_103 ? T_125 : T_126;
  assign T_128 = io_req_bits_in2[31:0];
  assign rhs_in = {T_127,T_128};
  assign T_129 = remainder[128:64];
  assign T_131 = T_129 - divisor;
  assign subtractor = T_131[64:0];
  assign less = subtractor[64];
  assign T_132 = remainder[63:0];
  assign GEN_36 = {{63'd0}, 1'h0};
  assign T_134 = GEN_36 - T_132;
  assign negated_remainder = T_134[63:0];
  assign T_135 = state == 3'h1;
  assign T_136 = remainder[63];
  assign T_137 = T_136 | isMul;
  assign GEN_0 = T_137 ? {{66'd0}, negated_remainder} : remainder;
  assign T_138 = divisor[63];
  assign T_139 = T_138 | isMul;
  assign GEN_1 = T_139 ? subtractor : divisor;
  assign GEN_2 = T_135 ? GEN_0 : remainder;
  assign GEN_3 = T_135 ? GEN_1 : divisor;
  assign GEN_4 = T_135 ? 3'h2 : state;
  assign T_140 = state == 3'h4;
  assign GEN_5 = T_140 ? {{66'd0}, negated_remainder} : GEN_2;
  assign GEN_6 = T_140 ? 3'h5 : GEN_4;
  assign T_141 = state == 3'h3;
  assign T_142 = remainder[128:65];
  assign T_143 = neg_out ? 3'h4 : 3'h5;
  assign GEN_7 = T_141 ? {{66'd0}, T_142} : GEN_5;
  assign GEN_8 = T_141 ? T_143 : GEN_6;
  assign T_144 = state == 3'h2;
  assign T_145 = T_144 & isMul;
  assign T_146 = remainder[129:65];
  assign T_148 = {T_146,T_132};
  assign T_149 = T_148[63:0];
  assign T_150 = T_148[128:64];
  assign T_151 = $signed(T_150);
  assign T_152 = $signed(divisor);
  assign T_153 = T_149[7:0];
  assign GEN_37 = {{57'd0}, T_153};
  assign T_154 = $signed(T_152) * $signed({1'b0,GEN_37});
  assign GEN_38 = {{8{T_151[64]}},T_151};
  assign T_155 = $signed(T_154) + $signed(GEN_38);
  assign T_156 = T_155[72:0];
  assign T_157 = $signed(T_156);
  assign T_158 = T_149[63:8];
  assign T_159 = $unsigned(T_157);
  assign T_160 = {T_159,T_158};
  assign GEN_39 = {{3'd0}, 4'h8};
  assign T_163 = count * GEN_39;
  assign T_164 = T_163[5:0];
  assign GEN_40 = $signed(65'h10000000000000000);
  assign T_165 = $signed(GEN_40) >>> T_164;
  assign T_166 = T_165[63:0];
  assign GEN_41 = {{4'd0}, 3'h7};
  assign T_169 = count != GEN_41;
  assign GEN_42 = {{6'd0}, 1'h0};
  assign T_172 = count != GEN_42;
  assign T_173 = T_169 & T_172;
  assign T_175 = isHi == 1'h0;
  assign T_176 = T_173 & T_175;
  assign T_177 = ~ T_166;
  assign T_178 = T_149 & T_177;
  assign T_180 = T_178 == GEN_36;
  assign T_181 = T_176 & T_180;
  assign GEN_45 = {{4'd0}, 7'h40};
  assign T_185 = GEN_45 - T_163;
  assign T_186 = T_185[10:0];
  assign T_187 = T_186[5:0];
  assign T_188 = T_148 >> T_187;
  assign T_189 = T_160[128:64];
  assign T_190 = T_181 ? T_188 : T_160;
  assign T_191 = T_190[63:0];
  assign T_192 = {T_189,T_191};
  assign T_193 = T_192[128:64];
  assign T_195 = T_192[63:0];
  assign T_196 = {T_193,1'h0};
  assign T_197 = {T_196,T_195};
  assign GEN_46 = {{6'd0}, 1'h1};
  assign T_199 = count + GEN_46;
  assign T_200 = T_199[6:0];
  assign T_202 = count == GEN_41;
  assign T_203 = T_181 | T_202;
  assign T_204 = isHi ? 3'h3 : 3'h5;
  assign GEN_9 = T_203 ? T_204 : GEN_8;
  assign GEN_10 = T_145 ? T_197 : GEN_7;
  assign GEN_11 = T_145 ? T_200 : count;
  assign GEN_12 = T_145 ? GEN_9 : GEN_8;
  assign T_207 = isMul == 1'h0;
  assign T_208 = T_144 & T_207;
  assign T_210 = count == 7'h40;
  assign T_212 = isHi ? 3'h3 : T_143;
  assign GEN_13 = T_210 ? T_212 : GEN_12;
  assign T_216 = remainder[127:64];
  assign T_217 = subtractor[63:0];
  assign T_218 = less ? T_216 : T_217;
  assign T_221 = less == 1'h0;
  assign T_222 = {T_218,T_132};
  assign T_223 = {T_222,T_221};
  assign T_224 = divisor[63:0];
  assign T_225 = T_224[63];
  assign T_227 = T_224[62];
  assign T_229 = T_224[61];
  assign T_231 = T_224[60];
  assign T_233 = T_224[59];
  assign T_235 = T_224[58];
  assign T_237 = T_224[57];
  assign T_239 = T_224[56];
  assign T_241 = T_224[55];
  assign T_243 = T_224[54];
  assign T_245 = T_224[53];
  assign T_247 = T_224[52];
  assign T_249 = T_224[51];
  assign T_251 = T_224[50];
  assign T_253 = T_224[49];
  assign T_255 = T_224[48];
  assign T_257 = T_224[47];
  assign T_259 = T_224[46];
  assign T_261 = T_224[45];
  assign T_263 = T_224[44];
  assign T_265 = T_224[43];
  assign T_267 = T_224[42];
  assign T_269 = T_224[41];
  assign T_271 = T_224[40];
  assign T_273 = T_224[39];
  assign T_275 = T_224[38];
  assign T_277 = T_224[37];
  assign T_279 = T_224[36];
  assign T_281 = T_224[35];
  assign T_283 = T_224[34];
  assign T_285 = T_224[33];
  assign T_287 = T_224[32];
  assign T_289 = T_224[31];
  assign T_291 = T_224[30];
  assign T_293 = T_224[29];
  assign T_295 = T_224[28];
  assign T_297 = T_224[27];
  assign T_299 = T_224[26];
  assign T_301 = T_224[25];
  assign T_303 = T_224[24];
  assign T_305 = T_224[23];
  assign T_307 = T_224[22];
  assign T_309 = T_224[21];
  assign T_311 = T_224[20];
  assign T_313 = T_224[19];
  assign T_315 = T_224[18];
  assign T_317 = T_224[17];
  assign T_319 = T_224[16];
  assign T_321 = T_224[15];
  assign T_323 = T_224[14];
  assign T_325 = T_224[13];
  assign T_327 = T_224[12];
  assign T_329 = T_224[11];
  assign T_331 = T_224[10];
  assign T_333 = T_224[9];
  assign T_335 = T_224[8];
  assign T_337 = T_224[7];
  assign T_339 = T_224[6];
  assign T_341 = T_224[5];
  assign T_343 = T_224[4];
  assign T_345 = T_224[3];
  assign T_347 = T_224[2];
  assign T_349 = T_224[1];
  assign T_351 = T_347 ? 2'h2 : {{1'd0}, T_349};
  assign T_352 = T_345 ? 2'h3 : T_351;
  assign T_353 = T_343 ? 3'h4 : {{1'd0}, T_352};
  assign T_354 = T_341 ? 3'h5 : T_353;
  assign T_355 = T_339 ? 3'h6 : T_354;
  assign T_356 = T_337 ? 3'h7 : T_355;
  assign T_357 = T_335 ? 4'h8 : {{1'd0}, T_356};
  assign T_358 = T_333 ? 4'h9 : T_357;
  assign T_359 = T_331 ? 4'ha : T_358;
  assign T_360 = T_329 ? 4'hb : T_359;
  assign T_361 = T_327 ? 4'hc : T_360;
  assign T_362 = T_325 ? 4'hd : T_361;
  assign T_363 = T_323 ? 4'he : T_362;
  assign T_364 = T_321 ? 4'hf : T_363;
  assign T_365 = T_319 ? 5'h10 : {{1'd0}, T_364};
  assign T_366 = T_317 ? 5'h11 : T_365;
  assign T_367 = T_315 ? 5'h12 : T_366;
  assign T_368 = T_313 ? 5'h13 : T_367;
  assign T_369 = T_311 ? 5'h14 : T_368;
  assign T_370 = T_309 ? 5'h15 : T_369;
  assign T_371 = T_307 ? 5'h16 : T_370;
  assign T_372 = T_305 ? 5'h17 : T_371;
  assign T_373 = T_303 ? 5'h18 : T_372;
  assign T_374 = T_301 ? 5'h19 : T_373;
  assign T_375 = T_299 ? 5'h1a : T_374;
  assign T_376 = T_297 ? 5'h1b : T_375;
  assign T_377 = T_295 ? 5'h1c : T_376;
  assign T_378 = T_293 ? 5'h1d : T_377;
  assign T_379 = T_291 ? 5'h1e : T_378;
  assign T_380 = T_289 ? 5'h1f : T_379;
  assign T_381 = T_287 ? 6'h20 : {{1'd0}, T_380};
  assign T_382 = T_285 ? 6'h21 : T_381;
  assign T_383 = T_283 ? 6'h22 : T_382;
  assign T_384 = T_281 ? 6'h23 : T_383;
  assign T_385 = T_279 ? 6'h24 : T_384;
  assign T_386 = T_277 ? 6'h25 : T_385;
  assign T_387 = T_275 ? 6'h26 : T_386;
  assign T_388 = T_273 ? 6'h27 : T_387;
  assign T_389 = T_271 ? 6'h28 : T_388;
  assign T_390 = T_269 ? 6'h29 : T_389;
  assign T_391 = T_267 ? 6'h2a : T_390;
  assign T_392 = T_265 ? 6'h2b : T_391;
  assign T_393 = T_263 ? 6'h2c : T_392;
  assign T_394 = T_261 ? 6'h2d : T_393;
  assign T_395 = T_259 ? 6'h2e : T_394;
  assign T_396 = T_257 ? 6'h2f : T_395;
  assign T_397 = T_255 ? 6'h30 : T_396;
  assign T_398 = T_253 ? 6'h31 : T_397;
  assign T_399 = T_251 ? 6'h32 : T_398;
  assign T_400 = T_249 ? 6'h33 : T_399;
  assign T_401 = T_247 ? 6'h34 : T_400;
  assign T_402 = T_245 ? 6'h35 : T_401;
  assign T_403 = T_243 ? 6'h36 : T_402;
  assign T_404 = T_241 ? 6'h37 : T_403;
  assign T_405 = T_239 ? 6'h38 : T_404;
  assign T_406 = T_237 ? 6'h39 : T_405;
  assign T_407 = T_235 ? 6'h3a : T_406;
  assign T_408 = T_233 ? 6'h3b : T_407;
  assign T_409 = T_231 ? 6'h3c : T_408;
  assign T_410 = T_229 ? 6'h3d : T_409;
  assign T_411 = T_227 ? 6'h3e : T_410;
  assign T_412 = T_225 ? 6'h3f : T_411;
  assign T_414 = T_132[63];
  assign T_416 = T_132[62];
  assign T_418 = T_132[61];
  assign T_420 = T_132[60];
  assign T_422 = T_132[59];
  assign T_424 = T_132[58];
  assign T_426 = T_132[57];
  assign T_428 = T_132[56];
  assign T_430 = T_132[55];
  assign T_432 = T_132[54];
  assign T_434 = T_132[53];
  assign T_436 = T_132[52];
  assign T_438 = T_132[51];
  assign T_440 = T_132[50];
  assign T_442 = T_132[49];
  assign T_444 = T_132[48];
  assign T_446 = T_132[47];
  assign T_448 = T_132[46];
  assign T_450 = T_132[45];
  assign T_452 = T_132[44];
  assign T_454 = T_132[43];
  assign T_456 = T_132[42];
  assign T_458 = T_132[41];
  assign T_460 = T_132[40];
  assign T_462 = T_132[39];
  assign T_464 = T_132[38];
  assign T_466 = T_132[37];
  assign T_468 = T_132[36];
  assign T_470 = T_132[35];
  assign T_472 = T_132[34];
  assign T_474 = T_132[33];
  assign T_476 = T_132[32];
  assign T_478 = T_132[31];
  assign T_480 = T_132[30];
  assign T_482 = T_132[29];
  assign T_484 = T_132[28];
  assign T_486 = T_132[27];
  assign T_488 = T_132[26];
  assign T_490 = T_132[25];
  assign T_492 = T_132[24];
  assign T_494 = T_132[23];
  assign T_496 = T_132[22];
  assign T_498 = T_132[21];
  assign T_500 = T_132[20];
  assign T_502 = T_132[19];
  assign T_504 = T_132[18];
  assign T_506 = T_132[17];
  assign T_508 = T_132[16];
  assign T_510 = T_132[15];
  assign T_512 = T_132[14];
  assign T_514 = T_132[13];
  assign T_516 = T_132[12];
  assign T_518 = T_132[11];
  assign T_520 = T_132[10];
  assign T_522 = T_132[9];
  assign T_524 = T_132[8];
  assign T_526 = T_132[7];
  assign T_528 = T_132[6];
  assign T_530 = T_132[5];
  assign T_532 = T_132[4];
  assign T_534 = T_132[3];
  assign T_536 = T_132[2];
  assign T_538 = T_132[1];
  assign T_540 = T_536 ? 2'h2 : {{1'd0}, T_538};
  assign T_541 = T_534 ? 2'h3 : T_540;
  assign T_542 = T_532 ? 3'h4 : {{1'd0}, T_541};
  assign T_543 = T_530 ? 3'h5 : T_542;
  assign T_544 = T_528 ? 3'h6 : T_543;
  assign T_545 = T_526 ? 3'h7 : T_544;
  assign T_546 = T_524 ? 4'h8 : {{1'd0}, T_545};
  assign T_547 = T_522 ? 4'h9 : T_546;
  assign T_548 = T_520 ? 4'ha : T_547;
  assign T_549 = T_518 ? 4'hb : T_548;
  assign T_550 = T_516 ? 4'hc : T_549;
  assign T_551 = T_514 ? 4'hd : T_550;
  assign T_552 = T_512 ? 4'he : T_551;
  assign T_553 = T_510 ? 4'hf : T_552;
  assign T_554 = T_508 ? 5'h10 : {{1'd0}, T_553};
  assign T_555 = T_506 ? 5'h11 : T_554;
  assign T_556 = T_504 ? 5'h12 : T_555;
  assign T_557 = T_502 ? 5'h13 : T_556;
  assign T_558 = T_500 ? 5'h14 : T_557;
  assign T_559 = T_498 ? 5'h15 : T_558;
  assign T_560 = T_496 ? 5'h16 : T_559;
  assign T_561 = T_494 ? 5'h17 : T_560;
  assign T_562 = T_492 ? 5'h18 : T_561;
  assign T_563 = T_490 ? 5'h19 : T_562;
  assign T_564 = T_488 ? 5'h1a : T_563;
  assign T_565 = T_486 ? 5'h1b : T_564;
  assign T_566 = T_484 ? 5'h1c : T_565;
  assign T_567 = T_482 ? 5'h1d : T_566;
  assign T_568 = T_480 ? 5'h1e : T_567;
  assign T_569 = T_478 ? 5'h1f : T_568;
  assign T_570 = T_476 ? 6'h20 : {{1'd0}, T_569};
  assign T_571 = T_474 ? 6'h21 : T_570;
  assign T_572 = T_472 ? 6'h22 : T_571;
  assign T_573 = T_470 ? 6'h23 : T_572;
  assign T_574 = T_468 ? 6'h24 : T_573;
  assign T_575 = T_466 ? 6'h25 : T_574;
  assign T_576 = T_464 ? 6'h26 : T_575;
  assign T_577 = T_462 ? 6'h27 : T_576;
  assign T_578 = T_460 ? 6'h28 : T_577;
  assign T_579 = T_458 ? 6'h29 : T_578;
  assign T_580 = T_456 ? 6'h2a : T_579;
  assign T_581 = T_454 ? 6'h2b : T_580;
  assign T_582 = T_452 ? 6'h2c : T_581;
  assign T_583 = T_450 ? 6'h2d : T_582;
  assign T_584 = T_448 ? 6'h2e : T_583;
  assign T_585 = T_446 ? 6'h2f : T_584;
  assign T_586 = T_444 ? 6'h30 : T_585;
  assign T_587 = T_442 ? 6'h31 : T_586;
  assign T_588 = T_440 ? 6'h32 : T_587;
  assign T_589 = T_438 ? 6'h33 : T_588;
  assign T_590 = T_436 ? 6'h34 : T_589;
  assign T_591 = T_434 ? 6'h35 : T_590;
  assign T_592 = T_432 ? 6'h36 : T_591;
  assign T_593 = T_430 ? 6'h37 : T_592;
  assign T_594 = T_428 ? 6'h38 : T_593;
  assign T_595 = T_426 ? 6'h39 : T_594;
  assign T_596 = T_424 ? 6'h3a : T_595;
  assign T_597 = T_422 ? 6'h3b : T_596;
  assign T_598 = T_420 ? 6'h3c : T_597;
  assign T_599 = T_418 ? 6'h3d : T_598;
  assign T_600 = T_416 ? 6'h3e : T_599;
  assign T_601 = T_414 ? 6'h3f : T_600;
  assign T_603 = 6'h3f + T_412;
  assign T_604 = T_603[5:0];
  assign T_605 = T_604 - T_601;
  assign T_606 = T_605[5:0];
  assign T_607 = T_412 > T_601;
  assign T_609 = count == GEN_42;
  assign T_610 = T_609 & less;
  assign GEN_50 = {{5'd0}, 1'h0};
  assign T_612 = T_606 > GEN_50;
  assign T_613 = T_612 | T_607;
  assign T_614 = T_610 & T_613;
  assign T_619 = T_607 ? 6'h3f : T_606;
  assign GEN_51 = {{63'd0}, T_132};
  assign T_621 = GEN_51 << T_619;
  assign GEN_14 = T_614 ? {{2'd0}, T_621} : T_223;
  assign GEN_15 = T_614 ? {{1'd0}, T_619} : T_200;
  assign T_626 = T_609 & T_221;
  assign T_629 = T_626 & T_175;
  assign GEN_16 = T_629 ? 1'h0 : neg_out;
  assign GEN_17 = T_208 ? GEN_13 : GEN_12;
  assign GEN_18 = T_208 ? GEN_15 : GEN_11;
  assign GEN_19 = T_208 ? {{1'd0}, GEN_14} : GEN_10;
  assign GEN_20 = T_208 ? GEN_16 : neg_out;
  assign T_631 = io_resp_ready & io_resp_valid;
  assign T_632 = T_631 | io_kill;
  assign GEN_21 = T_632 ? 3'h0 : GEN_17;
  assign T_633 = io_req_ready & io_req_valid;
  assign T_635 = T_71 == 1'h0;
  assign T_636 = rhs_sign & T_635;
  assign T_637 = lhs_sign | T_636;
  assign T_638 = T_637 ? 3'h1 : 3'h2;
  assign T_642 = lhs_sign != rhs_sign;
  assign T_643 = T_83 ? lhs_sign : T_642;
  assign T_644 = T_635 & T_643;
  assign T_645 = {rhs_sign,rhs_in};
  assign GEN_22 = T_633 ? T_638 : GEN_21;
  assign GEN_23 = T_633 ? T_71 : isMul;
  assign GEN_24 = T_633 ? T_83 : isHi;
  assign GEN_25 = T_633 ? {{6'd0}, 1'h0} : GEN_18;
  assign GEN_26 = T_633 ? T_644 : GEN_20;
  assign GEN_27 = T_633 ? T_645 : GEN_3;
  assign GEN_28 = T_633 ? {{66'd0}, lhs_in} : GEN_19;
  assign GEN_29 = T_633 ? io_req_bits_fn : req_fn;
  assign GEN_30 = T_633 ? io_req_bits_dw : req_dw;
  assign GEN_31 = T_633 ? io_req_bits_in1 : req_in1;
  assign GEN_32 = T_633 ? io_req_bits_in2 : req_in2;
  assign GEN_33 = T_633 ? io_req_bits_tag : req_tag;
  assign T_650 = 1'h0 == req_dw;
  assign T_652 = remainder[31];
  assign GEN_53 = {{31'd0}, T_652};
  assign T_654 = 32'h0 - GEN_53;
  assign T_655 = T_654[31:0];
  assign T_656 = remainder[31:0];
  assign T_657 = {T_655,T_656};
  assign T_659 = T_650 ? T_657 : T_132;
  assign T_660 = state == 3'h5;
  assign T_661 = state == 3'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_43 = {1{$random}};
  state = GEN_43[2:0];
  GEN_44 = {1{$random}};
  req_fn = GEN_44[3:0];
  GEN_47 = {1{$random}};
  req_dw = GEN_47[0:0];
  GEN_48 = {2{$random}};
  req_in1 = GEN_48[63:0];
  GEN_49 = {2{$random}};
  req_in2 = GEN_49[63:0];
  GEN_52 = {1{$random}};
  req_tag = GEN_52[4:0];
  GEN_54 = {1{$random}};
  count = GEN_54[6:0];
  GEN_55 = {1{$random}};
  neg_out = GEN_55[0:0];
  GEN_56 = {1{$random}};
  isMul = GEN_56[0:0];
  GEN_57 = {1{$random}};
  isHi = GEN_57[0:0];
  GEN_58 = {3{$random}};
  divisor = GEN_58[64:0];
  GEN_59 = {5{$random}};
  remainder = GEN_59[129:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      req_fn <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      req_dw <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      req_in1 <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      req_in2 <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      req_tag <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      count <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      neg_out <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      isMul <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      isHi <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      divisor <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      remainder <= GEN_28;
    end
  end
endmodule
module Rocket(
  input   clk,
  input   reset,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_msip,
  output  io_imem_req_valid,
  output [39:0] io_imem_req_bits_pc,
  output  io_imem_resp_ready,
  input   io_imem_resp_valid,
  input  [39:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_data_0,
  input   io_imem_resp_bits_mask,
  input   io_imem_resp_bits_xcpt_if,
  input   io_imem_btb_resp_valid,
  input   io_imem_btb_resp_bits_taken,
  input   io_imem_btb_resp_bits_mask,
  input   io_imem_btb_resp_bits_bridx,
  input  [38:0] io_imem_btb_resp_bits_target,
  input  [5:0] io_imem_btb_resp_bits_entry,
  input  [6:0] io_imem_btb_resp_bits_bht_history,
  input  [1:0] io_imem_btb_resp_bits_bht_value,
  output  io_imem_btb_update_valid,
  output  io_imem_btb_update_bits_prediction_valid,
  output  io_imem_btb_update_bits_prediction_bits_taken,
  output  io_imem_btb_update_bits_prediction_bits_mask,
  output  io_imem_btb_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_btb_update_bits_prediction_bits_target,
  output [5:0] io_imem_btb_update_bits_prediction_bits_entry,
  output [6:0] io_imem_btb_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_btb_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_btb_update_bits_pc,
  output [38:0] io_imem_btb_update_bits_target,
  output  io_imem_btb_update_bits_taken,
  output  io_imem_btb_update_bits_isJump,
  output  io_imem_btb_update_bits_isReturn,
  output [38:0] io_imem_btb_update_bits_br_pc,
  output  io_imem_bht_update_valid,
  output  io_imem_bht_update_bits_prediction_valid,
  output  io_imem_bht_update_bits_prediction_bits_taken,
  output  io_imem_bht_update_bits_prediction_bits_mask,
  output  io_imem_bht_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_bht_update_bits_prediction_bits_target,
  output [5:0] io_imem_bht_update_bits_prediction_bits_entry,
  output [6:0] io_imem_bht_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_bht_update_bits_prediction_bits_bht_value,
  output [38:0] io_imem_bht_update_bits_pc,
  output  io_imem_bht_update_bits_taken,
  output  io_imem_bht_update_bits_mispredict,
  output  io_imem_ras_update_valid,
  output  io_imem_ras_update_bits_isCall,
  output  io_imem_ras_update_bits_isReturn,
  output [38:0] io_imem_ras_update_bits_returnAddr,
  output  io_imem_ras_update_bits_prediction_valid,
  output  io_imem_ras_update_bits_prediction_bits_taken,
  output  io_imem_ras_update_bits_prediction_bits_mask,
  output  io_imem_ras_update_bits_prediction_bits_bridx,
  output [38:0] io_imem_ras_update_bits_prediction_bits_target,
  output [5:0] io_imem_ras_update_bits_prediction_bits_entry,
  output [6:0] io_imem_ras_update_bits_prediction_bits_bht_history,
  output [1:0] io_imem_ras_update_bits_prediction_bits_bht_value,
  output  io_imem_flush_icache,
  output  io_imem_flush_tlb,
  input  [39:0] io_imem_npc,
  input   io_dmem_req_ready,
  output  io_dmem_req_valid,
  output [39:0] io_dmem_req_bits_addr,
  output [8:0] io_dmem_req_bits_tag,
  output [4:0] io_dmem_req_bits_cmd,
  output [2:0] io_dmem_req_bits_typ,
  output  io_dmem_req_bits_phys,
  output [63:0] io_dmem_req_bits_data,
  output  io_dmem_s1_kill,
  output [63:0] io_dmem_s1_data,
  input   io_dmem_s2_nack,
  input   io_dmem_resp_valid,
  input  [39:0] io_dmem_resp_bits_addr,
  input  [8:0] io_dmem_resp_bits_tag,
  input  [4:0] io_dmem_resp_bits_cmd,
  input  [2:0] io_dmem_resp_bits_typ,
  input  [63:0] io_dmem_resp_bits_data,
  input   io_dmem_resp_bits_replay,
  input   io_dmem_resp_bits_has_data,
  input  [63:0] io_dmem_resp_bits_data_word_bypass,
  input  [63:0] io_dmem_resp_bits_store_data,
  input   io_dmem_replay_next,
  input   io_dmem_xcpt_ma_ld,
  input   io_dmem_xcpt_ma_st,
  input   io_dmem_xcpt_pf_ld,
  input   io_dmem_xcpt_pf_st,
  output  io_dmem_invalidate_lr,
  input   io_dmem_ordered,
  output [19:0] io_ptw_ptbr,
  output  io_ptw_invalidate,
  output  io_ptw_status_debug,
  output [1:0] io_ptw_status_prv,
  output  io_ptw_status_sd,
  output [30:0] io_ptw_status_zero3,
  output  io_ptw_status_sd_rv32,
  output [1:0] io_ptw_status_zero2,
  output [4:0] io_ptw_status_vm,
  output [4:0] io_ptw_status_zero1,
  output  io_ptw_status_pum,
  output  io_ptw_status_mprv,
  output [1:0] io_ptw_status_xs,
  output [1:0] io_ptw_status_fs,
  output [1:0] io_ptw_status_mpp,
  output [1:0] io_ptw_status_hpp,
  output  io_ptw_status_spp,
  output  io_ptw_status_mpie,
  output  io_ptw_status_hpie,
  output  io_ptw_status_spie,
  output  io_ptw_status_upie,
  output  io_ptw_status_mie,
  output  io_ptw_status_hie,
  output  io_ptw_status_sie,
  output  io_ptw_status_uie,
  output [31:0] io_fpu_inst,
  output [63:0] io_fpu_fromint_data,
  output [2:0] io_fpu_fcsr_rm,
  input   io_fpu_fcsr_flags_valid,
  input  [4:0] io_fpu_fcsr_flags_bits,
  input  [63:0] io_fpu_store_data,
  input  [63:0] io_fpu_toint_data,
  output  io_fpu_dmem_resp_val,
  output [2:0] io_fpu_dmem_resp_type,
  output [4:0] io_fpu_dmem_resp_tag,
  output [63:0] io_fpu_dmem_resp_data,
  output  io_fpu_valid,
  input   io_fpu_fcsr_rdy,
  input   io_fpu_nack_mem,
  input   io_fpu_illegal_rm,
  output  io_fpu_killx,
  output  io_fpu_killm,
  input  [4:0] io_fpu_dec_cmd,
  input   io_fpu_dec_ldst,
  input   io_fpu_dec_wen,
  input   io_fpu_dec_ren1,
  input   io_fpu_dec_ren2,
  input   io_fpu_dec_ren3,
  input   io_fpu_dec_swap12,
  input   io_fpu_dec_swap23,
  input   io_fpu_dec_single,
  input   io_fpu_dec_fromint,
  input   io_fpu_dec_toint,
  input   io_fpu_dec_fastpipe,
  input   io_fpu_dec_fma,
  input   io_fpu_dec_div,
  input   io_fpu_dec_sqrt,
  input   io_fpu_dec_round,
  input   io_fpu_dec_wflags,
  input   io_fpu_sboard_set,
  input   io_fpu_sboard_clr,
  input  [4:0] io_fpu_sboard_clra,
  input   io_fpu_cp_req_ready,
  output  io_fpu_cp_req_valid,
  output [4:0] io_fpu_cp_req_bits_cmd,
  output  io_fpu_cp_req_bits_ldst,
  output  io_fpu_cp_req_bits_wen,
  output  io_fpu_cp_req_bits_ren1,
  output  io_fpu_cp_req_bits_ren2,
  output  io_fpu_cp_req_bits_ren3,
  output  io_fpu_cp_req_bits_swap12,
  output  io_fpu_cp_req_bits_swap23,
  output  io_fpu_cp_req_bits_single,
  output  io_fpu_cp_req_bits_fromint,
  output  io_fpu_cp_req_bits_toint,
  output  io_fpu_cp_req_bits_fastpipe,
  output  io_fpu_cp_req_bits_fma,
  output  io_fpu_cp_req_bits_div,
  output  io_fpu_cp_req_bits_sqrt,
  output  io_fpu_cp_req_bits_round,
  output  io_fpu_cp_req_bits_wflags,
  output [2:0] io_fpu_cp_req_bits_rm,
  output [1:0] io_fpu_cp_req_bits_typ,
  output [64:0] io_fpu_cp_req_bits_in1,
  output [64:0] io_fpu_cp_req_bits_in2,
  output [64:0] io_fpu_cp_req_bits_in3,
  output  io_fpu_cp_resp_ready,
  input   io_fpu_cp_resp_valid,
  input  [64:0] io_fpu_cp_resp_bits_data,
  input  [4:0] io_fpu_cp_resp_bits_exc,
  input   io_rocc_cmd_ready,
  output  io_rocc_cmd_valid,
  output [6:0] io_rocc_cmd_bits_inst_funct,
  output [4:0] io_rocc_cmd_bits_inst_rs2,
  output [4:0] io_rocc_cmd_bits_inst_rs1,
  output  io_rocc_cmd_bits_inst_xd,
  output  io_rocc_cmd_bits_inst_xs1,
  output  io_rocc_cmd_bits_inst_xs2,
  output [4:0] io_rocc_cmd_bits_inst_rd,
  output [6:0] io_rocc_cmd_bits_inst_opcode,
  output [63:0] io_rocc_cmd_bits_rs1,
  output [63:0] io_rocc_cmd_bits_rs2,
  output  io_rocc_resp_ready,
  input   io_rocc_resp_valid,
  input  [4:0] io_rocc_resp_bits_rd,
  input  [63:0] io_rocc_resp_bits_data,
  output  io_rocc_mem_req_ready,
  input   io_rocc_mem_req_valid,
  input  [39:0] io_rocc_mem_req_bits_addr,
  input  [8:0] io_rocc_mem_req_bits_tag,
  input  [4:0] io_rocc_mem_req_bits_cmd,
  input  [2:0] io_rocc_mem_req_bits_typ,
  input   io_rocc_mem_req_bits_phys,
  input  [63:0] io_rocc_mem_req_bits_data,
  input   io_rocc_mem_s1_kill,
  input  [63:0] io_rocc_mem_s1_data,
  output  io_rocc_mem_s2_nack,
  output  io_rocc_mem_resp_valid,
  output [39:0] io_rocc_mem_resp_bits_addr,
  output [8:0] io_rocc_mem_resp_bits_tag,
  output [4:0] io_rocc_mem_resp_bits_cmd,
  output [2:0] io_rocc_mem_resp_bits_typ,
  output [63:0] io_rocc_mem_resp_bits_data,
  output  io_rocc_mem_resp_bits_replay,
  output  io_rocc_mem_resp_bits_has_data,
  output [63:0] io_rocc_mem_resp_bits_data_word_bypass,
  output [63:0] io_rocc_mem_resp_bits_store_data,
  output  io_rocc_mem_replay_next,
  output  io_rocc_mem_xcpt_ma_ld,
  output  io_rocc_mem_xcpt_ma_st,
  output  io_rocc_mem_xcpt_pf_ld,
  output  io_rocc_mem_xcpt_pf_st,
  input   io_rocc_mem_invalidate_lr,
  output  io_rocc_mem_ordered,
  input   io_rocc_busy,
  output  io_rocc_status_debug,
  output [1:0] io_rocc_status_prv,
  output  io_rocc_status_sd,
  output [30:0] io_rocc_status_zero3,
  output  io_rocc_status_sd_rv32,
  output [1:0] io_rocc_status_zero2,
  output [4:0] io_rocc_status_vm,
  output [4:0] io_rocc_status_zero1,
  output  io_rocc_status_pum,
  output  io_rocc_status_mprv,
  output [1:0] io_rocc_status_xs,
  output [1:0] io_rocc_status_fs,
  output [1:0] io_rocc_status_mpp,
  output [1:0] io_rocc_status_hpp,
  output  io_rocc_status_spp,
  output  io_rocc_status_mpie,
  output  io_rocc_status_hpie,
  output  io_rocc_status_spie,
  output  io_rocc_status_upie,
  output  io_rocc_status_mie,
  output  io_rocc_status_hie,
  output  io_rocc_status_sie,
  output  io_rocc_status_uie,
  input   io_rocc_interrupt,
  output  io_rocc_autl_acquire_ready,
  input   io_rocc_autl_acquire_valid,
  input  [25:0] io_rocc_autl_acquire_bits_addr_block,
  input  [1:0] io_rocc_autl_acquire_bits_client_xact_id,
  input  [2:0] io_rocc_autl_acquire_bits_addr_beat,
  input   io_rocc_autl_acquire_bits_is_builtin_type,
  input  [2:0] io_rocc_autl_acquire_bits_a_type,
  input  [11:0] io_rocc_autl_acquire_bits_union,
  input  [63:0] io_rocc_autl_acquire_bits_data,
  input   io_rocc_autl_grant_ready,
  output  io_rocc_autl_grant_valid,
  output [2:0] io_rocc_autl_grant_bits_addr_beat,
  output [1:0] io_rocc_autl_grant_bits_client_xact_id,
  output [2:0] io_rocc_autl_grant_bits_manager_xact_id,
  output  io_rocc_autl_grant_bits_is_builtin_type,
  output [3:0] io_rocc_autl_grant_bits_g_type,
  output [63:0] io_rocc_autl_grant_bits_data,
  output  io_rocc_fpu_req_ready,
  input   io_rocc_fpu_req_valid,
  input  [4:0] io_rocc_fpu_req_bits_cmd,
  input   io_rocc_fpu_req_bits_ldst,
  input   io_rocc_fpu_req_bits_wen,
  input   io_rocc_fpu_req_bits_ren1,
  input   io_rocc_fpu_req_bits_ren2,
  input   io_rocc_fpu_req_bits_ren3,
  input   io_rocc_fpu_req_bits_swap12,
  input   io_rocc_fpu_req_bits_swap23,
  input   io_rocc_fpu_req_bits_single,
  input   io_rocc_fpu_req_bits_fromint,
  input   io_rocc_fpu_req_bits_toint,
  input   io_rocc_fpu_req_bits_fastpipe,
  input   io_rocc_fpu_req_bits_fma,
  input   io_rocc_fpu_req_bits_div,
  input   io_rocc_fpu_req_bits_sqrt,
  input   io_rocc_fpu_req_bits_round,
  input   io_rocc_fpu_req_bits_wflags,
  input  [2:0] io_rocc_fpu_req_bits_rm,
  input  [1:0] io_rocc_fpu_req_bits_typ,
  input  [64:0] io_rocc_fpu_req_bits_in1,
  input  [64:0] io_rocc_fpu_req_bits_in2,
  input  [64:0] io_rocc_fpu_req_bits_in3,
  input   io_rocc_fpu_resp_ready,
  output  io_rocc_fpu_resp_valid,
  output [64:0] io_rocc_fpu_resp_bits_data,
  output [4:0] io_rocc_fpu_resp_bits_exc,
  output  io_rocc_exception,
  output [11:0] io_rocc_csr_waddr,
  output [63:0] io_rocc_csr_wdata,
  output  io_rocc_csr_wen,
  output  io_rocc_host_id
);
  reg  ex_ctrl_legal;
  reg [31:0] GEN_295;
  reg  ex_ctrl_fp;
  reg [31:0] GEN_296;
  reg  ex_ctrl_rocc;
  reg [31:0] GEN_297;
  reg  ex_ctrl_branch;
  reg [31:0] GEN_298;
  reg  ex_ctrl_jal;
  reg [31:0] GEN_299;
  reg  ex_ctrl_jalr;
  reg [31:0] GEN_300;
  reg  ex_ctrl_rxs2;
  reg [31:0] GEN_301;
  reg  ex_ctrl_rxs1;
  reg [31:0] GEN_302;
  reg [1:0] ex_ctrl_sel_alu2;
  reg [31:0] GEN_303;
  reg [1:0] ex_ctrl_sel_alu1;
  reg [31:0] GEN_304;
  reg [2:0] ex_ctrl_sel_imm;
  reg [31:0] GEN_305;
  reg  ex_ctrl_alu_dw;
  reg [31:0] GEN_306;
  reg [3:0] ex_ctrl_alu_fn;
  reg [31:0] GEN_307;
  reg  ex_ctrl_mem;
  reg [31:0] GEN_308;
  reg [4:0] ex_ctrl_mem_cmd;
  reg [31:0] GEN_309;
  reg [2:0] ex_ctrl_mem_type;
  reg [31:0] GEN_310;
  reg  ex_ctrl_rfs1;
  reg [31:0] GEN_311;
  reg  ex_ctrl_rfs2;
  reg [31:0] GEN_312;
  reg  ex_ctrl_rfs3;
  reg [31:0] GEN_313;
  reg  ex_ctrl_wfd;
  reg [31:0] GEN_314;
  reg  ex_ctrl_div;
  reg [31:0] GEN_315;
  reg  ex_ctrl_wxd;
  reg [31:0] GEN_316;
  reg [2:0] ex_ctrl_csr;
  reg [31:0] GEN_317;
  reg  ex_ctrl_fence_i;
  reg [31:0] GEN_318;
  reg  ex_ctrl_fence;
  reg [31:0] GEN_319;
  reg  ex_ctrl_amo;
  reg [31:0] GEN_320;
  reg  mem_ctrl_legal;
  reg [31:0] GEN_321;
  reg  mem_ctrl_fp;
  reg [31:0] GEN_322;
  reg  mem_ctrl_rocc;
  reg [31:0] GEN_323;
  reg  mem_ctrl_branch;
  reg [31:0] GEN_324;
  reg  mem_ctrl_jal;
  reg [31:0] GEN_325;
  reg  mem_ctrl_jalr;
  reg [31:0] GEN_326;
  reg  mem_ctrl_rxs2;
  reg [31:0] GEN_327;
  reg  mem_ctrl_rxs1;
  reg [31:0] GEN_328;
  reg [1:0] mem_ctrl_sel_alu2;
  reg [31:0] GEN_329;
  reg [1:0] mem_ctrl_sel_alu1;
  reg [31:0] GEN_330;
  reg [2:0] mem_ctrl_sel_imm;
  reg [31:0] GEN_331;
  reg  mem_ctrl_alu_dw;
  reg [31:0] GEN_332;
  reg [3:0] mem_ctrl_alu_fn;
  reg [31:0] GEN_333;
  reg  mem_ctrl_mem;
  reg [31:0] GEN_334;
  reg [4:0] mem_ctrl_mem_cmd;
  reg [31:0] GEN_335;
  reg [2:0] mem_ctrl_mem_type;
  reg [31:0] GEN_336;
  reg  mem_ctrl_rfs1;
  reg [31:0] GEN_337;
  reg  mem_ctrl_rfs2;
  reg [31:0] GEN_338;
  reg  mem_ctrl_rfs3;
  reg [31:0] GEN_339;
  reg  mem_ctrl_wfd;
  reg [31:0] GEN_340;
  reg  mem_ctrl_div;
  reg [31:0] GEN_341;
  reg  mem_ctrl_wxd;
  reg [31:0] GEN_342;
  reg [2:0] mem_ctrl_csr;
  reg [31:0] GEN_343;
  reg  mem_ctrl_fence_i;
  reg [31:0] GEN_344;
  reg  mem_ctrl_fence;
  reg [31:0] GEN_345;
  reg  mem_ctrl_amo;
  reg [31:0] GEN_346;
  reg  wb_ctrl_legal;
  reg [31:0] GEN_347;
  reg  wb_ctrl_fp;
  reg [31:0] GEN_348;
  reg  wb_ctrl_rocc;
  reg [31:0] GEN_349;
  reg  wb_ctrl_branch;
  reg [31:0] GEN_350;
  reg  wb_ctrl_jal;
  reg [31:0] GEN_351;
  reg  wb_ctrl_jalr;
  reg [31:0] GEN_352;
  reg  wb_ctrl_rxs2;
  reg [31:0] GEN_353;
  reg  wb_ctrl_rxs1;
  reg [31:0] GEN_354;
  reg [1:0] wb_ctrl_sel_alu2;
  reg [31:0] GEN_355;
  reg [1:0] wb_ctrl_sel_alu1;
  reg [31:0] GEN_356;
  reg [2:0] wb_ctrl_sel_imm;
  reg [31:0] GEN_357;
  reg  wb_ctrl_alu_dw;
  reg [31:0] GEN_358;
  reg [3:0] wb_ctrl_alu_fn;
  reg [31:0] GEN_359;
  reg  wb_ctrl_mem;
  reg [31:0] GEN_360;
  reg [4:0] wb_ctrl_mem_cmd;
  reg [31:0] GEN_361;
  reg [2:0] wb_ctrl_mem_type;
  reg [31:0] GEN_362;
  reg  wb_ctrl_rfs1;
  reg [31:0] GEN_363;
  reg  wb_ctrl_rfs2;
  reg [31:0] GEN_364;
  reg  wb_ctrl_rfs3;
  reg [31:0] GEN_365;
  reg  wb_ctrl_wfd;
  reg [31:0] GEN_366;
  reg  wb_ctrl_div;
  reg [31:0] GEN_367;
  reg  wb_ctrl_wxd;
  reg [31:0] GEN_368;
  reg [2:0] wb_ctrl_csr;
  reg [31:0] GEN_369;
  reg  wb_ctrl_fence_i;
  reg [31:0] GEN_370;
  reg  wb_ctrl_fence;
  reg [31:0] GEN_371;
  reg  wb_ctrl_amo;
  reg [31:0] GEN_372;
  reg  ex_reg_xcpt_interrupt;
  reg [31:0] GEN_373;
  reg  ex_reg_valid;
  reg [31:0] GEN_374;
  reg  ex_reg_btb_hit;
  reg [31:0] GEN_375;
  reg  ex_reg_btb_resp_taken;
  reg [31:0] GEN_376;
  reg  ex_reg_btb_resp_mask;
  reg [31:0] GEN_377;
  reg  ex_reg_btb_resp_bridx;
  reg [31:0] GEN_378;
  reg [38:0] ex_reg_btb_resp_target;
  reg [63:0] GEN_379;
  reg [5:0] ex_reg_btb_resp_entry;
  reg [31:0] GEN_380;
  reg [6:0] ex_reg_btb_resp_bht_history;
  reg [31:0] GEN_381;
  reg [1:0] ex_reg_btb_resp_bht_value;
  reg [31:0] GEN_382;
  reg  ex_reg_xcpt;
  reg [31:0] GEN_383;
  reg  ex_reg_flush_pipe;
  reg [31:0] GEN_384;
  reg  ex_reg_load_use;
  reg [31:0] GEN_385;
  reg [63:0] ex_reg_cause;
  reg [63:0] GEN_386;
  reg [39:0] ex_reg_pc;
  reg [63:0] GEN_387;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_388;
  reg  mem_reg_xcpt_interrupt;
  reg [31:0] GEN_389;
  reg  mem_reg_valid;
  reg [31:0] GEN_390;
  reg  mem_reg_btb_hit;
  reg [31:0] GEN_391;
  reg  mem_reg_btb_resp_taken;
  reg [31:0] GEN_392;
  reg  mem_reg_btb_resp_mask;
  reg [31:0] GEN_393;
  reg  mem_reg_btb_resp_bridx;
  reg [31:0] GEN_394;
  reg [38:0] mem_reg_btb_resp_target;
  reg [63:0] GEN_395;
  reg [5:0] mem_reg_btb_resp_entry;
  reg [31:0] GEN_396;
  reg [6:0] mem_reg_btb_resp_bht_history;
  reg [31:0] GEN_397;
  reg [1:0] mem_reg_btb_resp_bht_value;
  reg [31:0] GEN_398;
  reg  mem_reg_xcpt;
  reg [31:0] GEN_399;
  reg  mem_reg_replay;
  reg [31:0] GEN_400;
  reg  mem_reg_flush_pipe;
  reg [31:0] GEN_401;
  reg [63:0] mem_reg_cause;
  reg [63:0] GEN_402;
  reg  mem_reg_slow_bypass;
  reg [31:0] GEN_403;
  reg  mem_reg_load;
  reg [31:0] GEN_404;
  reg  mem_reg_store;
  reg [31:0] GEN_405;
  reg [39:0] mem_reg_pc;
  reg [63:0] GEN_406;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_407;
  reg [63:0] mem_reg_wdata;
  reg [63:0] GEN_408;
  reg [63:0] mem_reg_rs2;
  reg [63:0] GEN_409;
  wire  take_pc_mem;
  reg  wb_reg_valid;
  reg [31:0] GEN_410;
  reg  wb_reg_xcpt;
  reg [31:0] GEN_411;
  reg  wb_reg_mem_xcpt;
  reg [31:0] GEN_412;
  reg  wb_reg_replay;
  reg [31:0] GEN_413;
  reg [63:0] wb_reg_cause;
  reg [63:0] GEN_414;
  reg  wb_reg_rocc_pending;
  reg [31:0] GEN_415;
  reg [39:0] wb_reg_pc;
  reg [63:0] GEN_416;
  reg [31:0] wb_reg_inst;
  reg [31:0] GEN_417;
  reg [63:0] wb_reg_wdata;
  reg [63:0] GEN_418;
  reg [63:0] wb_reg_rs2;
  reg [63:0] GEN_419;
  wire  take_pc_wb;
  wire  take_pc_mem_wb;
  wire  id_ctrl_legal;
  wire  id_ctrl_fp;
  wire  id_ctrl_rocc;
  wire  id_ctrl_branch;
  wire  id_ctrl_jal;
  wire  id_ctrl_jalr;
  wire  id_ctrl_rxs2;
  wire  id_ctrl_rxs1;
  wire [1:0] id_ctrl_sel_alu2;
  wire [1:0] id_ctrl_sel_alu1;
  wire [2:0] id_ctrl_sel_imm;
  wire  id_ctrl_alu_dw;
  wire [3:0] id_ctrl_alu_fn;
  wire  id_ctrl_mem;
  wire [4:0] id_ctrl_mem_cmd;
  wire [2:0] id_ctrl_mem_type;
  wire  id_ctrl_rfs1;
  wire  id_ctrl_rfs2;
  wire  id_ctrl_rfs3;
  wire  id_ctrl_wfd;
  wire  id_ctrl_div;
  wire  id_ctrl_wxd;
  wire [2:0] id_ctrl_csr;
  wire  id_ctrl_fence_i;
  wire  id_ctrl_fence;
  wire  id_ctrl_amo;
  wire [31:0] T_6584;
  wire  T_6586;
  wire [31:0] T_6588;
  wire  T_6590;
  wire [31:0] T_6592;
  wire  T_6594;
  wire [31:0] T_6596;
  wire  T_6598;
  wire [31:0] T_6600;
  wire  T_6602;
  wire [31:0] T_6604;
  wire  T_6606;
  wire [31:0] T_6608;
  wire  T_6610;
  wire [31:0] T_6612;
  wire  T_6614;
  wire [31:0] T_6616;
  wire  T_6618;
  wire [31:0] T_6620;
  wire  T_6622;
  wire [31:0] T_6624;
  wire  T_6626;
  wire [31:0] T_6628;
  wire  T_6630;
  wire [31:0] T_6632;
  wire  T_6634;
  wire [31:0] T_6636;
  wire  T_6638;
  wire [31:0] T_6640;
  wire  T_6642;
  wire  T_6646;
  wire [31:0] T_6648;
  wire  T_6650;
  wire  T_6654;
  wire [31:0] T_6656;
  wire  T_6658;
  wire [31:0] T_6660;
  wire  T_6662;
  wire  T_6666;
  wire [31:0] T_6668;
  wire  T_6670;
  wire [31:0] T_6672;
  wire  T_6674;
  wire [31:0] T_6676;
  wire  T_6678;
  wire [31:0] T_6680;
  wire  T_6682;
  wire [31:0] T_6684;
  wire  T_6686;
  wire  T_6688;
  wire [31:0] T_6690;
  wire  T_6692;
  wire [31:0] T_6694;
  wire  T_6696;
  wire [31:0] T_6698;
  wire  T_6700;
  wire [31:0] T_6702;
  wire  T_6704;
  wire  T_6708;
  wire [31:0] T_6710;
  wire  T_6712;
  wire  T_6714;
  wire [31:0] T_6716;
  wire  T_6718;
  wire [31:0] T_6720;
  wire  T_6722;
  wire [31:0] T_6724;
  wire  T_6726;
  wire [31:0] T_6728;
  wire  T_6730;
  wire [31:0] T_6732;
  wire  T_6734;
  wire [31:0] T_6736;
  wire  T_6738;
  wire [31:0] T_6740;
  wire  T_6742;
  wire  T_6745;
  wire  T_6746;
  wire  T_6747;
  wire  T_6748;
  wire  T_6749;
  wire  T_6750;
  wire  T_6751;
  wire  T_6752;
  wire  T_6753;
  wire  T_6754;
  wire  T_6755;
  wire  T_6756;
  wire  T_6757;
  wire  T_6758;
  wire  T_6759;
  wire  T_6760;
  wire  T_6761;
  wire  T_6762;
  wire  T_6763;
  wire  T_6764;
  wire  T_6765;
  wire  T_6766;
  wire  T_6767;
  wire  T_6768;
  wire  T_6769;
  wire  T_6770;
  wire  T_6771;
  wire  T_6772;
  wire  T_6773;
  wire  T_6774;
  wire  T_6775;
  wire  T_6776;
  wire  T_6777;
  wire  T_6778;
  wire  T_6779;
  wire  T_6780;
  wire  T_6781;
  wire  T_6782;
  wire  T_6783;
  wire  T_6784;
  wire [31:0] T_6786;
  wire  T_6788;
  wire [31:0] T_6790;
  wire  T_6792;
  wire  T_6795;
  wire [31:0] T_6798;
  wire  T_6800;
  wire [31:0] T_6804;
  wire  T_6806;
  wire [31:0] T_6810;
  wire  T_6812;
  wire [31:0] T_6816;
  wire  T_6818;
  wire [31:0] T_6820;
  wire  T_6822;
  wire [31:0] T_6824;
  wire  T_6826;
  wire  T_6829;
  wire  T_6830;
  wire [31:0] T_6832;
  wire  T_6834;
  wire [31:0] T_6836;
  wire  T_6838;
  wire [31:0] T_6840;
  wire  T_6842;
  wire [31:0] T_6844;
  wire  T_6846;
  wire [31:0] T_6848;
  wire  T_6850;
  wire  T_6853;
  wire  T_6854;
  wire  T_6855;
  wire  T_6856;
  wire [31:0] T_6858;
  wire  T_6860;
  wire [31:0] T_6862;
  wire  T_6864;
  wire [31:0] T_6866;
  wire  T_6868;
  wire [31:0] T_6870;
  wire  T_6872;
  wire [31:0] T_6874;
  wire  T_6876;
  wire  T_6879;
  wire  T_6880;
  wire  T_6881;
  wire  T_6882;
  wire  T_6886;
  wire [31:0] T_6888;
  wire  T_6890;
  wire [31:0] T_6892;
  wire  T_6894;
  wire  T_6897;
  wire  T_6898;
  wire  T_6899;
  wire [1:0] T_6900;
  wire [31:0] T_6902;
  wire  T_6904;
  wire [31:0] T_6906;
  wire  T_6908;
  wire [31:0] T_6910;
  wire  T_6912;
  wire  T_6915;
  wire  T_6916;
  wire  T_6917;
  wire  T_6918;
  wire  T_6922;
  wire  T_6925;
  wire [1:0] T_6926;
  wire  T_6930;
  wire  T_6934;
  wire  T_6937;
  wire [31:0] T_6939;
  wire  T_6941;
  wire  T_6944;
  wire [31:0] T_6946;
  wire  T_6948;
  wire [31:0] T_6950;
  wire  T_6952;
  wire  T_6956;
  wire  T_6959;
  wire  T_6960;
  wire [1:0] T_6961;
  wire [2:0] T_6962;
  wire [31:0] T_6964;
  wire  T_6966;
  wire [31:0] T_6968;
  wire  T_6970;
  wire  T_6973;
  wire [31:0] T_6975;
  wire  T_6977;
  wire [31:0] T_6979;
  wire  T_6981;
  wire [31:0] T_6983;
  wire  T_6985;
  wire  T_6988;
  wire  T_6989;
  wire [31:0] T_6991;
  wire  T_6993;
  wire [31:0] T_6995;
  wire  T_6997;
  wire  T_7001;
  wire [31:0] T_7003;
  wire  T_7005;
  wire [31:0] T_7007;
  wire  T_7009;
  wire [31:0] T_7011;
  wire  T_7013;
  wire  T_7016;
  wire  T_7017;
  wire  T_7018;
  wire  T_7019;
  wire  T_7020;
  wire [31:0] T_7022;
  wire  T_7024;
  wire [31:0] T_7026;
  wire  T_7028;
  wire [31:0] T_7030;
  wire  T_7032;
  wire [31:0] T_7034;
  wire  T_7036;
  wire  T_7039;
  wire  T_7040;
  wire  T_7041;
  wire  T_7045;
  wire [31:0] T_7047;
  wire  T_7049;
  wire  T_7052;
  wire  T_7053;
  wire  T_7054;
  wire [1:0] T_7055;
  wire [2:0] T_7056;
  wire [3:0] T_7057;
  wire [31:0] T_7059;
  wire  T_7061;
  wire [31:0] T_7063;
  wire  T_7065;
  wire [31:0] T_7067;
  wire  T_7069;
  wire  T_7072;
  wire  T_7073;
  wire  T_7074;
  wire  T_7075;
  wire  T_7076;
  wire  T_7077;
  wire  T_7078;
  wire [31:0] T_7080;
  wire  T_7082;
  wire [31:0] T_7084;
  wire  T_7086;
  wire [31:0] T_7088;
  wire  T_7090;
  wire [31:0] T_7092;
  wire  T_7094;
  wire  T_7097;
  wire  T_7098;
  wire  T_7099;
  wire [31:0] T_7101;
  wire  T_7103;
  wire [31:0] T_7105;
  wire  T_7107;
  wire  T_7110;
  wire [31:0] T_7112;
  wire  T_7114;
  wire [31:0] T_7116;
  wire  T_7118;
  wire [31:0] T_7120;
  wire  T_7122;
  wire  T_7125;
  wire  T_7126;
  wire  T_7127;
  wire [31:0] T_7129;
  wire  T_7131;
  wire [1:0] T_7135;
  wire [2:0] T_7136;
  wire [3:0] T_7137;
  wire [4:0] T_7138;
  wire [31:0] T_7140;
  wire  T_7142;
  wire [31:0] T_7146;
  wire  T_7148;
  wire [31:0] T_7152;
  wire  T_7154;
  wire [1:0] T_7157;
  wire [2:0] T_7158;
  wire [31:0] T_7160;
  wire  T_7162;
  wire [31:0] T_7164;
  wire  T_7166;
  wire [31:0] T_7168;
  wire  T_7170;
  wire  T_7173;
  wire  T_7174;
  wire [31:0] T_7176;
  wire  T_7178;
  wire [31:0] T_7180;
  wire  T_7182;
  wire [31:0] T_7184;
  wire  T_7186;
  wire  T_7189;
  wire  T_7190;
  wire  T_7191;
  wire [31:0] T_7195;
  wire  T_7197;
  wire  T_7201;
  wire  T_7204;
  wire  T_7205;
  wire  T_7206;
  wire [31:0] T_7208;
  wire  T_7210;
  wire  T_7216;
  wire  T_7220;
  wire [31:0] T_7222;
  wire  T_7224;
  wire  T_7228;
  wire [31:0] T_7230;
  wire  T_7232;
  wire [31:0] T_7234;
  wire  T_7236;
  wire [31:0] T_7238;
  wire  T_7240;
  wire  T_7243;
  wire  T_7244;
  wire  T_7245;
  wire  T_7246;
  wire  T_7247;
  wire  T_7248;
  wire [31:0] T_7250;
  wire  T_7252;
  wire [31:0] T_7256;
  wire  T_7258;
  wire [31:0] T_7262;
  wire  T_7264;
  wire [1:0] T_7267;
  wire [2:0] T_7268;
  wire [31:0] T_7270;
  wire  T_7272;
  wire  T_7278;
  wire [31:0] T_7282;
  wire  T_7284;
  wire [4:0] id_raddr3;
  wire [4:0] id_raddr2;
  wire [4:0] id_raddr1;
  wire [4:0] id_waddr;
  wire  id_load_use;
  reg  id_reg_fence;
  reg [31:0] GEN_420;
  reg [63:0] T_7291 [0:30];
  reg [63:0] GEN_421;
  wire [63:0] T_7291_T_7301_data;
  wire [4:0] T_7291_T_7301_addr;
  wire  T_7291_T_7301_en;
  wire [63:0] T_7291_T_7312_data;
  wire [4:0] T_7291_T_7312_addr;
  wire  T_7291_T_7312_en;
  wire [63:0] T_7291_T_7961_data;
  wire [4:0] T_7291_T_7961_addr;
  wire  T_7291_T_7961_mask;
  wire  T_7291_T_7961_en;
  wire [63:0] T_7293;
  wire [4:0] GEN_173;
  wire  T_7296;
  wire [4:0] T_7300;
  wire [63:0] T_7302;
  wire [63:0] T_7304;
  wire [4:0] T_7311;
  wire [63:0] T_7313;
  wire  ctrl_killd;
  wire  csr_clk;
  wire  csr_reset;
  wire  csr_io_prci_reset;
  wire  csr_io_prci_id;
  wire  csr_io_prci_interrupts_mtip;
  wire  csr_io_prci_interrupts_meip;
  wire  csr_io_prci_interrupts_seip;
  wire  csr_io_prci_interrupts_debug;
  wire  csr_io_prci_interrupts_msip;
  wire [11:0] csr_io_rw_addr;
  wire [2:0] csr_io_rw_cmd;
  wire [63:0] csr_io_rw_rdata;
  wire [63:0] csr_io_rw_wdata;
  wire  csr_io_csr_stall;
  wire  csr_io_csr_xcpt;
  wire  csr_io_eret;
  wire [1:0] csr_io_prv;
  wire  csr_io_status_debug;
  wire [1:0] csr_io_status_prv;
  wire  csr_io_status_sd;
  wire [30:0] csr_io_status_zero3;
  wire  csr_io_status_sd_rv32;
  wire [1:0] csr_io_status_zero2;
  wire [4:0] csr_io_status_vm;
  wire [4:0] csr_io_status_zero1;
  wire  csr_io_status_pum;
  wire  csr_io_status_mprv;
  wire [1:0] csr_io_status_xs;
  wire [1:0] csr_io_status_fs;
  wire [1:0] csr_io_status_mpp;
  wire [1:0] csr_io_status_hpp;
  wire  csr_io_status_spp;
  wire  csr_io_status_mpie;
  wire  csr_io_status_hpie;
  wire  csr_io_status_spie;
  wire  csr_io_status_upie;
  wire  csr_io_status_mie;
  wire  csr_io_status_hie;
  wire  csr_io_status_sie;
  wire  csr_io_status_uie;
  wire [31:0] csr_io_ptbr;
  wire [39:0] csr_io_evec;
  wire  csr_io_exception;
  wire  csr_io_retire;
  wire  csr_io_uarch_counters_0;
  wire  csr_io_uarch_counters_1;
  wire  csr_io_uarch_counters_2;
  wire  csr_io_uarch_counters_3;
  wire  csr_io_uarch_counters_4;
  wire  csr_io_uarch_counters_5;
  wire  csr_io_uarch_counters_6;
  wire  csr_io_uarch_counters_7;
  wire  csr_io_uarch_counters_8;
  wire  csr_io_uarch_counters_9;
  wire  csr_io_uarch_counters_10;
  wire  csr_io_uarch_counters_11;
  wire  csr_io_uarch_counters_12;
  wire  csr_io_uarch_counters_13;
  wire  csr_io_uarch_counters_14;
  wire  csr_io_uarch_counters_15;
  wire [63:0] csr_io_cause;
  wire [39:0] csr_io_pc;
  wire [39:0] csr_io_badaddr;
  wire  csr_io_fatc;
  wire [63:0] csr_io_time;
  wire [2:0] csr_io_fcsr_rm;
  wire  csr_io_fcsr_flags_valid;
  wire [4:0] csr_io_fcsr_flags_bits;
  wire  csr_io_rocc_cmd_ready;
  wire  csr_io_rocc_cmd_valid;
  wire [6:0] csr_io_rocc_cmd_bits_inst_funct;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rs1;
  wire  csr_io_rocc_cmd_bits_inst_xd;
  wire  csr_io_rocc_cmd_bits_inst_xs1;
  wire  csr_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] csr_io_rocc_cmd_bits_inst_rd;
  wire [6:0] csr_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] csr_io_rocc_cmd_bits_rs1;
  wire [63:0] csr_io_rocc_cmd_bits_rs2;
  wire  csr_io_rocc_resp_ready;
  wire  csr_io_rocc_resp_valid;
  wire [4:0] csr_io_rocc_resp_bits_rd;
  wire [63:0] csr_io_rocc_resp_bits_data;
  wire  csr_io_rocc_mem_req_ready;
  wire  csr_io_rocc_mem_req_valid;
  wire [39:0] csr_io_rocc_mem_req_bits_addr;
  wire [8:0] csr_io_rocc_mem_req_bits_tag;
  wire [4:0] csr_io_rocc_mem_req_bits_cmd;
  wire [2:0] csr_io_rocc_mem_req_bits_typ;
  wire  csr_io_rocc_mem_req_bits_phys;
  wire [63:0] csr_io_rocc_mem_req_bits_data;
  wire  csr_io_rocc_mem_s1_kill;
  wire [63:0] csr_io_rocc_mem_s1_data;
  wire  csr_io_rocc_mem_s2_nack;
  wire  csr_io_rocc_mem_resp_valid;
  wire [39:0] csr_io_rocc_mem_resp_bits_addr;
  wire [8:0] csr_io_rocc_mem_resp_bits_tag;
  wire [4:0] csr_io_rocc_mem_resp_bits_cmd;
  wire [2:0] csr_io_rocc_mem_resp_bits_typ;
  wire [63:0] csr_io_rocc_mem_resp_bits_data;
  wire  csr_io_rocc_mem_resp_bits_replay;
  wire  csr_io_rocc_mem_resp_bits_has_data;
  wire [63:0] csr_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] csr_io_rocc_mem_resp_bits_store_data;
  wire  csr_io_rocc_mem_replay_next;
  wire  csr_io_rocc_mem_xcpt_ma_ld;
  wire  csr_io_rocc_mem_xcpt_ma_st;
  wire  csr_io_rocc_mem_xcpt_pf_ld;
  wire  csr_io_rocc_mem_xcpt_pf_st;
  wire  csr_io_rocc_mem_invalidate_lr;
  wire  csr_io_rocc_mem_ordered;
  wire  csr_io_rocc_busy;
  wire  csr_io_rocc_status_debug;
  wire [1:0] csr_io_rocc_status_prv;
  wire  csr_io_rocc_status_sd;
  wire [30:0] csr_io_rocc_status_zero3;
  wire  csr_io_rocc_status_sd_rv32;
  wire [1:0] csr_io_rocc_status_zero2;
  wire [4:0] csr_io_rocc_status_vm;
  wire [4:0] csr_io_rocc_status_zero1;
  wire  csr_io_rocc_status_pum;
  wire  csr_io_rocc_status_mprv;
  wire [1:0] csr_io_rocc_status_xs;
  wire [1:0] csr_io_rocc_status_fs;
  wire [1:0] csr_io_rocc_status_mpp;
  wire [1:0] csr_io_rocc_status_hpp;
  wire  csr_io_rocc_status_spp;
  wire  csr_io_rocc_status_mpie;
  wire  csr_io_rocc_status_hpie;
  wire  csr_io_rocc_status_spie;
  wire  csr_io_rocc_status_upie;
  wire  csr_io_rocc_status_mie;
  wire  csr_io_rocc_status_hie;
  wire  csr_io_rocc_status_sie;
  wire  csr_io_rocc_status_uie;
  wire  csr_io_rocc_interrupt;
  wire  csr_io_rocc_autl_acquire_ready;
  wire  csr_io_rocc_autl_acquire_valid;
  wire [25:0] csr_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] csr_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_acquire_bits_addr_beat;
  wire  csr_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] csr_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] csr_io_rocc_autl_acquire_bits_union;
  wire [63:0] csr_io_rocc_autl_acquire_bits_data;
  wire  csr_io_rocc_autl_grant_ready;
  wire  csr_io_rocc_autl_grant_valid;
  wire [2:0] csr_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] csr_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] csr_io_rocc_autl_grant_bits_manager_xact_id;
  wire  csr_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] csr_io_rocc_autl_grant_bits_g_type;
  wire [63:0] csr_io_rocc_autl_grant_bits_data;
  wire  csr_io_rocc_fpu_req_ready;
  wire  csr_io_rocc_fpu_req_valid;
  wire [4:0] csr_io_rocc_fpu_req_bits_cmd;
  wire  csr_io_rocc_fpu_req_bits_ldst;
  wire  csr_io_rocc_fpu_req_bits_wen;
  wire  csr_io_rocc_fpu_req_bits_ren1;
  wire  csr_io_rocc_fpu_req_bits_ren2;
  wire  csr_io_rocc_fpu_req_bits_ren3;
  wire  csr_io_rocc_fpu_req_bits_swap12;
  wire  csr_io_rocc_fpu_req_bits_swap23;
  wire  csr_io_rocc_fpu_req_bits_single;
  wire  csr_io_rocc_fpu_req_bits_fromint;
  wire  csr_io_rocc_fpu_req_bits_toint;
  wire  csr_io_rocc_fpu_req_bits_fastpipe;
  wire  csr_io_rocc_fpu_req_bits_fma;
  wire  csr_io_rocc_fpu_req_bits_div;
  wire  csr_io_rocc_fpu_req_bits_sqrt;
  wire  csr_io_rocc_fpu_req_bits_round;
  wire  csr_io_rocc_fpu_req_bits_wflags;
  wire [2:0] csr_io_rocc_fpu_req_bits_rm;
  wire [1:0] csr_io_rocc_fpu_req_bits_typ;
  wire [64:0] csr_io_rocc_fpu_req_bits_in1;
  wire [64:0] csr_io_rocc_fpu_req_bits_in2;
  wire [64:0] csr_io_rocc_fpu_req_bits_in3;
  wire  csr_io_rocc_fpu_resp_ready;
  wire  csr_io_rocc_fpu_resp_valid;
  wire [64:0] csr_io_rocc_fpu_resp_bits_data;
  wire [4:0] csr_io_rocc_fpu_resp_bits_exc;
  wire  csr_io_rocc_exception;
  wire [11:0] csr_io_rocc_csr_waddr;
  wire [63:0] csr_io_rocc_csr_wdata;
  wire  csr_io_rocc_csr_wen;
  wire  csr_io_rocc_host_id;
  wire  csr_io_interrupt;
  wire [63:0] csr_io_interrupt_cause;
  wire [3:0] csr_io_bp_0_control_tdrtype;
  wire [4:0] csr_io_bp_0_control_bpamaskmax;
  wire [35:0] csr_io_bp_0_control_reserved;
  wire [7:0] csr_io_bp_0_control_bpaction;
  wire [3:0] csr_io_bp_0_control_bpmatch;
  wire  csr_io_bp_0_control_m;
  wire  csr_io_bp_0_control_h;
  wire  csr_io_bp_0_control_s;
  wire  csr_io_bp_0_control_u;
  wire  csr_io_bp_0_control_r;
  wire  csr_io_bp_0_control_w;
  wire  csr_io_bp_0_control_x;
  wire [38:0] csr_io_bp_0_address;
  wire  id_csr_en;
  wire  id_system_insn;
  wire  T_7315;
  wire  T_7316;
  wire  T_7317;
  wire  id_csr_ren;
  wire [2:0] id_csr;
  wire [11:0] id_csr_addr;
  wire  T_7321;
  wire  T_7322;
  wire [11:0] T_7377;
  wire  T_7379;
  wire [11:0] T_7381;
  wire  T_7383;
  wire  T_7386;
  wire  T_7389;
  wire  T_7390;
  wire  id_csr_flush;
  wire  T_7392;
  wire [1:0] GEN_176;
  wire  T_7394;
  wire  T_7396;
  wire  T_7397;
  wire  T_7398;
  wire  T_7400;
  wire  T_7402;
  wire  T_7403;
  wire  id_illegal_insn;
  wire  id_amo_aq;
  wire  id_amo_rl;
  wire  T_7404;
  wire  id_fence_next;
  wire  T_7406;
  wire  id_mem_busy;
  wire  T_7412;
  wire  T_7414;
  wire  T_7415;
  wire  T_7417;
  wire  T_7418;
  wire  T_7419;
  wire  T_7420;
  wire  T_7421;
  wire  T_7422;
  wire  T_7423;
  wire  bpu_clk;
  wire  bpu_reset;
  wire  bpu_io_status_debug;
  wire [1:0] bpu_io_status_prv;
  wire  bpu_io_status_sd;
  wire [30:0] bpu_io_status_zero3;
  wire  bpu_io_status_sd_rv32;
  wire [1:0] bpu_io_status_zero2;
  wire [4:0] bpu_io_status_vm;
  wire [4:0] bpu_io_status_zero1;
  wire  bpu_io_status_pum;
  wire  bpu_io_status_mprv;
  wire [1:0] bpu_io_status_xs;
  wire [1:0] bpu_io_status_fs;
  wire [1:0] bpu_io_status_mpp;
  wire [1:0] bpu_io_status_hpp;
  wire  bpu_io_status_spp;
  wire  bpu_io_status_mpie;
  wire  bpu_io_status_hpie;
  wire  bpu_io_status_spie;
  wire  bpu_io_status_upie;
  wire  bpu_io_status_mie;
  wire  bpu_io_status_hie;
  wire  bpu_io_status_sie;
  wire  bpu_io_status_uie;
  wire [3:0] bpu_io_bp_0_control_tdrtype;
  wire [4:0] bpu_io_bp_0_control_bpamaskmax;
  wire [35:0] bpu_io_bp_0_control_reserved;
  wire [7:0] bpu_io_bp_0_control_bpaction;
  wire [3:0] bpu_io_bp_0_control_bpmatch;
  wire  bpu_io_bp_0_control_m;
  wire  bpu_io_bp_0_control_h;
  wire  bpu_io_bp_0_control_s;
  wire  bpu_io_bp_0_control_u;
  wire  bpu_io_bp_0_control_r;
  wire  bpu_io_bp_0_control_w;
  wire  bpu_io_bp_0_control_x;
  wire [38:0] bpu_io_bp_0_address;
  wire [38:0] bpu_io_pc;
  wire [38:0] bpu_io_ea;
  wire  bpu_io_xcpt_if;
  wire  bpu_io_xcpt_ld;
  wire  bpu_io_xcpt_st;
  wire  T_7427;
  wire  T_7428;
  wire  id_xcpt;
  wire [1:0] T_7429;
  wire [1:0] T_7430;
  wire [63:0] id_cause;
  wire [4:0] ex_waddr;
  wire [4:0] mem_waddr;
  wire [4:0] wb_waddr;
  wire  T_7434;
  wire  T_7435;
  wire  T_7437;
  wire  T_7438;
  wire  T_7440;
  wire  T_7442;
  wire  T_7443;
  wire  T_7444;
  wire  T_7445;
  wire  T_7447;
  wire  T_7448;
  wire  T_7450;
  wire  T_7451;
  wire  T_7452;
  wire  T_7453;
  wire  T_7455;
  wire [63:0] bypass_mux_0;
  wire [63:0] bypass_mux_1;
  wire [63:0] bypass_mux_2;
  wire [63:0] bypass_mux_3;
  reg  ex_reg_rs_bypass_0;
  reg [31:0] GEN_422;
  reg  ex_reg_rs_bypass_1;
  reg [31:0] GEN_423;
  reg [1:0] ex_reg_rs_lsb_0;
  reg [31:0] GEN_424;
  reg [1:0] ex_reg_rs_lsb_1;
  reg [31:0] GEN_425;
  reg [61:0] ex_reg_rs_msb_0;
  reg [63:0] GEN_426;
  reg [61:0] ex_reg_rs_msb_1;
  reg [63:0] GEN_427;
  wire [63:0] T_7483;
  wire [63:0] GEN_0;
  wire [1:0] GEN_180;
  wire [63:0] GEN_2;
  wire [63:0] GEN_3;
  wire [63:0] GEN_4;
  wire [63:0] T_7484;
  wire [63:0] T_7485;
  wire [63:0] GEN_1;
  wire [63:0] GEN_5;
  wire [63:0] GEN_6;
  wire [63:0] GEN_7;
  wire [63:0] T_7486;
  wire  T_7487;
  wire  T_7489;
  wire  T_7490;
  wire  T_7491;
  wire  T_7492;
  wire [10:0] T_7493;
  wire [10:0] T_7494;
  wire [10:0] T_7495;
  wire  T_7496;
  wire  T_7497;
  wire  T_7498;
  wire [7:0] T_7499;
  wire [7:0] T_7500;
  wire [7:0] T_7501;
  wire  T_7504;
  wire  T_7506;
  wire  T_7507;
  wire  T_7508;
  wire  T_7509;
  wire  T_7510;
  wire  T_7511;
  wire  T_7512;
  wire  T_7513;
  wire  T_7514;
  wire [5:0] T_7519;
  wire [5:0] T_7520;
  wire  T_7523;
  wire  T_7525;
  wire [3:0] T_7526;
  wire [3:0] T_7528;
  wire [3:0] T_7529;
  wire [3:0] T_7530;
  wire [3:0] T_7531;
  wire [3:0] T_7532;
  wire  T_7535;
  wire  T_7538;
  wire  T_7541;
  wire  T_7543;
  wire  T_7545;
  wire [9:0] T_7546;
  wire [10:0] T_7547;
  wire  T_7548;
  wire [7:0] T_7549;
  wire [8:0] T_7550;
  wire [10:0] T_7551;
  wire  T_7552;
  wire [11:0] T_7553;
  wire [20:0] T_7554;
  wire [31:0] T_7555;
  wire [31:0] ex_imm;
  wire [63:0] T_7557;
  wire [39:0] T_7558;
  wire  T_7559;
  wire  GEN_182;
  wire [39:0] T_7560;
  wire  T_7561;
  wire [63:0] ex_op1;
  wire [63:0] T_7563;
  wire  T_7565;
  wire [3:0] T_7566;
  wire  T_7567;
  wire [31:0] T_7568;
  wire  T_7569;
  wire [63:0] ex_op2;
  wire  alu_clk;
  wire  alu_reset;
  wire  alu_io_dw;
  wire [3:0] alu_io_fn;
  wire [63:0] alu_io_in2;
  wire [63:0] alu_io_in1;
  wire [63:0] alu_io_out;
  wire [63:0] alu_io_adder_out;
  wire  alu_io_cmp_out;
  wire [63:0] T_7570;
  wire [63:0] T_7571;
  wire  div_clk;
  wire  div_reset;
  wire  div_io_req_ready;
  wire  div_io_req_valid;
  wire [3:0] div_io_req_bits_fn;
  wire  div_io_req_bits_dw;
  wire [63:0] div_io_req_bits_in1;
  wire [63:0] div_io_req_bits_in2;
  wire [4:0] div_io_req_bits_tag;
  wire  div_io_kill;
  wire  div_io_resp_ready;
  wire  div_io_resp_valid;
  wire [63:0] div_io_resp_bits_data;
  wire [4:0] div_io_resp_bits_tag;
  wire  T_7572;
  wire  T_7574;
  wire  T_7577;
  wire  T_7579;
  wire  T_7580;
  wire  T_7581;
  wire [63:0] GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire [38:0] GEN_12;
  wire [5:0] GEN_13;
  wire [6:0] GEN_14;
  wire [1:0] GEN_15;
  wire  T_7584;
  wire  T_7585;
  wire  T_7586;
  wire  T_7587;
  wire [1:0] T_7592;
  wire [1:0] T_7593;
  wire [1:0] T_7594;
  wire  T_7596;
  wire  T_7597;
  wire [1:0] T_7598;
  wire [61:0] T_7599;
  wire [1:0] GEN_16;
  wire [61:0] GEN_17;
  wire  T_7600;
  wire  T_7601;
  wire  T_7602;
  wire [1:0] T_7607;
  wire [1:0] T_7608;
  wire [1:0] T_7609;
  wire  T_7611;
  wire  T_7612;
  wire [1:0] T_7613;
  wire [61:0] T_7614;
  wire [1:0] GEN_18;
  wire [61:0] GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire [1:0] GEN_28;
  wire [1:0] GEN_29;
  wire [2:0] GEN_30;
  wire  GEN_31;
  wire [3:0] GEN_32;
  wire  GEN_33;
  wire [4:0] GEN_34;
  wire [2:0] GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire [2:0] GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire [38:0] GEN_50;
  wire [5:0] GEN_51;
  wire [6:0] GEN_52;
  wire [1:0] GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire [1:0] GEN_57;
  wire [61:0] GEN_58;
  wire  GEN_59;
  wire [1:0] GEN_60;
  wire [61:0] GEN_61;
  wire  T_7617;
  wire [31:0] GEN_62;
  wire [39:0] GEN_63;
  wire  T_7619;
  wire  wb_dcache_miss;
  wire  T_7621;
  wire  T_7622;
  wire  T_7624;
  wire  T_7625;
  wire  replay_ex_structural;
  wire  replay_ex_load_use;
  wire  T_7626;
  wire  replay_ex;
  wire  T_7627;
  wire  T_7629;
  wire  ctrl_killx;
  wire  T_7630;
  wire [2:0] T_7636_0;
  wire [2:0] T_7636_1;
  wire [2:0] T_7636_2;
  wire [2:0] T_7636_3;
  wire  T_7638;
  wire  T_7639;
  wire  T_7640;
  wire  T_7641;
  wire  T_7644;
  wire  T_7645;
  wire  T_7646;
  wire  ex_slow_bypass;
  wire  T_7647;
  wire  T_7648;
  wire  ex_xcpt;
  wire [63:0] ex_cause;
  wire  mem_br_taken;
  wire [39:0] T_7650;
  wire  T_7651;
  wire  T_7654;
  wire  T_7655;
  wire  T_7656;
  wire [10:0] T_7658;
  wire [10:0] T_7659;
  wire [10:0] T_7660;
  wire [7:0] T_7664;
  wire [7:0] T_7665;
  wire [7:0] T_7666;
  wire  T_7672;
  wire  T_7673;
  wire  T_7675;
  wire  T_7676;
  wire  T_7677;
  wire  T_7678;
  wire  T_7679;
  wire [5:0] T_7684;
  wire [3:0] T_7691;
  wire [3:0] T_7694;
  wire [9:0] T_7711;
  wire [10:0] T_7712;
  wire  T_7713;
  wire [7:0] T_7714;
  wire [8:0] T_7715;
  wire [10:0] T_7716;
  wire  T_7717;
  wire [11:0] T_7718;
  wire [20:0] T_7719;
  wire [31:0] T_7720;
  wire [31:0] T_7721;
  wire [7:0] T_7736;
  wire  T_7747;
  wire  T_7748;
  wire  T_7749;
  wire [9:0] T_7781;
  wire [10:0] T_7782;
  wire  T_7783;
  wire [7:0] T_7784;
  wire [8:0] T_7785;
  wire [20:0] T_7789;
  wire [31:0] T_7790;
  wire [31:0] T_7791;
  wire [3:0] GEN_184;
  wire [31:0] T_7793;
  wire [31:0] T_7794;
  wire [39:0] GEN_185;
  wire [40:0] T_7795;
  wire [39:0] T_7796;
  wire [39:0] mem_br_target;
  wire [63:0] T_7797;
  wire [63:0] T_7798;
  wire [63:0] mem_int_wdata;
  wire [25:0] T_7799;
  wire [1:0] T_7800;
  wire [1:0] T_7801;
  wire [25:0] GEN_186;
  wire  T_7803;
  wire [25:0] GEN_187;
  wire  T_7805;
  wire  T_7806;
  wire [1:0] GEN_189;
  wire  T_7808;
  wire [25:0] T_7809;
  wire  GEN_190;
  wire [25:0] GEN_191;
  wire  T_7811;
  wire [1:0] GEN_192;
  wire [25:0] GEN_193;
  wire  T_7814;
  wire  T_7815;
  wire [1:0] GEN_195;
  wire  T_7817;
  wire  T_7818;
  wire  T_7819;
  wire  T_7820;
  wire [38:0] T_7821;
  wire [39:0] T_7822;
  wire [39:0] T_7823;
  wire [39:0] T_7824;
  wire [39:0] GEN_197;
  wire [39:0] T_7826;
  wire [39:0] T_7827;
  wire [39:0] mem_npc;
  wire  T_7828;
  wire  mem_wrong_npc;
  wire  mem_npc_misaligned;
  wire  T_7831;
  wire  mem_cfi;
  wire  T_7833;
  wire  mem_cfi_taken;
  wire  mem_misprediction;
  wire  T_7834;
  wire  want_take_pc_mem;
  wire  T_7836;
  wire  T_7837;
  wire  T_7839;
  wire  T_7842;
  wire  T_7845;
  wire  T_7848;
  wire [63:0] GEN_64;
  wire  T_7849;
  wire  T_7850;
  wire  T_7851;
  wire  T_7852;
  wire  T_7854;
  wire  T_7855;
  wire  T_7856;
  wire  T_7857;
  wire  T_7858;
  wire  T_7859;
  wire  T_7860;
  wire  T_7862;
  wire  T_7866;
  wire  T_7867;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire [38:0] GEN_68;
  wire [5:0] GEN_69;
  wire [6:0] GEN_70;
  wire [1:0] GEN_71;
  wire  T_7868;
  wire  T_7869;
  wire [63:0] GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire [1:0] GEN_81;
  wire [1:0] GEN_82;
  wire [2:0] GEN_83;
  wire  GEN_84;
  wire [3:0] GEN_85;
  wire  GEN_86;
  wire [4:0] GEN_87;
  wire [2:0] GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire [2:0] GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire [38:0] GEN_105;
  wire [5:0] GEN_106;
  wire [6:0] GEN_107;
  wire [1:0] GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire [31:0] GEN_111;
  wire [39:0] GEN_112;
  wire [63:0] GEN_113;
  wire [63:0] GEN_114;
  wire  T_7870;
  wire  T_7872;
  wire  T_7874;
  wire  T_7876;
  wire  T_7878;
  wire  T_7880;
  wire  T_7882;
  wire  T_7884;
  wire  T_7885;
  wire  T_7886;
  wire  T_7887;
  wire  T_7888;
  wire  mem_new_xcpt;
  wire [2:0] T_7889;
  wire [2:0] T_7890;
  wire [2:0] T_7891;
  wire [2:0] T_7892;
  wire [2:0] T_7893;
  wire [2:0] mem_new_cause;
  wire  T_7894;
  wire  T_7895;
  wire  mem_xcpt;
  wire [63:0] mem_cause;
  wire  dcache_kill_mem;
  wire  T_7897;
  wire  fpu_kill_mem;
  wire  T_7898;
  wire  replay_mem;
  wire  T_7899;
  wire  T_7900;
  wire  T_7902;
  wire  killm_common;
  wire  T_7903;
  reg  T_7904;
  reg [31:0] GEN_428;
  wire  T_7905;
  wire  T_7906;
  wire  ctrl_killm;
  wire  T_7908;
  wire  T_7910;
  wire  T_7911;
  wire  T_7914;
  wire  T_7918;
  wire  T_7919;
  wire [63:0] GEN_115;
  wire  T_7920;
  wire  T_7921;
  wire  T_7922;
  wire [63:0] T_7923;
  wire [63:0] GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire [1:0] GEN_125;
  wire [1:0] GEN_126;
  wire [2:0] GEN_127;
  wire  GEN_128;
  wire [3:0] GEN_129;
  wire  GEN_130;
  wire [4:0] GEN_131;
  wire [2:0] GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire [2:0] GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire [63:0] GEN_143;
  wire [63:0] GEN_144;
  wire [31:0] GEN_145;
  wire [39:0] GEN_146;
  wire  T_7924;
  wire  wb_set_sboard;
  wire  replay_wb_common;
  wire  T_7927;
  wire  wb_rocc_val;
  wire  T_7930;
  wire  T_7931;
  wire  replay_wb;
  wire  wb_xcpt;
  wire  T_7932;
  wire  T_7933;
  wire  GEN_147;
  wire  GEN_148;
  wire  T_7937;
  wire  dmem_resp_xpu;
  wire [7:0] dmem_resp_waddr;
  wire  dmem_resp_valid;
  wire  dmem_resp_replay;
  wire  T_7941;
  wire  T_7943;
  wire [63:0] ll_wdata;
  wire [7:0] ll_waddr;
  wire  T_7944;
  wire  ll_wen;
  wire  T_7945;
  wire  GEN_149;
  wire [7:0] GEN_150;
  wire  GEN_151;
  wire  T_7949;
  wire  T_7950;
  wire  T_7952;
  wire  wb_valid;
  wire  wb_wen;
  wire  rf_wen;
  wire [7:0] rf_waddr;
  wire  T_7953;
  wire  T_7954;
  wire [63:0] T_7955;
  wire [63:0] T_7956;
  wire [63:0] rf_wdata;
  wire [7:0] GEN_198;
  wire  T_7958;
  wire [4:0] T_7959;
  wire [4:0] T_7960;
  wire [7:0] GEN_199;
  wire  T_7962;
  wire [63:0] GEN_152;
  wire [7:0] GEN_200;
  wire  T_7963;
  wire [63:0] GEN_153;
  wire [63:0] GEN_159;
  wire [63:0] GEN_160;
  wire  GEN_163;
  wire [63:0] GEN_166;
  wire [63:0] GEN_167;
  wire [25:0] T_7964;
  wire [1:0] T_7965;
  wire [1:0] T_7966;
  wire  T_7968;
  wire  T_7970;
  wire  T_7971;
  wire  T_7973;
  wire [25:0] T_7974;
  wire  T_7976;
  wire  T_7979;
  wire  T_7980;
  wire  T_7982;
  wire  T_7983;
  wire  T_7984;
  wire  T_7985;
  wire [38:0] T_7986;
  wire [39:0] T_7987;
  wire [39:0] T_7988;
  wire [11:0] T_8005;
  wire [2:0] T_8006;
  wire  T_8008;
  wire  T_8009;
  wire  T_8011;
  wire  T_8012;
  wire  T_8014;
  wire  T_8015;
  reg [31:0] T_8017;
  reg [31:0] GEN_429;
  wire [255:0] GEN_214;
  wire [255:0] T_8020;
  wire [255:0] T_8022;
  wire [255:0] T_8023;
  wire [255:0] GEN_215;
  wire [255:0] T_8024;
  wire [255:0] GEN_168;
  wire [31:0] T_8026;
  wire  T_8027;
  wire  T_8028;
  wire [31:0] T_8029;
  wire  T_8030;
  wire  T_8031;
  wire [31:0] T_8032;
  wire  T_8033;
  wire  T_8034;
  wire  T_8035;
  wire  id_sboard_hazard;
  wire  T_8036;
  wire [31:0] GEN_216;
  wire [31:0] T_8038;
  wire [31:0] T_8040;
  wire [255:0] GEN_217;
  wire [255:0] T_8041;
  wire  T_8042;
  wire [255:0] GEN_169;
  wire  T_8043;
  wire  T_8044;
  wire  T_8045;
  wire  T_8046;
  wire  T_8047;
  wire  ex_cannot_bypass;
  wire  T_8048;
  wire  T_8049;
  wire  T_8050;
  wire  T_8051;
  wire  T_8052;
  wire  T_8053;
  wire  T_8054;
  wire  T_8055;
  wire  data_hazard_ex;
  wire  T_8057;
  wire  T_8059;
  wire  T_8060;
  wire  T_8061;
  wire  T_8063;
  wire  T_8064;
  wire  T_8065;
  wire  T_8066;
  wire  fp_data_hazard_ex;
  wire  T_8067;
  wire  T_8068;
  wire  id_ex_hazard;
  wire  T_8070;
  wire  T_8071;
  wire  T_8072;
  wire  T_8073;
  wire  T_8074;
  wire  mem_cannot_bypass;
  wire  T_8075;
  wire  T_8076;
  wire  T_8077;
  wire  T_8078;
  wire  T_8079;
  wire  T_8080;
  wire  T_8081;
  wire  T_8082;
  wire  data_hazard_mem;
  wire  T_8084;
  wire  T_8086;
  wire  T_8087;
  wire  T_8088;
  wire  T_8090;
  wire  T_8091;
  wire  T_8092;
  wire  T_8093;
  wire  fp_data_hazard_mem;
  wire  T_8094;
  wire  T_8095;
  wire  id_mem_hazard;
  wire  T_8096;
  wire  T_8097;
  wire  T_8098;
  wire  T_8099;
  wire  T_8100;
  wire  T_8101;
  wire  T_8102;
  wire  T_8103;
  wire  T_8104;
  wire  T_8105;
  wire  data_hazard_wb;
  wire  T_8107;
  wire  T_8109;
  wire  T_8110;
  wire  T_8111;
  wire  T_8113;
  wire  T_8114;
  wire  T_8115;
  wire  T_8116;
  wire  fp_data_hazard_wb;
  wire  T_8117;
  wire  T_8118;
  wire  id_wb_hazard;
  reg [31:0] T_8120;
  reg [31:0] GEN_430;
  wire  T_8122;
  wire  T_8123;
  wire  T_8124;
  wire [31:0] T_8128;
  wire [31:0] T_8129;
  wire [31:0] GEN_170;
  wire  T_8131;
  wire [255:0] T_8133;
  wire [255:0] T_8135;
  wire [255:0] T_8136;
  wire [255:0] GEN_220;
  wire [255:0] T_8137;
  wire  T_8138;
  wire [255:0] GEN_171;
  wire [31:0] T_8140;
  wire [31:0] T_8142;
  wire [31:0] T_8143;
  wire [255:0] GEN_222;
  wire [255:0] T_8144;
  wire  T_8145;
  wire [255:0] GEN_172;
  wire  T_8147;
  wire  T_8148;
  wire [31:0] T_8149;
  wire  T_8150;
  wire  T_8151;
  wire [31:0] T_8152;
  wire  T_8153;
  wire  T_8154;
  wire [31:0] T_8155;
  wire  T_8156;
  wire  T_8157;
  wire [31:0] T_8158;
  wire  T_8159;
  wire  T_8160;
  wire  T_8161;
  wire  T_8162;
  wire  T_8163;
  wire  id_stall_fpu;
  reg  dcache_blocked;
  reg [31:0] GEN_431;
  wire  T_8167;
  wire  T_8168;
  wire  T_8169;
  wire  T_8170;
  wire  T_8171;
  wire  T_8172;
  wire  T_8173;
  wire  T_8174;
  wire  T_8175;
  wire  T_8183;
  wire  ctrl_stalld;
  wire  T_8185;
  wire  T_8186;
  wire  T_8187;
  wire  T_8188;
  wire  T_8189;
  wire [39:0] T_8190;
  wire [39:0] T_8191;
  wire  T_8192;
  wire  T_8194;
  wire  T_8195;
  wire  T_8197;
  wire  T_8198;
  wire  T_8199;
  wire  T_8202;
  wire  T_8203;
  wire  T_8204;
  wire  T_8207;
  wire  T_8208;
  wire [4:0] T_8209;
  wire [4:0] T_8212;
  wire [4:0] GEN_223;
  wire  T_8213;
  wire  T_8214;
  wire  T_8215;
  wire  T_8218;
  wire  T_8219;
  wire  T_8222;
  wire  T_8225;
  wire  T_8226;
  wire  T_8227;
  wire  T_8230;
  wire  T_8231;
  wire  T_8232;
  wire [5:0] ex_dcache_tag;
  wire [25:0] T_8234;
  wire [1:0] T_8235;
  wire [1:0] T_8236;
  wire  T_8238;
  wire  T_8240;
  wire  T_8241;
  wire  T_8243;
  wire [25:0] T_8244;
  wire  T_8246;
  wire  T_8249;
  wire  T_8250;
  wire  T_8252;
  wire  T_8253;
  wire  T_8254;
  wire  T_8255;
  wire [38:0] T_8256;
  wire [39:0] T_8257;
  wire [63:0] T_8259;
  wire  T_8262;
  wire [6:0] T_8281_funct;
  wire [4:0] T_8281_rs2;
  wire [4:0] T_8281_rs1;
  wire  T_8281_xd;
  wire  T_8281_xs1;
  wire  T_8281_xs2;
  wire [4:0] T_8281_rd;
  wire [6:0] T_8281_opcode;
  wire [31:0] T_8291;
  wire [6:0] T_8292;
  wire [4:0] T_8293;
  wire  T_8294;
  wire  T_8295;
  wire  T_8296;
  wire [4:0] T_8297;
  wire [4:0] T_8298;
  wire [6:0] T_8299;
  wire [31:0] T_8300;
  wire [7:0] T_8302;
  wire [4:0] T_8303;
  reg [63:0] T_8304;
  reg [63:0] GEN_432;
  reg [63:0] T_8305;
  reg [63:0] GEN_433;
  wire [4:0] T_8306;
  reg [63:0] T_8307;
  reg [63:0] GEN_434;
  reg [63:0] T_8308;
  reg [63:0] GEN_435;
  wire  T_8310;
  reg  GEN_154;
  reg [31:0] GEN_436;
  reg [63:0] GEN_155;
  reg [63:0] GEN_437;
  reg  GEN_156;
  reg [31:0] GEN_438;
  reg [4:0] GEN_157;
  reg [31:0] GEN_439;
  reg  GEN_158;
  reg [31:0] GEN_440;
  reg  GEN_161;
  reg [31:0] GEN_441;
  reg  GEN_162;
  reg [31:0] GEN_442;
  reg  GEN_164;
  reg [31:0] GEN_443;
  reg  GEN_165;
  reg [31:0] GEN_444;
  reg  GEN_174;
  reg [31:0] GEN_445;
  reg  GEN_175;
  reg [31:0] GEN_446;
  reg  GEN_177;
  reg [31:0] GEN_447;
  reg  GEN_178;
  reg [31:0] GEN_448;
  reg  GEN_179;
  reg [31:0] GEN_449;
  reg  GEN_181;
  reg [31:0] GEN_450;
  reg  GEN_183;
  reg [31:0] GEN_451;
  reg  GEN_188;
  reg [31:0] GEN_452;
  reg  GEN_194;
  reg [31:0] GEN_453;
  reg  GEN_196;
  reg [31:0] GEN_454;
  reg  GEN_201;
  reg [31:0] GEN_455;
  reg [2:0] GEN_202;
  reg [31:0] GEN_456;
  reg [1:0] GEN_203;
  reg [31:0] GEN_457;
  reg [64:0] GEN_204;
  reg [95:0] GEN_458;
  reg [64:0] GEN_205;
  reg [95:0] GEN_459;
  reg [64:0] GEN_206;
  reg [95:0] GEN_460;
  reg  GEN_207;
  reg [31:0] GEN_461;
  reg  GEN_208;
  reg [31:0] GEN_462;
  reg  GEN_209;
  reg [31:0] GEN_463;
  reg  GEN_210;
  reg [31:0] GEN_464;
  reg  GEN_211;
  reg [31:0] GEN_465;
  reg [39:0] GEN_212;
  reg [63:0] GEN_466;
  reg [8:0] GEN_213;
  reg [31:0] GEN_467;
  reg [4:0] GEN_218;
  reg [31:0] GEN_468;
  reg [2:0] GEN_219;
  reg [31:0] GEN_469;
  reg [63:0] GEN_221;
  reg [63:0] GEN_470;
  reg  GEN_224;
  reg [31:0] GEN_471;
  reg  GEN_225;
  reg [31:0] GEN_472;
  reg [63:0] GEN_226;
  reg [63:0] GEN_473;
  reg [63:0] GEN_227;
  reg [63:0] GEN_474;
  reg  GEN_228;
  reg [31:0] GEN_475;
  reg  GEN_229;
  reg [31:0] GEN_476;
  reg  GEN_230;
  reg [31:0] GEN_477;
  reg  GEN_231;
  reg [31:0] GEN_478;
  reg  GEN_232;
  reg [31:0] GEN_479;
  reg  GEN_233;
  reg [31:0] GEN_480;
  reg  GEN_234;
  reg [31:0] GEN_481;
  reg  GEN_235;
  reg [31:0] GEN_482;
  reg [2:0] GEN_236;
  reg [31:0] GEN_483;
  reg [1:0] GEN_237;
  reg [31:0] GEN_484;
  reg [2:0] GEN_238;
  reg [31:0] GEN_485;
  reg  GEN_239;
  reg [31:0] GEN_486;
  reg [3:0] GEN_240;
  reg [31:0] GEN_487;
  reg [63:0] GEN_241;
  reg [63:0] GEN_488;
  reg  GEN_242;
  reg [31:0] GEN_489;
  reg  GEN_243;
  reg [31:0] GEN_490;
  reg [64:0] GEN_244;
  reg [95:0] GEN_491;
  reg [4:0] GEN_245;
  reg [31:0] GEN_492;
  reg  GEN_246;
  reg [31:0] GEN_493;
  reg  GEN_247;
  reg [31:0] GEN_494;
  reg  GEN_248;
  reg [31:0] GEN_495;
  reg [4:0] GEN_249;
  reg [31:0] GEN_496;
  reg [63:0] GEN_250;
  reg [63:0] GEN_497;
  reg  GEN_251;
  reg [31:0] GEN_498;
  reg [39:0] GEN_252;
  reg [63:0] GEN_499;
  reg [8:0] GEN_253;
  reg [31:0] GEN_500;
  reg [4:0] GEN_254;
  reg [31:0] GEN_501;
  reg [2:0] GEN_255;
  reg [31:0] GEN_502;
  reg  GEN_256;
  reg [31:0] GEN_503;
  reg [63:0] GEN_257;
  reg [63:0] GEN_504;
  reg  GEN_258;
  reg [31:0] GEN_505;
  reg [63:0] GEN_259;
  reg [63:0] GEN_506;
  reg  GEN_260;
  reg [31:0] GEN_507;
  reg  GEN_261;
  reg [31:0] GEN_508;
  reg  GEN_262;
  reg [31:0] GEN_509;
  reg [25:0] GEN_263;
  reg [31:0] GEN_510;
  reg [1:0] GEN_264;
  reg [31:0] GEN_511;
  reg [2:0] GEN_265;
  reg [31:0] GEN_512;
  reg  GEN_266;
  reg [31:0] GEN_513;
  reg [2:0] GEN_267;
  reg [31:0] GEN_514;
  reg [11:0] GEN_268;
  reg [31:0] GEN_515;
  reg [63:0] GEN_269;
  reg [63:0] GEN_516;
  reg  GEN_270;
  reg [31:0] GEN_517;
  reg  GEN_271;
  reg [31:0] GEN_518;
  reg [4:0] GEN_272;
  reg [31:0] GEN_519;
  reg  GEN_273;
  reg [31:0] GEN_520;
  reg  GEN_274;
  reg [31:0] GEN_521;
  reg  GEN_275;
  reg [31:0] GEN_522;
  reg  GEN_276;
  reg [31:0] GEN_523;
  reg  GEN_277;
  reg [31:0] GEN_524;
  reg  GEN_278;
  reg [31:0] GEN_525;
  reg  GEN_279;
  reg [31:0] GEN_526;
  reg  GEN_280;
  reg [31:0] GEN_527;
  reg  GEN_281;
  reg [31:0] GEN_528;
  reg  GEN_282;
  reg [31:0] GEN_529;
  reg  GEN_283;
  reg [31:0] GEN_530;
  reg  GEN_284;
  reg [31:0] GEN_531;
  reg  GEN_285;
  reg [31:0] GEN_532;
  reg  GEN_286;
  reg [31:0] GEN_533;
  reg  GEN_287;
  reg [31:0] GEN_534;
  reg  GEN_288;
  reg [31:0] GEN_535;
  reg [2:0] GEN_289;
  reg [31:0] GEN_536;
  reg [1:0] GEN_290;
  reg [31:0] GEN_537;
  reg [64:0] GEN_291;
  reg [95:0] GEN_538;
  reg [64:0] GEN_292;
  reg [95:0] GEN_539;
  reg [64:0] GEN_293;
  reg [95:0] GEN_540;
  reg  GEN_294;
  reg [31:0] GEN_541;
  CSRFile csr (
    .clk(csr_clk),
    .reset(csr_reset),
    .io_prci_reset(csr_io_prci_reset),
    .io_prci_id(csr_io_prci_id),
    .io_prci_interrupts_mtip(csr_io_prci_interrupts_mtip),
    .io_prci_interrupts_meip(csr_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(csr_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(csr_io_prci_interrupts_debug),
    .io_prci_interrupts_msip(csr_io_prci_interrupts_msip),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_csr_stall(csr_io_csr_stall),
    .io_csr_xcpt(csr_io_csr_xcpt),
    .io_eret(csr_io_eret),
    .io_prv(csr_io_prv),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero3(csr_io_status_zero3),
    .io_status_sd_rv32(csr_io_status_sd_rv32),
    .io_status_zero2(csr_io_status_zero2),
    .io_status_vm(csr_io_status_vm),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_pum(csr_io_status_pum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_ptbr(csr_io_ptbr),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_uarch_counters_0(csr_io_uarch_counters_0),
    .io_uarch_counters_1(csr_io_uarch_counters_1),
    .io_uarch_counters_2(csr_io_uarch_counters_2),
    .io_uarch_counters_3(csr_io_uarch_counters_3),
    .io_uarch_counters_4(csr_io_uarch_counters_4),
    .io_uarch_counters_5(csr_io_uarch_counters_5),
    .io_uarch_counters_6(csr_io_uarch_counters_6),
    .io_uarch_counters_7(csr_io_uarch_counters_7),
    .io_uarch_counters_8(csr_io_uarch_counters_8),
    .io_uarch_counters_9(csr_io_uarch_counters_9),
    .io_uarch_counters_10(csr_io_uarch_counters_10),
    .io_uarch_counters_11(csr_io_uarch_counters_11),
    .io_uarch_counters_12(csr_io_uarch_counters_12),
    .io_uarch_counters_13(csr_io_uarch_counters_13),
    .io_uarch_counters_14(csr_io_uarch_counters_14),
    .io_uarch_counters_15(csr_io_uarch_counters_15),
    .io_cause(csr_io_cause),
    .io_pc(csr_io_pc),
    .io_badaddr(csr_io_badaddr),
    .io_fatc(csr_io_fatc),
    .io_time(csr_io_time),
    .io_fcsr_rm(csr_io_fcsr_rm),
    .io_fcsr_flags_valid(csr_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(csr_io_fcsr_flags_bits),
    .io_rocc_cmd_ready(csr_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(csr_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(csr_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(csr_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(csr_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(csr_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(csr_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(csr_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(csr_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(csr_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(csr_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(csr_io_rocc_cmd_bits_rs2),
    .io_rocc_resp_ready(csr_io_rocc_resp_ready),
    .io_rocc_resp_valid(csr_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(csr_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(csr_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(csr_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(csr_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(csr_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(csr_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(csr_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(csr_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(csr_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(csr_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(csr_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(csr_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(csr_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(csr_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(csr_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(csr_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(csr_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(csr_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(csr_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(csr_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(csr_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(csr_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(csr_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(csr_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(csr_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(csr_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(csr_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(csr_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(csr_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(csr_io_rocc_mem_ordered),
    .io_rocc_busy(csr_io_rocc_busy),
    .io_rocc_status_debug(csr_io_rocc_status_debug),
    .io_rocc_status_prv(csr_io_rocc_status_prv),
    .io_rocc_status_sd(csr_io_rocc_status_sd),
    .io_rocc_status_zero3(csr_io_rocc_status_zero3),
    .io_rocc_status_sd_rv32(csr_io_rocc_status_sd_rv32),
    .io_rocc_status_zero2(csr_io_rocc_status_zero2),
    .io_rocc_status_vm(csr_io_rocc_status_vm),
    .io_rocc_status_zero1(csr_io_rocc_status_zero1),
    .io_rocc_status_pum(csr_io_rocc_status_pum),
    .io_rocc_status_mprv(csr_io_rocc_status_mprv),
    .io_rocc_status_xs(csr_io_rocc_status_xs),
    .io_rocc_status_fs(csr_io_rocc_status_fs),
    .io_rocc_status_mpp(csr_io_rocc_status_mpp),
    .io_rocc_status_hpp(csr_io_rocc_status_hpp),
    .io_rocc_status_spp(csr_io_rocc_status_spp),
    .io_rocc_status_mpie(csr_io_rocc_status_mpie),
    .io_rocc_status_hpie(csr_io_rocc_status_hpie),
    .io_rocc_status_spie(csr_io_rocc_status_spie),
    .io_rocc_status_upie(csr_io_rocc_status_upie),
    .io_rocc_status_mie(csr_io_rocc_status_mie),
    .io_rocc_status_hie(csr_io_rocc_status_hie),
    .io_rocc_status_sie(csr_io_rocc_status_sie),
    .io_rocc_status_uie(csr_io_rocc_status_uie),
    .io_rocc_interrupt(csr_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(csr_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(csr_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(csr_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(csr_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(csr_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(csr_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(csr_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(csr_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(csr_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(csr_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(csr_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(csr_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(csr_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(csr_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(csr_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(csr_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(csr_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(csr_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(csr_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(csr_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(csr_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(csr_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(csr_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(csr_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(csr_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(csr_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(csr_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(csr_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(csr_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(csr_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(csr_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(csr_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(csr_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(csr_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(csr_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(csr_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(csr_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(csr_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(csr_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(csr_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(csr_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(csr_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(csr_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(csr_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(csr_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(csr_io_rocc_exception),
    .io_rocc_csr_waddr(csr_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(csr_io_rocc_csr_wdata),
    .io_rocc_csr_wen(csr_io_rocc_csr_wen),
    .io_rocc_host_id(csr_io_rocc_host_id),
    .io_interrupt(csr_io_interrupt),
    .io_interrupt_cause(csr_io_interrupt_cause),
    .io_bp_0_control_tdrtype(csr_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(csr_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(csr_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(csr_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(csr_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(csr_io_bp_0_control_m),
    .io_bp_0_control_h(csr_io_bp_0_control_h),
    .io_bp_0_control_s(csr_io_bp_0_control_s),
    .io_bp_0_control_u(csr_io_bp_0_control_u),
    .io_bp_0_control_r(csr_io_bp_0_control_r),
    .io_bp_0_control_w(csr_io_bp_0_control_w),
    .io_bp_0_control_x(csr_io_bp_0_control_x),
    .io_bp_0_address(csr_io_bp_0_address)
  );
  BreakpointUnit bpu (
    .clk(bpu_clk),
    .reset(bpu_reset),
    .io_status_debug(bpu_io_status_debug),
    .io_status_prv(bpu_io_status_prv),
    .io_status_sd(bpu_io_status_sd),
    .io_status_zero3(bpu_io_status_zero3),
    .io_status_sd_rv32(bpu_io_status_sd_rv32),
    .io_status_zero2(bpu_io_status_zero2),
    .io_status_vm(bpu_io_status_vm),
    .io_status_zero1(bpu_io_status_zero1),
    .io_status_pum(bpu_io_status_pum),
    .io_status_mprv(bpu_io_status_mprv),
    .io_status_xs(bpu_io_status_xs),
    .io_status_fs(bpu_io_status_fs),
    .io_status_mpp(bpu_io_status_mpp),
    .io_status_hpp(bpu_io_status_hpp),
    .io_status_spp(bpu_io_status_spp),
    .io_status_mpie(bpu_io_status_mpie),
    .io_status_hpie(bpu_io_status_hpie),
    .io_status_spie(bpu_io_status_spie),
    .io_status_upie(bpu_io_status_upie),
    .io_status_mie(bpu_io_status_mie),
    .io_status_hie(bpu_io_status_hie),
    .io_status_sie(bpu_io_status_sie),
    .io_status_uie(bpu_io_status_uie),
    .io_bp_0_control_tdrtype(bpu_io_bp_0_control_tdrtype),
    .io_bp_0_control_bpamaskmax(bpu_io_bp_0_control_bpamaskmax),
    .io_bp_0_control_reserved(bpu_io_bp_0_control_reserved),
    .io_bp_0_control_bpaction(bpu_io_bp_0_control_bpaction),
    .io_bp_0_control_bpmatch(bpu_io_bp_0_control_bpmatch),
    .io_bp_0_control_m(bpu_io_bp_0_control_m),
    .io_bp_0_control_h(bpu_io_bp_0_control_h),
    .io_bp_0_control_s(bpu_io_bp_0_control_s),
    .io_bp_0_control_u(bpu_io_bp_0_control_u),
    .io_bp_0_control_r(bpu_io_bp_0_control_r),
    .io_bp_0_control_w(bpu_io_bp_0_control_w),
    .io_bp_0_control_x(bpu_io_bp_0_control_x),
    .io_bp_0_address(bpu_io_bp_0_address),
    .io_pc(bpu_io_pc),
    .io_ea(bpu_io_ea),
    .io_xcpt_if(bpu_io_xcpt_if),
    .io_xcpt_ld(bpu_io_xcpt_ld),
    .io_xcpt_st(bpu_io_xcpt_st)
  );
  ALU alu (
    .clk(alu_clk),
    .reset(alu_reset),
    .io_dw(alu_io_dw),
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    .io_cmp_out(alu_io_cmp_out)
  );
  MulDiv div (
    .clk(div_clk),
    .reset(div_reset),
    .io_req_ready(div_io_req_ready),
    .io_req_valid(div_io_req_valid),
    .io_req_bits_fn(div_io_req_bits_fn),
    .io_req_bits_dw(div_io_req_bits_dw),
    .io_req_bits_in1(div_io_req_bits_in1),
    .io_req_bits_in2(div_io_req_bits_in2),
    .io_req_bits_tag(div_io_req_bits_tag),
    .io_kill(div_io_kill),
    .io_resp_ready(div_io_resp_ready),
    .io_resp_valid(div_io_resp_valid),
    .io_resp_bits_data(div_io_resp_bits_data),
    .io_resp_bits_tag(div_io_resp_bits_tag)
  );
  assign io_imem_req_valid = take_pc_mem_wb;
  assign io_imem_req_bits_pc = T_8191;
  assign io_imem_resp_ready = T_8199;
  assign io_imem_btb_update_valid = T_8207;
  assign io_imem_btb_update_bits_prediction_valid = mem_reg_btb_hit;
  assign io_imem_btb_update_bits_prediction_bits_taken = mem_reg_btb_resp_taken;
  assign io_imem_btb_update_bits_prediction_bits_mask = mem_reg_btb_resp_mask;
  assign io_imem_btb_update_bits_prediction_bits_bridx = mem_reg_btb_resp_bridx;
  assign io_imem_btb_update_bits_prediction_bits_target = mem_reg_btb_resp_target;
  assign io_imem_btb_update_bits_prediction_bits_entry = mem_reg_btb_resp_entry;
  assign io_imem_btb_update_bits_prediction_bits_bht_history = mem_reg_btb_resp_bht_history;
  assign io_imem_btb_update_bits_prediction_bits_bht_value = mem_reg_btb_resp_bht_value;
  assign io_imem_btb_update_bits_pc = mem_reg_pc[38:0];
  assign io_imem_btb_update_bits_target = io_imem_req_bits_pc[38:0];
  assign io_imem_btb_update_bits_taken = GEN_154;
  assign io_imem_btb_update_bits_isJump = T_8208;
  assign io_imem_btb_update_bits_isReturn = T_8214;
  assign io_imem_btb_update_bits_br_pc = mem_reg_pc[38:0];
  assign io_imem_bht_update_valid = T_8218;
  assign io_imem_bht_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_bht_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_bht_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_bht_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_bht_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_bht_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_bht_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_bht_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_bht_update_bits_pc = mem_reg_pc[38:0];
  assign io_imem_bht_update_bits_taken = mem_br_taken;
  assign io_imem_bht_update_bits_mispredict = mem_wrong_npc;
  assign io_imem_ras_update_valid = T_8225;
  assign io_imem_ras_update_bits_isCall = T_8227;
  assign io_imem_ras_update_bits_isReturn = io_imem_btb_update_bits_isReturn;
  assign io_imem_ras_update_bits_returnAddr = mem_int_wdata[38:0];
  assign io_imem_ras_update_bits_prediction_valid = io_imem_btb_update_bits_prediction_valid;
  assign io_imem_ras_update_bits_prediction_bits_taken = io_imem_btb_update_bits_prediction_bits_taken;
  assign io_imem_ras_update_bits_prediction_bits_mask = io_imem_btb_update_bits_prediction_bits_mask;
  assign io_imem_ras_update_bits_prediction_bits_bridx = io_imem_btb_update_bits_prediction_bits_bridx;
  assign io_imem_ras_update_bits_prediction_bits_target = io_imem_btb_update_bits_prediction_bits_target;
  assign io_imem_ras_update_bits_prediction_bits_entry = io_imem_btb_update_bits_prediction_bits_entry;
  assign io_imem_ras_update_bits_prediction_bits_bht_history = io_imem_btb_update_bits_prediction_bits_bht_history;
  assign io_imem_ras_update_bits_prediction_bits_bht_value = io_imem_btb_update_bits_prediction_bits_bht_value;
  assign io_imem_flush_icache = T_8195;
  assign io_imem_flush_tlb = csr_io_fatc;
  assign io_dmem_req_valid = T_8232;
  assign io_dmem_req_bits_addr = T_8257;
  assign io_dmem_req_bits_tag = {{3'd0}, ex_dcache_tag};
  assign io_dmem_req_bits_cmd = ex_ctrl_mem_cmd;
  assign io_dmem_req_bits_typ = ex_ctrl_mem_type;
  assign io_dmem_req_bits_phys = 1'h0;
  assign io_dmem_req_bits_data = GEN_155;
  assign io_dmem_s1_kill = T_7906;
  assign io_dmem_s1_data = T_8259;
  assign io_dmem_invalidate_lr = wb_xcpt;
  assign io_ptw_ptbr = csr_io_ptbr[19:0];
  assign io_ptw_invalidate = csr_io_fatc;
  assign io_ptw_status_debug = csr_io_status_debug;
  assign io_ptw_status_prv = csr_io_status_prv;
  assign io_ptw_status_sd = csr_io_status_sd;
  assign io_ptw_status_zero3 = csr_io_status_zero3;
  assign io_ptw_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_ptw_status_zero2 = csr_io_status_zero2;
  assign io_ptw_status_vm = csr_io_status_vm;
  assign io_ptw_status_zero1 = csr_io_status_zero1;
  assign io_ptw_status_pum = csr_io_status_pum;
  assign io_ptw_status_mprv = csr_io_status_mprv;
  assign io_ptw_status_xs = csr_io_status_xs;
  assign io_ptw_status_fs = csr_io_status_fs;
  assign io_ptw_status_mpp = csr_io_status_mpp;
  assign io_ptw_status_hpp = csr_io_status_hpp;
  assign io_ptw_status_spp = csr_io_status_spp;
  assign io_ptw_status_mpie = csr_io_status_mpie;
  assign io_ptw_status_hpie = csr_io_status_hpie;
  assign io_ptw_status_spie = csr_io_status_spie;
  assign io_ptw_status_upie = csr_io_status_upie;
  assign io_ptw_status_mie = csr_io_status_mie;
  assign io_ptw_status_hie = csr_io_status_hie;
  assign io_ptw_status_sie = csr_io_status_sie;
  assign io_ptw_status_uie = csr_io_status_uie;
  assign io_fpu_inst = io_imem_resp_bits_data_0;
  assign io_fpu_fromint_data = T_7484;
  assign io_fpu_fcsr_rm = csr_io_fcsr_rm;
  assign io_fpu_dmem_resp_val = T_8231;
  assign io_fpu_dmem_resp_type = io_dmem_resp_bits_typ;
  assign io_fpu_dmem_resp_tag = dmem_resp_waddr[4:0];
  assign io_fpu_dmem_resp_data = io_dmem_resp_bits_data_word_bypass;
  assign io_fpu_valid = T_8230;
  assign io_fpu_killx = ctrl_killx;
  assign io_fpu_killm = killm_common;
  assign io_fpu_cp_req_valid = GEN_156;
  assign io_fpu_cp_req_bits_cmd = GEN_157;
  assign io_fpu_cp_req_bits_ldst = GEN_158;
  assign io_fpu_cp_req_bits_wen = GEN_161;
  assign io_fpu_cp_req_bits_ren1 = GEN_162;
  assign io_fpu_cp_req_bits_ren2 = GEN_164;
  assign io_fpu_cp_req_bits_ren3 = GEN_165;
  assign io_fpu_cp_req_bits_swap12 = GEN_174;
  assign io_fpu_cp_req_bits_swap23 = GEN_175;
  assign io_fpu_cp_req_bits_single = GEN_177;
  assign io_fpu_cp_req_bits_fromint = GEN_178;
  assign io_fpu_cp_req_bits_toint = GEN_179;
  assign io_fpu_cp_req_bits_fastpipe = GEN_181;
  assign io_fpu_cp_req_bits_fma = GEN_183;
  assign io_fpu_cp_req_bits_div = GEN_188;
  assign io_fpu_cp_req_bits_sqrt = GEN_194;
  assign io_fpu_cp_req_bits_round = GEN_196;
  assign io_fpu_cp_req_bits_wflags = GEN_201;
  assign io_fpu_cp_req_bits_rm = GEN_202;
  assign io_fpu_cp_req_bits_typ = GEN_203;
  assign io_fpu_cp_req_bits_in1 = GEN_204;
  assign io_fpu_cp_req_bits_in2 = GEN_205;
  assign io_fpu_cp_req_bits_in3 = GEN_206;
  assign io_fpu_cp_resp_ready = GEN_207;
  assign io_rocc_cmd_valid = wb_rocc_val;
  assign io_rocc_cmd_bits_inst_funct = T_8281_funct;
  assign io_rocc_cmd_bits_inst_rs2 = T_8281_rs2;
  assign io_rocc_cmd_bits_inst_rs1 = T_8281_rs1;
  assign io_rocc_cmd_bits_inst_xd = T_8281_xd;
  assign io_rocc_cmd_bits_inst_xs1 = T_8281_xs1;
  assign io_rocc_cmd_bits_inst_xs2 = T_8281_xs2;
  assign io_rocc_cmd_bits_inst_rd = T_8281_rd;
  assign io_rocc_cmd_bits_inst_opcode = T_8281_opcode;
  assign io_rocc_cmd_bits_rs1 = wb_reg_wdata;
  assign io_rocc_cmd_bits_rs2 = wb_reg_rs2;
  assign io_rocc_resp_ready = GEN_208;
  assign io_rocc_mem_req_ready = GEN_209;
  assign io_rocc_mem_s2_nack = GEN_210;
  assign io_rocc_mem_resp_valid = GEN_211;
  assign io_rocc_mem_resp_bits_addr = GEN_212;
  assign io_rocc_mem_resp_bits_tag = GEN_213;
  assign io_rocc_mem_resp_bits_cmd = GEN_218;
  assign io_rocc_mem_resp_bits_typ = GEN_219;
  assign io_rocc_mem_resp_bits_data = GEN_221;
  assign io_rocc_mem_resp_bits_replay = GEN_224;
  assign io_rocc_mem_resp_bits_has_data = GEN_225;
  assign io_rocc_mem_resp_bits_data_word_bypass = GEN_226;
  assign io_rocc_mem_resp_bits_store_data = GEN_227;
  assign io_rocc_mem_replay_next = GEN_228;
  assign io_rocc_mem_xcpt_ma_ld = GEN_229;
  assign io_rocc_mem_xcpt_ma_st = GEN_230;
  assign io_rocc_mem_xcpt_pf_ld = GEN_231;
  assign io_rocc_mem_xcpt_pf_st = GEN_232;
  assign io_rocc_mem_ordered = GEN_233;
  assign io_rocc_status_debug = csr_io_status_debug;
  assign io_rocc_status_prv = csr_io_status_prv;
  assign io_rocc_status_sd = csr_io_status_sd;
  assign io_rocc_status_zero3 = csr_io_status_zero3;
  assign io_rocc_status_sd_rv32 = csr_io_status_sd_rv32;
  assign io_rocc_status_zero2 = csr_io_status_zero2;
  assign io_rocc_status_vm = csr_io_status_vm;
  assign io_rocc_status_zero1 = csr_io_status_zero1;
  assign io_rocc_status_pum = csr_io_status_pum;
  assign io_rocc_status_mprv = csr_io_status_mprv;
  assign io_rocc_status_xs = csr_io_status_xs;
  assign io_rocc_status_fs = csr_io_status_fs;
  assign io_rocc_status_mpp = csr_io_status_mpp;
  assign io_rocc_status_hpp = csr_io_status_hpp;
  assign io_rocc_status_spp = csr_io_status_spp;
  assign io_rocc_status_mpie = csr_io_status_mpie;
  assign io_rocc_status_hpie = csr_io_status_hpie;
  assign io_rocc_status_spie = csr_io_status_spie;
  assign io_rocc_status_upie = csr_io_status_upie;
  assign io_rocc_status_mie = csr_io_status_mie;
  assign io_rocc_status_hie = csr_io_status_hie;
  assign io_rocc_status_sie = csr_io_status_sie;
  assign io_rocc_status_uie = csr_io_status_uie;
  assign io_rocc_autl_acquire_ready = GEN_234;
  assign io_rocc_autl_grant_valid = GEN_235;
  assign io_rocc_autl_grant_bits_addr_beat = GEN_236;
  assign io_rocc_autl_grant_bits_client_xact_id = GEN_237;
  assign io_rocc_autl_grant_bits_manager_xact_id = GEN_238;
  assign io_rocc_autl_grant_bits_is_builtin_type = GEN_239;
  assign io_rocc_autl_grant_bits_g_type = GEN_240;
  assign io_rocc_autl_grant_bits_data = GEN_241;
  assign io_rocc_fpu_req_ready = GEN_242;
  assign io_rocc_fpu_resp_valid = GEN_243;
  assign io_rocc_fpu_resp_bits_data = GEN_244;
  assign io_rocc_fpu_resp_bits_exc = GEN_245;
  assign io_rocc_exception = T_8262;
  assign io_rocc_csr_waddr = csr_io_rocc_csr_waddr;
  assign io_rocc_csr_wdata = csr_io_rocc_csr_wdata;
  assign io_rocc_csr_wen = csr_io_rocc_csr_wen;
  assign io_rocc_host_id = GEN_246;
  assign take_pc_mem = T_7837;
  assign take_pc_wb = T_7933;
  assign take_pc_mem_wb = take_pc_wb | take_pc_mem;
  assign id_ctrl_legal = T_6784;
  assign id_ctrl_fp = T_6795;
  assign id_ctrl_rocc = 1'h0;
  assign id_ctrl_branch = T_6800;
  assign id_ctrl_jal = T_6806;
  assign id_ctrl_jalr = T_6812;
  assign id_ctrl_rxs2 = T_6830;
  assign id_ctrl_rxs1 = T_6856;
  assign id_ctrl_sel_alu2 = T_6900;
  assign id_ctrl_sel_alu1 = T_6926;
  assign id_ctrl_sel_imm = T_6962;
  assign id_ctrl_alu_dw = T_6973;
  assign id_ctrl_alu_fn = T_7057;
  assign id_ctrl_mem = T_7078;
  assign id_ctrl_mem_cmd = T_7138;
  assign id_ctrl_mem_type = T_7158;
  assign id_ctrl_rfs1 = T_7174;
  assign id_ctrl_rfs2 = T_7191;
  assign id_ctrl_rfs3 = T_7170;
  assign id_ctrl_wfd = T_7206;
  assign id_ctrl_div = T_7210;
  assign id_ctrl_wxd = T_7248;
  assign id_ctrl_csr = T_7268;
  assign id_ctrl_fence_i = T_7272;
  assign id_ctrl_fence = T_7278;
  assign id_ctrl_amo = T_7284;
  assign T_6584 = io_imem_resp_bits_data_0 & 32'h207f;
  assign T_6586 = T_6584 == 32'h3;
  assign T_6588 = io_imem_resp_bits_data_0 & 32'h106f;
  assign T_6590 = T_6588 == 32'h3;
  assign T_6592 = io_imem_resp_bits_data_0 & 32'h607f;
  assign T_6594 = T_6592 == 32'hf;
  assign T_6596 = io_imem_resp_bits_data_0 & 32'h7077;
  assign T_6598 = T_6596 == 32'h13;
  assign T_6600 = io_imem_resp_bits_data_0 & 32'h5f;
  assign T_6602 = T_6600 == 32'h17;
  assign T_6604 = io_imem_resp_bits_data_0 & 32'hfc00007f;
  assign T_6606 = T_6604 == 32'h33;
  assign T_6608 = io_imem_resp_bits_data_0 & 32'hbe007077;
  assign T_6610 = T_6608 == 32'h33;
  assign T_6612 = io_imem_resp_bits_data_0 & 32'h4000073;
  assign T_6614 = T_6612 == 32'h43;
  assign T_6616 = io_imem_resp_bits_data_0 & 32'he400007f;
  assign T_6618 = T_6616 == 32'h53;
  assign T_6620 = io_imem_resp_bits_data_0 & 32'h707b;
  assign T_6622 = T_6620 == 32'h63;
  assign T_6624 = io_imem_resp_bits_data_0 & 32'h7f;
  assign T_6626 = T_6624 == 32'h6f;
  assign T_6628 = io_imem_resp_bits_data_0 & 32'hffefffff;
  assign T_6630 = T_6628 == 32'h73;
  assign T_6632 = io_imem_resp_bits_data_0 & 32'hfc00305f;
  assign T_6634 = T_6632 == 32'h1013;
  assign T_6636 = io_imem_resp_bits_data_0 & 32'hfe00305f;
  assign T_6638 = T_6636 == 32'h101b;
  assign T_6640 = io_imem_resp_bits_data_0 & 32'h605b;
  assign T_6642 = T_6640 == 32'h2003;
  assign T_6646 = T_6584 == 32'h2013;
  assign T_6648 = io_imem_resp_bits_data_0 & 32'h1800607f;
  assign T_6650 = T_6648 == 32'h202f;
  assign T_6654 = T_6584 == 32'h2073;
  assign T_6656 = io_imem_resp_bits_data_0 & 32'hbc00707f;
  assign T_6658 = T_6656 == 32'h5013;
  assign T_6660 = io_imem_resp_bits_data_0 & 32'hbe00705f;
  assign T_6662 = T_6660 == 32'h501b;
  assign T_6666 = T_6608 == 32'h5033;
  assign T_6668 = io_imem_resp_bits_data_0 & 32'hfe004077;
  assign T_6670 = T_6668 == 32'h2004033;
  assign T_6672 = io_imem_resp_bits_data_0 & 32'he800607f;
  assign T_6674 = T_6672 == 32'h800202f;
  assign T_6676 = io_imem_resp_bits_data_0 & 32'hf9f0607f;
  assign T_6678 = T_6676 == 32'h1000202f;
  assign T_6680 = io_imem_resp_bits_data_0 & 32'hdfffffff;
  assign T_6682 = T_6680 == 32'h10200073;
  assign T_6684 = io_imem_resp_bits_data_0 & 32'hfff07fff;
  assign T_6686 = T_6684 == 32'h10400073;
  assign T_6688 = io_imem_resp_bits_data_0 == 32'h10500073;
  assign T_6690 = io_imem_resp_bits_data_0 & 32'hf400607f;
  assign T_6692 = T_6690 == 32'h20000053;
  assign T_6694 = io_imem_resp_bits_data_0 & 32'h7c00607f;
  assign T_6696 = T_6694 == 32'h20000053;
  assign T_6698 = io_imem_resp_bits_data_0 & 32'h7c00507f;
  assign T_6700 = T_6698 == 32'h20000053;
  assign T_6702 = io_imem_resp_bits_data_0 & 32'h7ff0007f;
  assign T_6704 = T_6702 == 32'h40100053;
  assign T_6708 = T_6702 == 32'h42000053;
  assign T_6710 = io_imem_resp_bits_data_0 & 32'hfdf0007f;
  assign T_6712 = T_6710 == 32'h58000053;
  assign T_6714 = io_imem_resp_bits_data_0 == 32'h7b200073;
  assign T_6716 = io_imem_resp_bits_data_0 & 32'hedc0007f;
  assign T_6718 = T_6716 == 32'hc0000053;
  assign T_6720 = io_imem_resp_bits_data_0 & 32'hfdf0607f;
  assign T_6722 = T_6720 == 32'he0000053;
  assign T_6724 = io_imem_resp_bits_data_0 & 32'hedf0707f;
  assign T_6726 = T_6724 == 32'he0000053;
  assign T_6728 = io_imem_resp_bits_data_0 & 32'h603f;
  assign T_6730 = T_6728 == 32'h23;
  assign T_6732 = io_imem_resp_bits_data_0 & 32'h306f;
  assign T_6734 = T_6732 == 32'h1063;
  assign T_6736 = io_imem_resp_bits_data_0 & 32'h407f;
  assign T_6738 = T_6736 == 32'h4063;
  assign T_6740 = io_imem_resp_bits_data_0 & 32'hfc007077;
  assign T_6742 = T_6740 == 32'h33;
  assign T_6745 = T_6586 | T_6590;
  assign T_6746 = T_6745 | T_6594;
  assign T_6747 = T_6746 | T_6598;
  assign T_6748 = T_6747 | T_6602;
  assign T_6749 = T_6748 | T_6606;
  assign T_6750 = T_6749 | T_6610;
  assign T_6751 = T_6750 | T_6614;
  assign T_6752 = T_6751 | T_6618;
  assign T_6753 = T_6752 | T_6622;
  assign T_6754 = T_6753 | T_6626;
  assign T_6755 = T_6754 | T_6630;
  assign T_6756 = T_6755 | T_6634;
  assign T_6757 = T_6756 | T_6638;
  assign T_6758 = T_6757 | T_6642;
  assign T_6759 = T_6758 | T_6646;
  assign T_6760 = T_6759 | T_6650;
  assign T_6761 = T_6760 | T_6654;
  assign T_6762 = T_6761 | T_6658;
  assign T_6763 = T_6762 | T_6662;
  assign T_6764 = T_6763 | T_6666;
  assign T_6765 = T_6764 | T_6670;
  assign T_6766 = T_6765 | T_6674;
  assign T_6767 = T_6766 | T_6678;
  assign T_6768 = T_6767 | T_6682;
  assign T_6769 = T_6768 | T_6686;
  assign T_6770 = T_6769 | T_6688;
  assign T_6771 = T_6770 | T_6692;
  assign T_6772 = T_6771 | T_6696;
  assign T_6773 = T_6772 | T_6700;
  assign T_6774 = T_6773 | T_6704;
  assign T_6775 = T_6774 | T_6708;
  assign T_6776 = T_6775 | T_6712;
  assign T_6777 = T_6776 | T_6714;
  assign T_6778 = T_6777 | T_6718;
  assign T_6779 = T_6778 | T_6722;
  assign T_6780 = T_6779 | T_6726;
  assign T_6781 = T_6780 | T_6730;
  assign T_6782 = T_6781 | T_6734;
  assign T_6783 = T_6782 | T_6738;
  assign T_6784 = T_6783 | T_6742;
  assign T_6786 = io_imem_resp_bits_data_0 & 32'h5c;
  assign T_6788 = T_6786 == 32'h4;
  assign T_6790 = io_imem_resp_bits_data_0 & 32'h60;
  assign T_6792 = T_6790 == 32'h40;
  assign T_6795 = T_6788 | T_6792;
  assign T_6798 = io_imem_resp_bits_data_0 & 32'h74;
  assign T_6800 = T_6798 == 32'h60;
  assign T_6804 = io_imem_resp_bits_data_0 & 32'h68;
  assign T_6806 = T_6804 == 32'h68;
  assign T_6810 = io_imem_resp_bits_data_0 & 32'h203c;
  assign T_6812 = T_6810 == 32'h24;
  assign T_6816 = io_imem_resp_bits_data_0 & 32'h64;
  assign T_6818 = T_6816 == 32'h20;
  assign T_6820 = io_imem_resp_bits_data_0 & 32'h34;
  assign T_6822 = T_6820 == 32'h20;
  assign T_6824 = io_imem_resp_bits_data_0 & 32'h2048;
  assign T_6826 = T_6824 == 32'h2008;
  assign T_6829 = T_6818 | T_6822;
  assign T_6830 = T_6829 | T_6826;
  assign T_6832 = io_imem_resp_bits_data_0 & 32'h44;
  assign T_6834 = T_6832 == 32'h0;
  assign T_6836 = io_imem_resp_bits_data_0 & 32'h4024;
  assign T_6838 = T_6836 == 32'h20;
  assign T_6840 = io_imem_resp_bits_data_0 & 32'h38;
  assign T_6842 = T_6840 == 32'h20;
  assign T_6844 = io_imem_resp_bits_data_0 & 32'h2050;
  assign T_6846 = T_6844 == 32'h2000;
  assign T_6848 = io_imem_resp_bits_data_0 & 32'h90000034;
  assign T_6850 = T_6848 == 32'h90000010;
  assign T_6853 = T_6834 | T_6838;
  assign T_6854 = T_6853 | T_6842;
  assign T_6855 = T_6854 | T_6846;
  assign T_6856 = T_6855 | T_6850;
  assign T_6858 = io_imem_resp_bits_data_0 & 32'h58;
  assign T_6860 = T_6858 == 32'h0;
  assign T_6862 = io_imem_resp_bits_data_0 & 32'h20;
  assign T_6864 = T_6862 == 32'h0;
  assign T_6866 = io_imem_resp_bits_data_0 & 32'hc;
  assign T_6868 = T_6866 == 32'h4;
  assign T_6870 = io_imem_resp_bits_data_0 & 32'h48;
  assign T_6872 = T_6870 == 32'h48;
  assign T_6874 = io_imem_resp_bits_data_0 & 32'h4050;
  assign T_6876 = T_6874 == 32'h4050;
  assign T_6879 = T_6860 | T_6864;
  assign T_6880 = T_6879 | T_6868;
  assign T_6881 = T_6880 | T_6872;
  assign T_6882 = T_6881 | T_6876;
  assign T_6886 = T_6870 == 32'h0;
  assign T_6888 = io_imem_resp_bits_data_0 & 32'h18;
  assign T_6890 = T_6888 == 32'h0;
  assign T_6892 = io_imem_resp_bits_data_0 & 32'h4008;
  assign T_6894 = T_6892 == 32'h4000;
  assign T_6897 = T_6886 | T_6834;
  assign T_6898 = T_6897 | T_6890;
  assign T_6899 = T_6898 | T_6894;
  assign T_6900 = {T_6899,T_6882};
  assign T_6902 = io_imem_resp_bits_data_0 & 32'h4004;
  assign T_6904 = T_6902 == 32'h0;
  assign T_6906 = io_imem_resp_bits_data_0 & 32'h50;
  assign T_6908 = T_6906 == 32'h0;
  assign T_6910 = io_imem_resp_bits_data_0 & 32'h24;
  assign T_6912 = T_6910 == 32'h0;
  assign T_6915 = T_6904 | T_6908;
  assign T_6916 = T_6915 | T_6834;
  assign T_6917 = T_6916 | T_6912;
  assign T_6918 = T_6917 | T_6890;
  assign T_6922 = T_6820 == 32'h14;
  assign T_6925 = T_6922 | T_6872;
  assign T_6926 = {T_6925,T_6918};
  assign T_6930 = T_6888 == 32'h8;
  assign T_6934 = T_6832 == 32'h40;
  assign T_6937 = T_6930 | T_6934;
  assign T_6939 = io_imem_resp_bits_data_0 & 32'h14;
  assign T_6941 = T_6939 == 32'h14;
  assign T_6944 = T_6930 | T_6941;
  assign T_6946 = io_imem_resp_bits_data_0 & 32'h30;
  assign T_6948 = T_6946 == 32'h0;
  assign T_6950 = io_imem_resp_bits_data_0 & 32'h201c;
  assign T_6952 = T_6950 == 32'h4;
  assign T_6956 = T_6939 == 32'h10;
  assign T_6959 = T_6948 | T_6952;
  assign T_6960 = T_6959 | T_6956;
  assign T_6961 = {T_6944,T_6937};
  assign T_6962 = {T_6960,T_6961};
  assign T_6964 = io_imem_resp_bits_data_0 & 32'h10;
  assign T_6966 = T_6964 == 32'h0;
  assign T_6968 = io_imem_resp_bits_data_0 & 32'h8;
  assign T_6970 = T_6968 == 32'h0;
  assign T_6973 = T_6966 | T_6970;
  assign T_6975 = io_imem_resp_bits_data_0 & 32'h3054;
  assign T_6977 = T_6975 == 32'h1010;
  assign T_6979 = io_imem_resp_bits_data_0 & 32'h1058;
  assign T_6981 = T_6979 == 32'h1040;
  assign T_6983 = io_imem_resp_bits_data_0 & 32'h7044;
  assign T_6985 = T_6983 == 32'h7000;
  assign T_6988 = T_6977 | T_6981;
  assign T_6989 = T_6988 | T_6985;
  assign T_6991 = io_imem_resp_bits_data_0 & 32'h4054;
  assign T_6993 = T_6991 == 32'h40;
  assign T_6995 = io_imem_resp_bits_data_0 & 32'h2058;
  assign T_6997 = T_6995 == 32'h2040;
  assign T_7001 = T_6975 == 32'h3010;
  assign T_7003 = io_imem_resp_bits_data_0 & 32'h6054;
  assign T_7005 = T_7003 == 32'h6010;
  assign T_7007 = io_imem_resp_bits_data_0 & 32'h40003034;
  assign T_7009 = T_7007 == 32'h40000030;
  assign T_7011 = io_imem_resp_bits_data_0 & 32'h40001054;
  assign T_7013 = T_7011 == 32'h40001010;
  assign T_7016 = T_6993 | T_6997;
  assign T_7017 = T_7016 | T_7001;
  assign T_7018 = T_7017 | T_7005;
  assign T_7019 = T_7018 | T_7009;
  assign T_7020 = T_7019 | T_7013;
  assign T_7022 = io_imem_resp_bits_data_0 & 32'h2054;
  assign T_7024 = T_7022 == 32'h2010;
  assign T_7026 = io_imem_resp_bits_data_0 & 32'h40004054;
  assign T_7028 = T_7026 == 32'h4010;
  assign T_7030 = io_imem_resp_bits_data_0 & 32'h5054;
  assign T_7032 = T_7030 == 32'h4010;
  assign T_7034 = io_imem_resp_bits_data_0 & 32'h4058;
  assign T_7036 = T_7034 == 32'h4040;
  assign T_7039 = T_7024 | T_7028;
  assign T_7040 = T_7039 | T_7032;
  assign T_7041 = T_7040 | T_7036;
  assign T_7045 = T_7003 == 32'h2010;
  assign T_7047 = io_imem_resp_bits_data_0 & 32'h40003054;
  assign T_7049 = T_7047 == 32'h40001010;
  assign T_7052 = T_7045 | T_7036;
  assign T_7053 = T_7052 | T_7009;
  assign T_7054 = T_7053 | T_7049;
  assign T_7055 = {T_7020,T_6989};
  assign T_7056 = {T_7041,T_7055};
  assign T_7057 = {T_7054,T_7056};
  assign T_7059 = io_imem_resp_bits_data_0 & 32'h405f;
  assign T_7061 = T_7059 == 32'h3;
  assign T_7063 = io_imem_resp_bits_data_0 & 32'h107f;
  assign T_7065 = T_7063 == 32'h3;
  assign T_7067 = io_imem_resp_bits_data_0 & 32'h707f;
  assign T_7069 = T_7067 == 32'h100f;
  assign T_7072 = T_7061 | T_6586;
  assign T_7073 = T_7072 | T_7065;
  assign T_7074 = T_7073 | T_7069;
  assign T_7075 = T_7074 | T_6642;
  assign T_7076 = T_7075 | T_6650;
  assign T_7077 = T_7076 | T_6674;
  assign T_7078 = T_7077 | T_6678;
  assign T_7080 = io_imem_resp_bits_data_0 & 32'h2008;
  assign T_7082 = T_7080 == 32'h8;
  assign T_7084 = io_imem_resp_bits_data_0 & 32'h28;
  assign T_7086 = T_7084 == 32'h20;
  assign T_7088 = io_imem_resp_bits_data_0 & 32'h18000020;
  assign T_7090 = T_7088 == 32'h18000020;
  assign T_7092 = io_imem_resp_bits_data_0 & 32'h20000020;
  assign T_7094 = T_7092 == 32'h20000020;
  assign T_7097 = T_7082 | T_7086;
  assign T_7098 = T_7097 | T_7090;
  assign T_7099 = T_7098 | T_7094;
  assign T_7101 = io_imem_resp_bits_data_0 & 32'h10002008;
  assign T_7103 = T_7101 == 32'h10002008;
  assign T_7105 = io_imem_resp_bits_data_0 & 32'h40002008;
  assign T_7107 = T_7105 == 32'h40002008;
  assign T_7110 = T_7103 | T_7107;
  assign T_7112 = io_imem_resp_bits_data_0 & 32'h8000008;
  assign T_7114 = T_7112 == 32'h8000008;
  assign T_7116 = io_imem_resp_bits_data_0 & 32'h10000008;
  assign T_7118 = T_7116 == 32'h10000008;
  assign T_7120 = io_imem_resp_bits_data_0 & 32'h80000008;
  assign T_7122 = T_7120 == 32'h80000008;
  assign T_7125 = T_7082 | T_7114;
  assign T_7126 = T_7125 | T_7118;
  assign T_7127 = T_7126 | T_7122;
  assign T_7129 = io_imem_resp_bits_data_0 & 32'h18002008;
  assign T_7131 = T_7129 == 32'h2008;
  assign T_7135 = {T_7110,T_7099};
  assign T_7136 = {T_7127,T_7135};
  assign T_7137 = {T_7131,T_7136};
  assign T_7138 = {1'h0,T_7137};
  assign T_7140 = io_imem_resp_bits_data_0 & 32'h1000;
  assign T_7142 = T_7140 == 32'h1000;
  assign T_7146 = io_imem_resp_bits_data_0 & 32'h2000;
  assign T_7148 = T_7146 == 32'h2000;
  assign T_7152 = io_imem_resp_bits_data_0 & 32'h4000;
  assign T_7154 = T_7152 == 32'h4000;
  assign T_7157 = {T_7148,T_7142};
  assign T_7158 = {T_7154,T_7157};
  assign T_7160 = io_imem_resp_bits_data_0 & 32'h80000060;
  assign T_7162 = T_7160 == 32'h40;
  assign T_7164 = io_imem_resp_bits_data_0 & 32'h10000060;
  assign T_7166 = T_7164 == 32'h40;
  assign T_7168 = io_imem_resp_bits_data_0 & 32'h70;
  assign T_7170 = T_7168 == 32'h40;
  assign T_7173 = T_7162 | T_7166;
  assign T_7174 = T_7173 | T_7170;
  assign T_7176 = io_imem_resp_bits_data_0 & 32'h7c;
  assign T_7178 = T_7176 == 32'h24;
  assign T_7180 = io_imem_resp_bits_data_0 & 32'h40000060;
  assign T_7182 = T_7180 == 32'h40;
  assign T_7184 = io_imem_resp_bits_data_0 & 32'h90000060;
  assign T_7186 = T_7184 == 32'h10000040;
  assign T_7189 = T_7178 | T_7182;
  assign T_7190 = T_7189 | T_7170;
  assign T_7191 = T_7190 | T_7186;
  assign T_7195 = io_imem_resp_bits_data_0 & 32'h3c;
  assign T_7197 = T_7195 == 32'h4;
  assign T_7201 = T_7164 == 32'h10000040;
  assign T_7204 = T_7197 | T_7162;
  assign T_7205 = T_7204 | T_7170;
  assign T_7206 = T_7205 | T_7201;
  assign T_7208 = io_imem_resp_bits_data_0 & 32'h2000074;
  assign T_7210 = T_7208 == 32'h2000030;
  assign T_7216 = T_6816 == 32'h0;
  assign T_7220 = T_6906 == 32'h10;
  assign T_7222 = io_imem_resp_bits_data_0 & 32'h2024;
  assign T_7224 = T_7222 == 32'h24;
  assign T_7228 = T_7084 == 32'h28;
  assign T_7230 = io_imem_resp_bits_data_0 & 32'h1030;
  assign T_7232 = T_7230 == 32'h1030;
  assign T_7234 = io_imem_resp_bits_data_0 & 32'h2030;
  assign T_7236 = T_7234 == 32'h2030;
  assign T_7238 = io_imem_resp_bits_data_0 & 32'h90000010;
  assign T_7240 = T_7238 == 32'h80000010;
  assign T_7243 = T_7216 | T_7220;
  assign T_7244 = T_7243 | T_7224;
  assign T_7245 = T_7244 | T_7228;
  assign T_7246 = T_7245 | T_7232;
  assign T_7247 = T_7246 | T_7236;
  assign T_7248 = T_7247 | T_7240;
  assign T_7250 = io_imem_resp_bits_data_0 & 32'h1070;
  assign T_7252 = T_7250 == 32'h1070;
  assign T_7256 = io_imem_resp_bits_data_0 & 32'h2070;
  assign T_7258 = T_7256 == 32'h2070;
  assign T_7262 = io_imem_resp_bits_data_0 & 32'h3070;
  assign T_7264 = T_7262 == 32'h70;
  assign T_7267 = {T_7258,T_7252};
  assign T_7268 = {T_7264,T_7267};
  assign T_7270 = io_imem_resp_bits_data_0 & 32'h3058;
  assign T_7272 = T_7270 == 32'h1008;
  assign T_7278 = T_7270 == 32'h8;
  assign T_7282 = io_imem_resp_bits_data_0 & 32'h6048;
  assign T_7284 = T_7282 == 32'h2008;
  assign id_raddr3 = io_imem_resp_bits_data_0[31:27];
  assign id_raddr2 = io_imem_resp_bits_data_0[24:20];
  assign id_raddr1 = io_imem_resp_bits_data_0[19:15];
  assign id_waddr = io_imem_resp_bits_data_0[11:7];
  assign id_load_use = T_8097;
  assign T_7291_T_7301_addr = T_7300;
  assign T_7291_T_7301_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_7291_T_7301_data = T_7291[T_7291_T_7301_addr];
  `else
  assign T_7291_T_7301_data = T_7291_T_7301_addr >= 5'h1f ? $random : T_7291[T_7291_T_7301_addr];
  `endif
  assign T_7291_T_7312_addr = T_7311;
  assign T_7291_T_7312_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_7291_T_7312_data = T_7291[T_7291_T_7312_addr];
  `else
  assign T_7291_T_7312_data = T_7291_T_7312_addr >= 5'h1f ? $random : T_7291[T_7291_T_7312_addr];
  `endif
  assign T_7291_T_7961_data = rf_wdata;
  assign T_7291_T_7961_addr = T_7960;
  assign T_7291_T_7961_mask = GEN_163;
  assign T_7291_T_7961_en = GEN_163;
  assign T_7293 = GEN_166;
  assign GEN_173 = {{4'd0}, 1'h0};
  assign T_7296 = id_raddr1 == GEN_173;
  assign T_7300 = ~ id_raddr1;
  assign T_7302 = T_7291_T_7301_data;
  assign T_7304 = GEN_167;
  assign T_7311 = ~ id_raddr2;
  assign T_7313 = T_7291_T_7312_data;
  assign ctrl_killd = T_8188;
  assign csr_clk = clk;
  assign csr_reset = reset;
  assign csr_io_prci_reset = io_prci_reset;
  assign csr_io_prci_id = io_prci_id;
  assign csr_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign csr_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign csr_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign csr_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign csr_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign csr_io_rw_addr = T_8005;
  assign csr_io_rw_cmd = T_8006;
  assign csr_io_rw_wdata = wb_reg_wdata;
  assign csr_io_exception = wb_reg_xcpt;
  assign csr_io_retire = wb_valid;
  assign csr_io_uarch_counters_0 = 1'h0;
  assign csr_io_uarch_counters_1 = 1'h0;
  assign csr_io_uarch_counters_2 = 1'h0;
  assign csr_io_uarch_counters_3 = 1'h0;
  assign csr_io_uarch_counters_4 = 1'h0;
  assign csr_io_uarch_counters_5 = 1'h0;
  assign csr_io_uarch_counters_6 = 1'h0;
  assign csr_io_uarch_counters_7 = 1'h0;
  assign csr_io_uarch_counters_8 = 1'h0;
  assign csr_io_uarch_counters_9 = 1'h0;
  assign csr_io_uarch_counters_10 = 1'h0;
  assign csr_io_uarch_counters_11 = 1'h0;
  assign csr_io_uarch_counters_12 = 1'h0;
  assign csr_io_uarch_counters_13 = 1'h0;
  assign csr_io_uarch_counters_14 = 1'h0;
  assign csr_io_uarch_counters_15 = 1'h0;
  assign csr_io_cause = wb_reg_cause;
  assign csr_io_pc = wb_reg_pc;
  assign csr_io_badaddr = T_7988;
  assign csr_io_fcsr_flags_valid = io_fpu_fcsr_flags_valid;
  assign csr_io_fcsr_flags_bits = io_fpu_fcsr_flags_bits;
  assign csr_io_rocc_cmd_ready = GEN_247;
  assign csr_io_rocc_resp_valid = GEN_248;
  assign csr_io_rocc_resp_bits_rd = GEN_249;
  assign csr_io_rocc_resp_bits_data = GEN_250;
  assign csr_io_rocc_mem_req_valid = GEN_251;
  assign csr_io_rocc_mem_req_bits_addr = GEN_252;
  assign csr_io_rocc_mem_req_bits_tag = GEN_253;
  assign csr_io_rocc_mem_req_bits_cmd = GEN_254;
  assign csr_io_rocc_mem_req_bits_typ = GEN_255;
  assign csr_io_rocc_mem_req_bits_phys = GEN_256;
  assign csr_io_rocc_mem_req_bits_data = GEN_257;
  assign csr_io_rocc_mem_s1_kill = GEN_258;
  assign csr_io_rocc_mem_s1_data = GEN_259;
  assign csr_io_rocc_mem_invalidate_lr = GEN_260;
  assign csr_io_rocc_busy = GEN_261;
  assign csr_io_rocc_interrupt = io_rocc_interrupt;
  assign csr_io_rocc_autl_acquire_valid = GEN_262;
  assign csr_io_rocc_autl_acquire_bits_addr_block = GEN_263;
  assign csr_io_rocc_autl_acquire_bits_client_xact_id = GEN_264;
  assign csr_io_rocc_autl_acquire_bits_addr_beat = GEN_265;
  assign csr_io_rocc_autl_acquire_bits_is_builtin_type = GEN_266;
  assign csr_io_rocc_autl_acquire_bits_a_type = GEN_267;
  assign csr_io_rocc_autl_acquire_bits_union = GEN_268;
  assign csr_io_rocc_autl_acquire_bits_data = GEN_269;
  assign csr_io_rocc_autl_grant_ready = GEN_270;
  assign csr_io_rocc_fpu_req_valid = GEN_271;
  assign csr_io_rocc_fpu_req_bits_cmd = GEN_272;
  assign csr_io_rocc_fpu_req_bits_ldst = GEN_273;
  assign csr_io_rocc_fpu_req_bits_wen = GEN_274;
  assign csr_io_rocc_fpu_req_bits_ren1 = GEN_275;
  assign csr_io_rocc_fpu_req_bits_ren2 = GEN_276;
  assign csr_io_rocc_fpu_req_bits_ren3 = GEN_277;
  assign csr_io_rocc_fpu_req_bits_swap12 = GEN_278;
  assign csr_io_rocc_fpu_req_bits_swap23 = GEN_279;
  assign csr_io_rocc_fpu_req_bits_single = GEN_280;
  assign csr_io_rocc_fpu_req_bits_fromint = GEN_281;
  assign csr_io_rocc_fpu_req_bits_toint = GEN_282;
  assign csr_io_rocc_fpu_req_bits_fastpipe = GEN_283;
  assign csr_io_rocc_fpu_req_bits_fma = GEN_284;
  assign csr_io_rocc_fpu_req_bits_div = GEN_285;
  assign csr_io_rocc_fpu_req_bits_sqrt = GEN_286;
  assign csr_io_rocc_fpu_req_bits_round = GEN_287;
  assign csr_io_rocc_fpu_req_bits_wflags = GEN_288;
  assign csr_io_rocc_fpu_req_bits_rm = GEN_289;
  assign csr_io_rocc_fpu_req_bits_typ = GEN_290;
  assign csr_io_rocc_fpu_req_bits_in1 = GEN_291;
  assign csr_io_rocc_fpu_req_bits_in2 = GEN_292;
  assign csr_io_rocc_fpu_req_bits_in3 = GEN_293;
  assign csr_io_rocc_fpu_resp_ready = GEN_294;
  assign id_csr_en = id_ctrl_csr != 3'h0;
  assign id_system_insn = id_ctrl_csr == 3'h4;
  assign T_7315 = id_ctrl_csr == 3'h2;
  assign T_7316 = id_ctrl_csr == 3'h3;
  assign T_7317 = T_7315 | T_7316;
  assign id_csr_ren = T_7317 & T_7296;
  assign id_csr = id_csr_ren ? 3'h5 : id_ctrl_csr;
  assign id_csr_addr = io_imem_resp_bits_data_0[31:20];
  assign T_7321 = id_csr_ren == 1'h0;
  assign T_7322 = id_csr_en & T_7321;
  assign T_7377 = id_csr_addr & 12'h46;
  assign T_7379 = T_7377 == 12'h40;
  assign T_7381 = id_csr_addr & 12'h644;
  assign T_7383 = T_7381 == 12'h240;
  assign T_7386 = T_7379 | T_7383;
  assign T_7389 = T_7386 == 1'h0;
  assign T_7390 = T_7322 & T_7389;
  assign id_csr_flush = id_system_insn | T_7390;
  assign T_7392 = id_ctrl_legal == 1'h0;
  assign GEN_176 = {{1'd0}, 1'h0};
  assign T_7394 = csr_io_status_fs != GEN_176;
  assign T_7396 = T_7394 == 1'h0;
  assign T_7397 = id_ctrl_fp & T_7396;
  assign T_7398 = T_7392 | T_7397;
  assign T_7400 = csr_io_status_xs != GEN_176;
  assign T_7402 = T_7400 == 1'h0;
  assign T_7403 = id_ctrl_rocc & T_7402;
  assign id_illegal_insn = T_7398 | T_7403;
  assign id_amo_aq = io_imem_resp_bits_data_0[26];
  assign id_amo_rl = io_imem_resp_bits_data_0[25];
  assign T_7404 = id_ctrl_amo & id_amo_rl;
  assign id_fence_next = id_ctrl_fence | T_7404;
  assign T_7406 = io_dmem_ordered == 1'h0;
  assign id_mem_busy = T_7406 | io_dmem_req_valid;
  assign T_7412 = wb_reg_valid & wb_ctrl_rocc;
  assign T_7414 = id_reg_fence & id_mem_busy;
  assign T_7415 = id_fence_next | T_7414;
  assign T_7417 = id_ctrl_amo & id_amo_aq;
  assign T_7418 = T_7417 | id_ctrl_fence_i;
  assign T_7419 = id_ctrl_mem | id_ctrl_rocc;
  assign T_7420 = id_reg_fence & T_7419;
  assign T_7421 = T_7418 | T_7420;
  assign T_7422 = T_7421 | id_csr_en;
  assign T_7423 = id_mem_busy & T_7422;
  assign bpu_clk = clk;
  assign bpu_reset = reset;
  assign bpu_io_status_debug = csr_io_status_debug;
  assign bpu_io_status_prv = csr_io_status_prv;
  assign bpu_io_status_sd = csr_io_status_sd;
  assign bpu_io_status_zero3 = csr_io_status_zero3;
  assign bpu_io_status_sd_rv32 = csr_io_status_sd_rv32;
  assign bpu_io_status_zero2 = csr_io_status_zero2;
  assign bpu_io_status_vm = csr_io_status_vm;
  assign bpu_io_status_zero1 = csr_io_status_zero1;
  assign bpu_io_status_pum = csr_io_status_pum;
  assign bpu_io_status_mprv = csr_io_status_mprv;
  assign bpu_io_status_xs = csr_io_status_xs;
  assign bpu_io_status_fs = csr_io_status_fs;
  assign bpu_io_status_mpp = csr_io_status_mpp;
  assign bpu_io_status_hpp = csr_io_status_hpp;
  assign bpu_io_status_spp = csr_io_status_spp;
  assign bpu_io_status_mpie = csr_io_status_mpie;
  assign bpu_io_status_hpie = csr_io_status_hpie;
  assign bpu_io_status_spie = csr_io_status_spie;
  assign bpu_io_status_upie = csr_io_status_upie;
  assign bpu_io_status_mie = csr_io_status_mie;
  assign bpu_io_status_hie = csr_io_status_hie;
  assign bpu_io_status_sie = csr_io_status_sie;
  assign bpu_io_status_uie = csr_io_status_uie;
  assign bpu_io_bp_0_control_tdrtype = csr_io_bp_0_control_tdrtype;
  assign bpu_io_bp_0_control_bpamaskmax = csr_io_bp_0_control_bpamaskmax;
  assign bpu_io_bp_0_control_reserved = csr_io_bp_0_control_reserved;
  assign bpu_io_bp_0_control_bpaction = csr_io_bp_0_control_bpaction;
  assign bpu_io_bp_0_control_bpmatch = csr_io_bp_0_control_bpmatch;
  assign bpu_io_bp_0_control_m = csr_io_bp_0_control_m;
  assign bpu_io_bp_0_control_h = csr_io_bp_0_control_h;
  assign bpu_io_bp_0_control_s = csr_io_bp_0_control_s;
  assign bpu_io_bp_0_control_u = csr_io_bp_0_control_u;
  assign bpu_io_bp_0_control_r = csr_io_bp_0_control_r;
  assign bpu_io_bp_0_control_w = csr_io_bp_0_control_w;
  assign bpu_io_bp_0_control_x = csr_io_bp_0_control_x;
  assign bpu_io_bp_0_address = csr_io_bp_0_address;
  assign bpu_io_pc = io_imem_resp_bits_pc[38:0];
  assign bpu_io_ea = mem_reg_wdata[38:0];
  assign T_7427 = csr_io_interrupt | bpu_io_xcpt_if;
  assign T_7428 = T_7427 | io_imem_resp_bits_xcpt_if;
  assign id_xcpt = T_7428 | id_illegal_insn;
  assign T_7429 = io_imem_resp_bits_xcpt_if ? {{1'd0}, 1'h1} : 2'h2;
  assign T_7430 = bpu_io_xcpt_if ? 2'h3 : T_7429;
  assign id_cause = csr_io_interrupt ? csr_io_interrupt_cause : {{62'd0}, T_7430};
  assign ex_waddr = ex_reg_inst[11:7];
  assign mem_waddr = mem_reg_inst[11:7];
  assign wb_waddr = wb_reg_inst[11:7];
  assign T_7434 = ex_reg_valid & ex_ctrl_wxd;
  assign T_7435 = mem_reg_valid & mem_ctrl_wxd;
  assign T_7437 = mem_ctrl_mem == 1'h0;
  assign T_7438 = T_7435 & T_7437;
  assign T_7440 = GEN_173 == id_raddr1;
  assign T_7442 = ex_waddr == id_raddr1;
  assign T_7443 = T_7434 & T_7442;
  assign T_7444 = mem_waddr == id_raddr1;
  assign T_7445 = T_7438 & T_7444;
  assign T_7447 = T_7435 & T_7444;
  assign T_7448 = GEN_173 == id_raddr2;
  assign T_7450 = ex_waddr == id_raddr2;
  assign T_7451 = T_7434 & T_7450;
  assign T_7452 = mem_waddr == id_raddr2;
  assign T_7453 = T_7438 & T_7452;
  assign T_7455 = T_7435 & T_7452;
  assign bypass_mux_0 = {{63'd0}, 1'h0};
  assign bypass_mux_1 = mem_reg_wdata;
  assign bypass_mux_2 = wb_reg_wdata;
  assign bypass_mux_3 = io_dmem_resp_bits_data_word_bypass;
  assign T_7483 = {ex_reg_rs_msb_0,ex_reg_rs_lsb_0};
  assign GEN_0 = GEN_4;
  assign GEN_180 = {{1'd0}, 1'h1};
  assign GEN_2 = GEN_180 == ex_reg_rs_lsb_0 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_3 = 2'h2 == ex_reg_rs_lsb_0 ? bypass_mux_2 : GEN_2;
  assign GEN_4 = 2'h3 == ex_reg_rs_lsb_0 ? bypass_mux_3 : GEN_3;
  assign T_7484 = ex_reg_rs_bypass_0 ? GEN_0 : T_7483;
  assign T_7485 = {ex_reg_rs_msb_1,ex_reg_rs_lsb_1};
  assign GEN_1 = GEN_7;
  assign GEN_5 = GEN_180 == ex_reg_rs_lsb_1 ? bypass_mux_1 : bypass_mux_0;
  assign GEN_6 = 2'h2 == ex_reg_rs_lsb_1 ? bypass_mux_2 : GEN_5;
  assign GEN_7 = 2'h3 == ex_reg_rs_lsb_1 ? bypass_mux_3 : GEN_6;
  assign T_7486 = ex_reg_rs_bypass_1 ? GEN_1 : T_7485;
  assign T_7487 = ex_ctrl_sel_imm == 3'h5;
  assign T_7489 = ex_reg_inst[31];
  assign T_7490 = $signed(T_7489);
  assign T_7491 = T_7487 ? $signed($signed(1'h0)) : $signed(T_7490);
  assign T_7492 = ex_ctrl_sel_imm == 3'h2;
  assign T_7493 = ex_reg_inst[30:20];
  assign T_7494 = $signed(T_7493);
  assign T_7495 = T_7492 ? $signed(T_7494) : $signed({11{T_7491}});
  assign T_7496 = ex_ctrl_sel_imm != 3'h2;
  assign T_7497 = ex_ctrl_sel_imm != 3'h3;
  assign T_7498 = T_7496 & T_7497;
  assign T_7499 = ex_reg_inst[19:12];
  assign T_7500 = $signed(T_7499);
  assign T_7501 = T_7498 ? $signed({8{T_7491}}) : $signed(T_7500);
  assign T_7504 = T_7492 | T_7487;
  assign T_7506 = ex_ctrl_sel_imm == 3'h3;
  assign T_7507 = ex_reg_inst[20];
  assign T_7508 = $signed(T_7507);
  assign T_7509 = ex_ctrl_sel_imm == 3'h1;
  assign T_7510 = ex_reg_inst[7];
  assign T_7511 = $signed(T_7510);
  assign T_7512 = T_7509 ? $signed(T_7511) : $signed(T_7491);
  assign T_7513 = T_7506 ? $signed(T_7508) : $signed(T_7512);
  assign T_7514 = T_7504 ? $signed($signed(1'h0)) : $signed(T_7513);
  assign T_7519 = ex_reg_inst[30:25];
  assign T_7520 = T_7504 ? {{5'd0}, 1'h0} : T_7519;
  assign T_7523 = ex_ctrl_sel_imm == 3'h0;
  assign T_7525 = T_7523 | T_7509;
  assign T_7526 = ex_reg_inst[11:8];
  assign T_7528 = ex_reg_inst[19:16];
  assign T_7529 = ex_reg_inst[24:21];
  assign T_7530 = T_7487 ? T_7528 : T_7529;
  assign T_7531 = T_7525 ? T_7526 : T_7530;
  assign T_7532 = T_7492 ? {{3'd0}, 1'h0} : T_7531;
  assign T_7535 = ex_ctrl_sel_imm == 3'h4;
  assign T_7538 = ex_reg_inst[15];
  assign T_7541 = T_7487 ? T_7538 : 1'h0;
  assign T_7543 = T_7535 ? T_7507 : T_7541;
  assign T_7545 = T_7523 ? T_7510 : T_7543;
  assign T_7546 = {T_7520,T_7532};
  assign T_7547 = {T_7546,T_7545};
  assign T_7548 = $unsigned(T_7514);
  assign T_7549 = $unsigned(T_7501);
  assign T_7550 = {T_7549,T_7548};
  assign T_7551 = $unsigned(T_7495);
  assign T_7552 = $unsigned(T_7491);
  assign T_7553 = {T_7552,T_7551};
  assign T_7554 = {T_7553,T_7550};
  assign T_7555 = {T_7554,T_7547};
  assign ex_imm = $signed(T_7555);
  assign T_7557 = $signed(T_7484);
  assign T_7558 = $signed(ex_reg_pc);
  assign T_7559 = 2'h2 == ex_ctrl_sel_alu1;
  assign GEN_182 = $signed(1'h0);
  assign T_7560 = T_7559 ? $signed(T_7558) : $signed({40{GEN_182}});
  assign T_7561 = 2'h1 == ex_ctrl_sel_alu1;
  assign ex_op1 = T_7561 ? $signed(T_7557) : $signed({{24{T_7560[39]}},T_7560});
  assign T_7563 = $signed(T_7486);
  assign T_7565 = 2'h1 == ex_ctrl_sel_alu2;
  assign T_7566 = T_7565 ? $signed($signed(4'h4)) : $signed({4{GEN_182}});
  assign T_7567 = 2'h3 == ex_ctrl_sel_alu2;
  assign T_7568 = T_7567 ? $signed(ex_imm) : $signed({{28{T_7566[3]}},T_7566});
  assign T_7569 = 2'h2 == ex_ctrl_sel_alu2;
  assign ex_op2 = T_7569 ? $signed(T_7563) : $signed({{32{T_7568[31]}},T_7568});
  assign alu_clk = clk;
  assign alu_reset = reset;
  assign alu_io_dw = ex_ctrl_alu_dw;
  assign alu_io_fn = ex_ctrl_alu_fn;
  assign alu_io_in2 = T_7570;
  assign alu_io_in1 = T_7571;
  assign T_7570 = $unsigned(ex_op2);
  assign T_7571 = $unsigned(ex_op1);
  assign div_clk = clk;
  assign div_reset = reset;
  assign div_io_req_valid = T_7572;
  assign div_io_req_bits_fn = ex_ctrl_alu_fn;
  assign div_io_req_bits_dw = ex_ctrl_alu_dw;
  assign div_io_req_bits_in1 = T_7484;
  assign div_io_req_bits_in2 = T_7486;
  assign div_io_req_bits_tag = ex_waddr;
  assign div_io_kill = T_7905;
  assign div_io_resp_ready = GEN_149;
  assign T_7572 = ex_reg_valid & ex_ctrl_div;
  assign T_7574 = ctrl_killd == 1'h0;
  assign T_7577 = T_7574 & id_xcpt;
  assign T_7579 = take_pc_mem_wb == 1'h0;
  assign T_7580 = csr_io_interrupt & T_7579;
  assign T_7581 = T_7580 & io_imem_resp_valid;
  assign GEN_8 = id_xcpt ? id_cause : ex_reg_cause;
  assign GEN_9 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_taken : ex_reg_btb_resp_taken;
  assign GEN_10 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_mask : ex_reg_btb_resp_mask;
  assign GEN_11 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bridx : ex_reg_btb_resp_bridx;
  assign GEN_12 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_target : ex_reg_btb_resp_target;
  assign GEN_13 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_entry : ex_reg_btb_resp_entry;
  assign GEN_14 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_history : ex_reg_btb_resp_bht_history;
  assign GEN_15 = io_imem_btb_resp_valid ? io_imem_btb_resp_bits_bht_value : ex_reg_btb_resp_bht_value;
  assign T_7584 = id_ctrl_fence_i | id_csr_flush;
  assign T_7585 = T_7440 | T_7443;
  assign T_7586 = T_7585 | T_7445;
  assign T_7587 = T_7586 | T_7447;
  assign T_7592 = T_7445 ? 2'h2 : 2'h3;
  assign T_7593 = T_7443 ? {{1'd0}, 1'h1} : T_7592;
  assign T_7594 = T_7440 ? {{1'd0}, 1'h0} : T_7593;
  assign T_7596 = T_7587 == 1'h0;
  assign T_7597 = id_ctrl_rxs1 & T_7596;
  assign T_7598 = T_7293[1:0];
  assign T_7599 = T_7293[63:2];
  assign GEN_16 = T_7597 ? T_7598 : T_7594;
  assign GEN_17 = T_7597 ? T_7599 : ex_reg_rs_msb_0;
  assign T_7600 = T_7448 | T_7451;
  assign T_7601 = T_7600 | T_7453;
  assign T_7602 = T_7601 | T_7455;
  assign T_7607 = T_7453 ? 2'h2 : 2'h3;
  assign T_7608 = T_7451 ? {{1'd0}, 1'h1} : T_7607;
  assign T_7609 = T_7448 ? {{1'd0}, 1'h0} : T_7608;
  assign T_7611 = T_7602 == 1'h0;
  assign T_7612 = id_ctrl_rxs2 & T_7611;
  assign T_7613 = T_7304[1:0];
  assign T_7614 = T_7304[63:2];
  assign GEN_18 = T_7612 ? T_7613 : T_7609;
  assign GEN_19 = T_7612 ? T_7614 : ex_reg_rs_msb_1;
  assign GEN_20 = T_7574 ? id_ctrl_legal : ex_ctrl_legal;
  assign GEN_21 = T_7574 ? id_ctrl_fp : ex_ctrl_fp;
  assign GEN_22 = T_7574 ? id_ctrl_rocc : ex_ctrl_rocc;
  assign GEN_23 = T_7574 ? id_ctrl_branch : ex_ctrl_branch;
  assign GEN_24 = T_7574 ? id_ctrl_jal : ex_ctrl_jal;
  assign GEN_25 = T_7574 ? id_ctrl_jalr : ex_ctrl_jalr;
  assign GEN_26 = T_7574 ? id_ctrl_rxs2 : ex_ctrl_rxs2;
  assign GEN_27 = T_7574 ? id_ctrl_rxs1 : ex_ctrl_rxs1;
  assign GEN_28 = T_7574 ? id_ctrl_sel_alu2 : ex_ctrl_sel_alu2;
  assign GEN_29 = T_7574 ? id_ctrl_sel_alu1 : ex_ctrl_sel_alu1;
  assign GEN_30 = T_7574 ? id_ctrl_sel_imm : ex_ctrl_sel_imm;
  assign GEN_31 = T_7574 ? id_ctrl_alu_dw : ex_ctrl_alu_dw;
  assign GEN_32 = T_7574 ? id_ctrl_alu_fn : ex_ctrl_alu_fn;
  assign GEN_33 = T_7574 ? id_ctrl_mem : ex_ctrl_mem;
  assign GEN_34 = T_7574 ? id_ctrl_mem_cmd : ex_ctrl_mem_cmd;
  assign GEN_35 = T_7574 ? id_ctrl_mem_type : ex_ctrl_mem_type;
  assign GEN_36 = T_7574 ? id_ctrl_rfs1 : ex_ctrl_rfs1;
  assign GEN_37 = T_7574 ? id_ctrl_rfs2 : ex_ctrl_rfs2;
  assign GEN_38 = T_7574 ? id_ctrl_rfs3 : ex_ctrl_rfs3;
  assign GEN_39 = T_7574 ? id_ctrl_wfd : ex_ctrl_wfd;
  assign GEN_40 = T_7574 ? id_ctrl_div : ex_ctrl_div;
  assign GEN_41 = T_7574 ? id_ctrl_wxd : ex_ctrl_wxd;
  assign GEN_42 = T_7574 ? id_csr : ex_ctrl_csr;
  assign GEN_43 = T_7574 ? id_ctrl_fence_i : ex_ctrl_fence_i;
  assign GEN_44 = T_7574 ? id_ctrl_fence : ex_ctrl_fence;
  assign GEN_45 = T_7574 ? id_ctrl_amo : ex_ctrl_amo;
  assign GEN_46 = T_7574 ? io_imem_btb_resp_valid : ex_reg_btb_hit;
  assign GEN_47 = T_7574 ? GEN_9 : ex_reg_btb_resp_taken;
  assign GEN_48 = T_7574 ? GEN_10 : ex_reg_btb_resp_mask;
  assign GEN_49 = T_7574 ? GEN_11 : ex_reg_btb_resp_bridx;
  assign GEN_50 = T_7574 ? GEN_12 : ex_reg_btb_resp_target;
  assign GEN_51 = T_7574 ? GEN_13 : ex_reg_btb_resp_entry;
  assign GEN_52 = T_7574 ? GEN_14 : ex_reg_btb_resp_bht_history;
  assign GEN_53 = T_7574 ? GEN_15 : ex_reg_btb_resp_bht_value;
  assign GEN_54 = T_7574 ? T_7584 : ex_reg_flush_pipe;
  assign GEN_55 = T_7574 ? id_load_use : ex_reg_load_use;
  assign GEN_56 = T_7574 ? T_7587 : ex_reg_rs_bypass_0;
  assign GEN_57 = T_7574 ? GEN_16 : ex_reg_rs_lsb_0;
  assign GEN_58 = T_7574 ? GEN_17 : ex_reg_rs_msb_0;
  assign GEN_59 = T_7574 ? T_7602 : ex_reg_rs_bypass_1;
  assign GEN_60 = T_7574 ? GEN_18 : ex_reg_rs_lsb_1;
  assign GEN_61 = T_7574 ? GEN_19 : ex_reg_rs_msb_1;
  assign T_7617 = T_7574 | csr_io_interrupt;
  assign GEN_62 = T_7617 ? io_imem_resp_bits_data_0 : ex_reg_inst;
  assign GEN_63 = T_7617 ? io_imem_resp_bits_pc : ex_reg_pc;
  assign T_7619 = io_dmem_resp_valid == 1'h0;
  assign wb_dcache_miss = wb_ctrl_mem & T_7619;
  assign T_7621 = io_dmem_req_ready == 1'h0;
  assign T_7622 = ex_ctrl_mem & T_7621;
  assign T_7624 = div_io_req_ready == 1'h0;
  assign T_7625 = ex_ctrl_div & T_7624;
  assign replay_ex_structural = T_7622 | T_7625;
  assign replay_ex_load_use = wb_dcache_miss & ex_reg_load_use;
  assign T_7626 = replay_ex_structural | replay_ex_load_use;
  assign replay_ex = ex_reg_valid & T_7626;
  assign T_7627 = take_pc_mem_wb | replay_ex;
  assign T_7629 = ex_reg_valid == 1'h0;
  assign ctrl_killx = T_7627 | T_7629;
  assign T_7630 = ex_ctrl_mem_cmd == 5'h7;
  assign T_7636_0 = 3'h0;
  assign T_7636_1 = 3'h4;
  assign T_7636_2 = 3'h1;
  assign T_7636_3 = 3'h5;
  assign T_7638 = T_7636_0 == ex_ctrl_mem_type;
  assign T_7639 = T_7636_1 == ex_ctrl_mem_type;
  assign T_7640 = T_7636_2 == ex_ctrl_mem_type;
  assign T_7641 = T_7636_3 == ex_ctrl_mem_type;
  assign T_7644 = T_7638 | T_7639;
  assign T_7645 = T_7644 | T_7640;
  assign T_7646 = T_7645 | T_7641;
  assign ex_slow_bypass = T_7630 | T_7646;
  assign T_7647 = ex_reg_xcpt_interrupt | ex_reg_xcpt;
  assign T_7648 = ex_ctrl_fp & io_fpu_illegal_rm;
  assign ex_xcpt = T_7647 | T_7648;
  assign ex_cause = T_7647 ? ex_reg_cause : {{62'd0}, 2'h2};
  assign mem_br_taken = mem_reg_wdata[0];
  assign T_7650 = $signed(mem_reg_pc);
  assign T_7651 = mem_ctrl_branch & mem_br_taken;
  assign T_7654 = mem_reg_inst[31];
  assign T_7655 = $signed(T_7654);
  assign T_7656 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7655);
  assign T_7658 = mem_reg_inst[30:20];
  assign T_7659 = $signed(T_7658);
  assign T_7660 = 1'h0 ? $signed(T_7659) : $signed({11{T_7656}});
  assign T_7664 = mem_reg_inst[19:12];
  assign T_7665 = $signed(T_7664);
  assign T_7666 = 1'h1 ? $signed({8{T_7656}}) : $signed(T_7665);
  assign T_7672 = mem_reg_inst[20];
  assign T_7673 = $signed(T_7672);
  assign T_7675 = mem_reg_inst[7];
  assign T_7676 = $signed(T_7675);
  assign T_7677 = 1'h1 ? $signed(T_7676) : $signed(T_7656);
  assign T_7678 = 1'h0 ? $signed(T_7673) : $signed(T_7677);
  assign T_7679 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7678);
  assign T_7684 = mem_reg_inst[30:25];
  assign T_7691 = mem_reg_inst[11:8];
  assign T_7694 = mem_reg_inst[24:21];
  assign T_7711 = {T_7684,T_7691};
  assign T_7712 = {T_7711,1'h0};
  assign T_7713 = $unsigned(T_7679);
  assign T_7714 = $unsigned(T_7666);
  assign T_7715 = {T_7714,T_7713};
  assign T_7716 = $unsigned(T_7660);
  assign T_7717 = $unsigned(T_7656);
  assign T_7718 = {T_7717,T_7716};
  assign T_7719 = {T_7718,T_7715};
  assign T_7720 = {T_7719,T_7712};
  assign T_7721 = $signed(T_7720);
  assign T_7736 = 1'h0 ? $signed({8{T_7656}}) : $signed(T_7665);
  assign T_7747 = 1'h0 ? $signed(T_7676) : $signed(T_7656);
  assign T_7748 = 1'h1 ? $signed(T_7673) : $signed(T_7747);
  assign T_7749 = 1'h0 ? $signed($signed(1'h0)) : $signed(T_7748);
  assign T_7781 = {T_7684,T_7694};
  assign T_7782 = {T_7781,1'h0};
  assign T_7783 = $unsigned(T_7749);
  assign T_7784 = $unsigned(T_7736);
  assign T_7785 = {T_7784,T_7783};
  assign T_7789 = {T_7718,T_7785};
  assign T_7790 = {T_7789,T_7782};
  assign T_7791 = $signed(T_7790);
  assign GEN_184 = $signed(4'h4);
  assign T_7793 = mem_ctrl_jal ? $signed(T_7791) : $signed({{28{GEN_184[3]}},GEN_184});
  assign T_7794 = T_7651 ? $signed(T_7721) : $signed(T_7793);
  assign GEN_185 = {{8{T_7794[31]}},T_7794};
  assign T_7795 = $signed(T_7650) + $signed(GEN_185);
  assign T_7796 = T_7795[39:0];
  assign mem_br_target = $signed(T_7796);
  assign T_7797 = $signed(mem_reg_wdata);
  assign T_7798 = mem_ctrl_jalr ? $signed({{24{mem_br_target[39]}},mem_br_target}) : $signed(T_7797);
  assign mem_int_wdata = $unsigned(T_7798);
  assign T_7799 = mem_reg_wdata[63:38];
  assign T_7800 = mem_reg_wdata[39:38];
  assign T_7801 = $signed(T_7800);
  assign GEN_186 = {{25'd0}, 1'h0};
  assign T_7803 = T_7799 == GEN_186;
  assign GEN_187 = {{25'd0}, 1'h1};
  assign T_7805 = T_7799 == GEN_187;
  assign T_7806 = T_7803 | T_7805;
  assign GEN_189 = {2{GEN_182}};
  assign T_7808 = $signed(T_7801) != $signed(GEN_189);
  assign T_7809 = $signed(T_7799);
  assign GEN_190 = $signed(1'h1);
  assign GEN_191 = {26{GEN_190}};
  assign T_7811 = $signed(T_7809) == $signed(GEN_191);
  assign GEN_192 = $signed(2'h2);
  assign GEN_193 = {{24{GEN_192[1]}},GEN_192};
  assign T_7814 = $signed(T_7809) == $signed(GEN_193);
  assign T_7815 = T_7811 | T_7814;
  assign GEN_195 = {2{GEN_190}};
  assign T_7817 = $signed(T_7801) == $signed(GEN_195);
  assign T_7818 = T_7801[0];
  assign T_7819 = T_7815 ? T_7817 : T_7818;
  assign T_7820 = T_7806 ? T_7808 : T_7819;
  assign T_7821 = mem_reg_wdata[38:0];
  assign T_7822 = {T_7820,T_7821};
  assign T_7823 = $signed(T_7822);
  assign T_7824 = mem_ctrl_jalr ? $signed(T_7823) : $signed(mem_br_target);
  assign GEN_197 = {{38{GEN_192[1]}},GEN_192};
  assign T_7826 = $signed(T_7824) & $signed(GEN_197);
  assign T_7827 = $signed(T_7826);
  assign mem_npc = $unsigned(T_7827);
  assign T_7828 = mem_npc != ex_reg_pc;
  assign mem_wrong_npc = T_7828 | T_7629;
  assign mem_npc_misaligned = mem_npc[1];
  assign T_7831 = mem_ctrl_branch | mem_ctrl_jalr;
  assign mem_cfi = T_7831 | mem_ctrl_jal;
  assign T_7833 = T_7651 | mem_ctrl_jalr;
  assign mem_cfi_taken = T_7833 | mem_ctrl_jal;
  assign mem_misprediction = mem_cfi & mem_wrong_npc;
  assign T_7834 = mem_misprediction | mem_reg_flush_pipe;
  assign want_take_pc_mem = mem_reg_valid & T_7834;
  assign T_7836 = mem_npc_misaligned == 1'h0;
  assign T_7837 = want_take_pc_mem & T_7836;
  assign T_7839 = ctrl_killx == 1'h0;
  assign T_7842 = T_7579 & replay_ex;
  assign T_7845 = T_7839 & ex_xcpt;
  assign T_7848 = T_7579 & ex_reg_xcpt_interrupt;
  assign GEN_64 = ex_xcpt ? ex_cause : mem_reg_cause;
  assign T_7849 = ex_reg_valid | ex_reg_xcpt_interrupt;
  assign T_7850 = ex_ctrl_mem_cmd == 5'h0;
  assign T_7851 = ex_ctrl_mem_cmd == 5'h6;
  assign T_7852 = T_7850 | T_7851;
  assign T_7854 = T_7852 | T_7630;
  assign T_7855 = ex_ctrl_mem_cmd[3];
  assign T_7856 = ex_ctrl_mem_cmd == 5'h4;
  assign T_7857 = T_7855 | T_7856;
  assign T_7858 = T_7854 | T_7857;
  assign T_7859 = ex_ctrl_mem & T_7858;
  assign T_7860 = ex_ctrl_mem_cmd == 5'h1;
  assign T_7862 = T_7860 | T_7630;
  assign T_7866 = T_7862 | T_7857;
  assign T_7867 = ex_ctrl_mem & T_7866;
  assign GEN_65 = ex_reg_btb_hit ? ex_reg_btb_resp_taken : mem_reg_btb_resp_taken;
  assign GEN_66 = ex_reg_btb_hit ? ex_reg_btb_resp_mask : mem_reg_btb_resp_mask;
  assign GEN_67 = ex_reg_btb_hit ? ex_reg_btb_resp_bridx : mem_reg_btb_resp_bridx;
  assign GEN_68 = ex_reg_btb_hit ? ex_reg_btb_resp_target : mem_reg_btb_resp_target;
  assign GEN_69 = ex_reg_btb_hit ? ex_reg_btb_resp_entry : mem_reg_btb_resp_entry;
  assign GEN_70 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_history : mem_reg_btb_resp_bht_history;
  assign GEN_71 = ex_reg_btb_hit ? ex_reg_btb_resp_bht_value : mem_reg_btb_resp_bht_value;
  assign T_7868 = ex_ctrl_mem | ex_ctrl_rocc;
  assign T_7869 = ex_ctrl_rxs2 & T_7868;
  assign GEN_72 = T_7869 ? T_7486 : mem_reg_rs2;
  assign GEN_73 = T_7849 ? ex_ctrl_legal : mem_ctrl_legal;
  assign GEN_74 = T_7849 ? ex_ctrl_fp : mem_ctrl_fp;
  assign GEN_75 = T_7849 ? ex_ctrl_rocc : mem_ctrl_rocc;
  assign GEN_76 = T_7849 ? ex_ctrl_branch : mem_ctrl_branch;
  assign GEN_77 = T_7849 ? ex_ctrl_jal : mem_ctrl_jal;
  assign GEN_78 = T_7849 ? ex_ctrl_jalr : mem_ctrl_jalr;
  assign GEN_79 = T_7849 ? ex_ctrl_rxs2 : mem_ctrl_rxs2;
  assign GEN_80 = T_7849 ? ex_ctrl_rxs1 : mem_ctrl_rxs1;
  assign GEN_81 = T_7849 ? ex_ctrl_sel_alu2 : mem_ctrl_sel_alu2;
  assign GEN_82 = T_7849 ? ex_ctrl_sel_alu1 : mem_ctrl_sel_alu1;
  assign GEN_83 = T_7849 ? ex_ctrl_sel_imm : mem_ctrl_sel_imm;
  assign GEN_84 = T_7849 ? ex_ctrl_alu_dw : mem_ctrl_alu_dw;
  assign GEN_85 = T_7849 ? ex_ctrl_alu_fn : mem_ctrl_alu_fn;
  assign GEN_86 = T_7849 ? ex_ctrl_mem : mem_ctrl_mem;
  assign GEN_87 = T_7849 ? ex_ctrl_mem_cmd : mem_ctrl_mem_cmd;
  assign GEN_88 = T_7849 ? ex_ctrl_mem_type : mem_ctrl_mem_type;
  assign GEN_89 = T_7849 ? ex_ctrl_rfs1 : mem_ctrl_rfs1;
  assign GEN_90 = T_7849 ? ex_ctrl_rfs2 : mem_ctrl_rfs2;
  assign GEN_91 = T_7849 ? ex_ctrl_rfs3 : mem_ctrl_rfs3;
  assign GEN_92 = T_7849 ? ex_ctrl_wfd : mem_ctrl_wfd;
  assign GEN_93 = T_7849 ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_94 = T_7849 ? ex_ctrl_wxd : mem_ctrl_wxd;
  assign GEN_95 = T_7849 ? ex_ctrl_csr : mem_ctrl_csr;
  assign GEN_96 = T_7849 ? ex_ctrl_fence_i : mem_ctrl_fence_i;
  assign GEN_97 = T_7849 ? ex_ctrl_fence : mem_ctrl_fence;
  assign GEN_98 = T_7849 ? ex_ctrl_amo : mem_ctrl_amo;
  assign GEN_99 = T_7849 ? T_7859 : mem_reg_load;
  assign GEN_100 = T_7849 ? T_7867 : mem_reg_store;
  assign GEN_101 = T_7849 ? ex_reg_btb_hit : mem_reg_btb_hit;
  assign GEN_102 = T_7849 ? GEN_65 : mem_reg_btb_resp_taken;
  assign GEN_103 = T_7849 ? GEN_66 : mem_reg_btb_resp_mask;
  assign GEN_104 = T_7849 ? GEN_67 : mem_reg_btb_resp_bridx;
  assign GEN_105 = T_7849 ? GEN_68 : mem_reg_btb_resp_target;
  assign GEN_106 = T_7849 ? GEN_69 : mem_reg_btb_resp_entry;
  assign GEN_107 = T_7849 ? GEN_70 : mem_reg_btb_resp_bht_history;
  assign GEN_108 = T_7849 ? GEN_71 : mem_reg_btb_resp_bht_value;
  assign GEN_109 = T_7849 ? ex_reg_flush_pipe : mem_reg_flush_pipe;
  assign GEN_110 = T_7849 ? ex_slow_bypass : mem_reg_slow_bypass;
  assign GEN_111 = T_7849 ? ex_reg_inst : mem_reg_inst;
  assign GEN_112 = T_7849 ? ex_reg_pc : mem_reg_pc;
  assign GEN_113 = T_7849 ? alu_io_out : mem_reg_wdata;
  assign GEN_114 = T_7849 ? GEN_72 : mem_reg_rs2;
  assign T_7870 = mem_reg_load & bpu_io_xcpt_ld;
  assign T_7872 = mem_reg_store & bpu_io_xcpt_st;
  assign T_7874 = want_take_pc_mem & mem_npc_misaligned;
  assign T_7876 = mem_ctrl_mem & io_dmem_xcpt_ma_st;
  assign T_7878 = mem_ctrl_mem & io_dmem_xcpt_ma_ld;
  assign T_7880 = mem_ctrl_mem & io_dmem_xcpt_pf_st;
  assign T_7882 = mem_ctrl_mem & io_dmem_xcpt_pf_ld;
  assign T_7884 = T_7870 | T_7872;
  assign T_7885 = T_7884 | T_7874;
  assign T_7886 = T_7885 | T_7876;
  assign T_7887 = T_7886 | T_7878;
  assign T_7888 = T_7887 | T_7880;
  assign mem_new_xcpt = T_7888 | T_7882;
  assign T_7889 = T_7880 ? 3'h7 : 3'h5;
  assign T_7890 = T_7878 ? 3'h4 : T_7889;
  assign T_7891 = T_7876 ? 3'h6 : T_7890;
  assign T_7892 = T_7874 ? {{2'd0}, 1'h0} : T_7891;
  assign T_7893 = T_7872 ? {{1'd0}, 2'h3} : T_7892;
  assign mem_new_cause = T_7870 ? {{1'd0}, 2'h3} : T_7893;
  assign T_7894 = mem_reg_xcpt_interrupt | mem_reg_xcpt;
  assign T_7895 = mem_reg_valid & mem_new_xcpt;
  assign mem_xcpt = T_7894 | T_7895;
  assign mem_cause = T_7894 ? mem_reg_cause : {{61'd0}, mem_new_cause};
  assign dcache_kill_mem = T_7435 & io_dmem_replay_next;
  assign T_7897 = mem_reg_valid & mem_ctrl_fp;
  assign fpu_kill_mem = T_7897 & io_fpu_nack_mem;
  assign T_7898 = dcache_kill_mem | mem_reg_replay;
  assign replay_mem = T_7898 | fpu_kill_mem;
  assign T_7899 = dcache_kill_mem | take_pc_wb;
  assign T_7900 = T_7899 | mem_reg_xcpt;
  assign T_7902 = mem_reg_valid == 1'h0;
  assign killm_common = T_7900 | T_7902;
  assign T_7903 = div_io_req_ready & div_io_req_valid;
  assign T_7905 = killm_common & T_7904;
  assign T_7906 = killm_common | mem_xcpt;
  assign ctrl_killm = T_7906 | fpu_kill_mem;
  assign T_7908 = ctrl_killm == 1'h0;
  assign T_7910 = take_pc_wb == 1'h0;
  assign T_7911 = replay_mem & T_7910;
  assign T_7914 = mem_xcpt & T_7910;
  assign T_7918 = T_7894 == 1'h0;
  assign T_7919 = T_7895 & T_7918;
  assign GEN_115 = mem_xcpt ? mem_cause : wb_reg_cause;
  assign T_7920 = mem_reg_valid | mem_reg_replay;
  assign T_7921 = T_7920 | mem_reg_xcpt_interrupt;
  assign T_7922 = mem_ctrl_fp & mem_ctrl_wxd;
  assign T_7923 = T_7922 ? io_fpu_toint_data : mem_int_wdata;
  assign GEN_116 = mem_ctrl_rocc ? mem_reg_rs2 : wb_reg_rs2;
  assign GEN_117 = T_7921 ? mem_ctrl_legal : wb_ctrl_legal;
  assign GEN_118 = T_7921 ? mem_ctrl_fp : wb_ctrl_fp;
  assign GEN_119 = T_7921 ? mem_ctrl_rocc : wb_ctrl_rocc;
  assign GEN_120 = T_7921 ? mem_ctrl_branch : wb_ctrl_branch;
  assign GEN_121 = T_7921 ? mem_ctrl_jal : wb_ctrl_jal;
  assign GEN_122 = T_7921 ? mem_ctrl_jalr : wb_ctrl_jalr;
  assign GEN_123 = T_7921 ? mem_ctrl_rxs2 : wb_ctrl_rxs2;
  assign GEN_124 = T_7921 ? mem_ctrl_rxs1 : wb_ctrl_rxs1;
  assign GEN_125 = T_7921 ? mem_ctrl_sel_alu2 : wb_ctrl_sel_alu2;
  assign GEN_126 = T_7921 ? mem_ctrl_sel_alu1 : wb_ctrl_sel_alu1;
  assign GEN_127 = T_7921 ? mem_ctrl_sel_imm : wb_ctrl_sel_imm;
  assign GEN_128 = T_7921 ? mem_ctrl_alu_dw : wb_ctrl_alu_dw;
  assign GEN_129 = T_7921 ? mem_ctrl_alu_fn : wb_ctrl_alu_fn;
  assign GEN_130 = T_7921 ? mem_ctrl_mem : wb_ctrl_mem;
  assign GEN_131 = T_7921 ? mem_ctrl_mem_cmd : wb_ctrl_mem_cmd;
  assign GEN_132 = T_7921 ? mem_ctrl_mem_type : wb_ctrl_mem_type;
  assign GEN_133 = T_7921 ? mem_ctrl_rfs1 : wb_ctrl_rfs1;
  assign GEN_134 = T_7921 ? mem_ctrl_rfs2 : wb_ctrl_rfs2;
  assign GEN_135 = T_7921 ? mem_ctrl_rfs3 : wb_ctrl_rfs3;
  assign GEN_136 = T_7921 ? mem_ctrl_wfd : wb_ctrl_wfd;
  assign GEN_137 = T_7921 ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_138 = T_7921 ? mem_ctrl_wxd : wb_ctrl_wxd;
  assign GEN_139 = T_7921 ? mem_ctrl_csr : wb_ctrl_csr;
  assign GEN_140 = T_7921 ? mem_ctrl_fence_i : wb_ctrl_fence_i;
  assign GEN_141 = T_7921 ? mem_ctrl_fence : wb_ctrl_fence;
  assign GEN_142 = T_7921 ? mem_ctrl_amo : wb_ctrl_amo;
  assign GEN_143 = T_7921 ? T_7923 : wb_reg_wdata;
  assign GEN_144 = T_7921 ? GEN_116 : wb_reg_rs2;
  assign GEN_145 = T_7921 ? mem_reg_inst : wb_reg_inst;
  assign GEN_146 = T_7921 ? mem_reg_pc : wb_reg_pc;
  assign T_7924 = wb_ctrl_div | wb_dcache_miss;
  assign wb_set_sboard = T_7924 | wb_ctrl_rocc;
  assign replay_wb_common = io_dmem_s2_nack | wb_reg_replay;
  assign T_7927 = replay_wb_common == 1'h0;
  assign wb_rocc_val = T_7412 & T_7927;
  assign T_7930 = io_rocc_cmd_ready == 1'h0;
  assign T_7931 = T_7412 & T_7930;
  assign replay_wb = replay_wb_common | T_7931;
  assign wb_xcpt = wb_reg_xcpt | csr_io_csr_xcpt;
  assign T_7932 = replay_wb | wb_xcpt;
  assign T_7933 = T_7932 | csr_io_eret;
  assign GEN_147 = wb_rocc_val ? T_7930 : wb_reg_rocc_pending;
  assign GEN_148 = wb_reg_xcpt ? 1'h0 : GEN_147;
  assign T_7937 = io_dmem_resp_bits_tag[0];
  assign dmem_resp_xpu = T_7937 == 1'h0;
  assign dmem_resp_waddr = io_dmem_resp_bits_tag[8:1];
  assign dmem_resp_valid = io_dmem_resp_valid & io_dmem_resp_bits_has_data;
  assign dmem_resp_replay = dmem_resp_valid & io_dmem_resp_bits_replay;
  assign T_7941 = wb_reg_valid & wb_ctrl_wxd;
  assign T_7943 = T_7941 == 1'h0;
  assign ll_wdata = div_io_resp_bits_data;
  assign ll_waddr = GEN_150;
  assign T_7944 = div_io_resp_ready & div_io_resp_valid;
  assign ll_wen = GEN_151;
  assign T_7945 = dmem_resp_replay & dmem_resp_xpu;
  assign GEN_149 = T_7945 ? 1'h0 : T_7943;
  assign GEN_150 = T_7945 ? dmem_resp_waddr : {{3'd0}, div_io_resp_bits_tag};
  assign GEN_151 = T_7945 ? 1'h1 : T_7944;
  assign T_7949 = replay_wb == 1'h0;
  assign T_7950 = wb_reg_valid & T_7949;
  assign T_7952 = csr_io_csr_xcpt == 1'h0;
  assign wb_valid = T_7950 & T_7952;
  assign wb_wen = wb_valid & wb_ctrl_wxd;
  assign rf_wen = wb_wen | ll_wen;
  assign rf_waddr = ll_wen ? ll_waddr : {{3'd0}, wb_waddr};
  assign T_7953 = dmem_resp_valid & dmem_resp_xpu;
  assign T_7954 = wb_ctrl_csr != 3'h0;
  assign T_7955 = T_7954 ? csr_io_rw_rdata : wb_reg_wdata;
  assign T_7956 = ll_wen ? ll_wdata : T_7955;
  assign rf_wdata = T_7953 ? io_dmem_resp_bits_data : T_7956;
  assign GEN_198 = {{7'd0}, 1'h0};
  assign T_7958 = rf_waddr != GEN_198;
  assign T_7959 = rf_waddr[4:0];
  assign T_7960 = ~ T_7959;
  assign GEN_199 = {{3'd0}, id_raddr1};
  assign T_7962 = rf_waddr == GEN_199;
  assign GEN_152 = T_7962 ? rf_wdata : T_7302;
  assign GEN_200 = {{3'd0}, id_raddr2};
  assign T_7963 = rf_waddr == GEN_200;
  assign GEN_153 = T_7963 ? rf_wdata : T_7313;
  assign GEN_159 = T_7958 ? GEN_152 : T_7302;
  assign GEN_160 = T_7958 ? GEN_153 : T_7313;
  assign GEN_163 = rf_wen ? T_7958 : 1'h0;
  assign GEN_166 = rf_wen ? GEN_159 : T_7302;
  assign GEN_167 = rf_wen ? GEN_160 : T_7313;
  assign T_7964 = wb_reg_wdata[63:38];
  assign T_7965 = wb_reg_wdata[39:38];
  assign T_7966 = $signed(T_7965);
  assign T_7968 = T_7964 == GEN_186;
  assign T_7970 = T_7964 == GEN_187;
  assign T_7971 = T_7968 | T_7970;
  assign T_7973 = $signed(T_7966) != $signed(GEN_189);
  assign T_7974 = $signed(T_7964);
  assign T_7976 = $signed(T_7974) == $signed(GEN_191);
  assign T_7979 = $signed(T_7974) == $signed(GEN_193);
  assign T_7980 = T_7976 | T_7979;
  assign T_7982 = $signed(T_7966) == $signed(GEN_195);
  assign T_7983 = T_7966[0];
  assign T_7984 = T_7980 ? T_7982 : T_7983;
  assign T_7985 = T_7971 ? T_7973 : T_7984;
  assign T_7986 = wb_reg_wdata[38:0];
  assign T_7987 = {T_7985,T_7986};
  assign T_7988 = wb_reg_mem_xcpt ? T_7987 : wb_reg_pc;
  assign T_8005 = wb_reg_inst[31:20];
  assign T_8006 = wb_reg_valid ? wb_ctrl_csr : 3'h0;
  assign T_8008 = id_raddr1 != GEN_173;
  assign T_8009 = id_ctrl_rxs1 & T_8008;
  assign T_8011 = id_raddr2 != GEN_173;
  assign T_8012 = id_ctrl_rxs2 & T_8011;
  assign T_8014 = id_waddr != GEN_173;
  assign T_8015 = id_ctrl_wxd & T_8014;
  assign GEN_214 = {{255'd0}, 1'h1};
  assign T_8020 = GEN_214 << ll_waddr;
  assign T_8022 = ll_wen ? T_8020 : {{255'd0}, 1'h0};
  assign T_8023 = ~ T_8022;
  assign GEN_215 = {{224'd0}, T_8017};
  assign T_8024 = GEN_215 & T_8023;
  assign GEN_168 = ll_wen ? T_8024 : {{224'd0}, T_8017};
  assign T_8026 = T_8017 >> id_raddr1;
  assign T_8027 = T_8026[0];
  assign T_8028 = T_8009 & T_8027;
  assign T_8029 = T_8017 >> id_raddr2;
  assign T_8030 = T_8029[0];
  assign T_8031 = T_8012 & T_8030;
  assign T_8032 = T_8017 >> id_waddr;
  assign T_8033 = T_8032[0];
  assign T_8034 = T_8015 & T_8033;
  assign T_8035 = T_8028 | T_8031;
  assign id_sboard_hazard = T_8035 | T_8034;
  assign T_8036 = wb_set_sboard & wb_wen;
  assign GEN_216 = {{31'd0}, 1'h1};
  assign T_8038 = GEN_216 << wb_waddr;
  assign T_8040 = T_8036 ? T_8038 : {{31'd0}, 1'h0};
  assign GEN_217 = {{224'd0}, T_8040};
  assign T_8041 = T_8024 | GEN_217;
  assign T_8042 = ll_wen | T_8036;
  assign GEN_169 = T_8042 ? T_8041 : GEN_168;
  assign T_8043 = ex_ctrl_csr != 3'h0;
  assign T_8044 = T_8043 | ex_ctrl_jalr;
  assign T_8045 = T_8044 | ex_ctrl_mem;
  assign T_8046 = T_8045 | ex_ctrl_div;
  assign T_8047 = T_8046 | ex_ctrl_fp;
  assign ex_cannot_bypass = T_8047 | ex_ctrl_rocc;
  assign T_8048 = id_raddr1 == ex_waddr;
  assign T_8049 = T_8009 & T_8048;
  assign T_8050 = id_raddr2 == ex_waddr;
  assign T_8051 = T_8012 & T_8050;
  assign T_8052 = id_waddr == ex_waddr;
  assign T_8053 = T_8015 & T_8052;
  assign T_8054 = T_8049 | T_8051;
  assign T_8055 = T_8054 | T_8053;
  assign data_hazard_ex = ex_ctrl_wxd & T_8055;
  assign T_8057 = io_fpu_dec_ren1 & T_8048;
  assign T_8059 = io_fpu_dec_ren2 & T_8050;
  assign T_8060 = id_raddr3 == ex_waddr;
  assign T_8061 = io_fpu_dec_ren3 & T_8060;
  assign T_8063 = io_fpu_dec_wen & T_8052;
  assign T_8064 = T_8057 | T_8059;
  assign T_8065 = T_8064 | T_8061;
  assign T_8066 = T_8065 | T_8063;
  assign fp_data_hazard_ex = ex_ctrl_wfd & T_8066;
  assign T_8067 = data_hazard_ex & ex_cannot_bypass;
  assign T_8068 = T_8067 | fp_data_hazard_ex;
  assign id_ex_hazard = ex_reg_valid & T_8068;
  assign T_8070 = mem_ctrl_csr != 3'h0;
  assign T_8071 = mem_ctrl_mem & mem_reg_slow_bypass;
  assign T_8072 = T_8070 | T_8071;
  assign T_8073 = T_8072 | mem_ctrl_div;
  assign T_8074 = T_8073 | mem_ctrl_fp;
  assign mem_cannot_bypass = T_8074 | mem_ctrl_rocc;
  assign T_8075 = id_raddr1 == mem_waddr;
  assign T_8076 = T_8009 & T_8075;
  assign T_8077 = id_raddr2 == mem_waddr;
  assign T_8078 = T_8012 & T_8077;
  assign T_8079 = id_waddr == mem_waddr;
  assign T_8080 = T_8015 & T_8079;
  assign T_8081 = T_8076 | T_8078;
  assign T_8082 = T_8081 | T_8080;
  assign data_hazard_mem = mem_ctrl_wxd & T_8082;
  assign T_8084 = io_fpu_dec_ren1 & T_8075;
  assign T_8086 = io_fpu_dec_ren2 & T_8077;
  assign T_8087 = id_raddr3 == mem_waddr;
  assign T_8088 = io_fpu_dec_ren3 & T_8087;
  assign T_8090 = io_fpu_dec_wen & T_8079;
  assign T_8091 = T_8084 | T_8086;
  assign T_8092 = T_8091 | T_8088;
  assign T_8093 = T_8092 | T_8090;
  assign fp_data_hazard_mem = mem_ctrl_wfd & T_8093;
  assign T_8094 = data_hazard_mem & mem_cannot_bypass;
  assign T_8095 = T_8094 | fp_data_hazard_mem;
  assign id_mem_hazard = mem_reg_valid & T_8095;
  assign T_8096 = mem_reg_valid & data_hazard_mem;
  assign T_8097 = T_8096 & mem_ctrl_mem;
  assign T_8098 = id_raddr1 == wb_waddr;
  assign T_8099 = T_8009 & T_8098;
  assign T_8100 = id_raddr2 == wb_waddr;
  assign T_8101 = T_8012 & T_8100;
  assign T_8102 = id_waddr == wb_waddr;
  assign T_8103 = T_8015 & T_8102;
  assign T_8104 = T_8099 | T_8101;
  assign T_8105 = T_8104 | T_8103;
  assign data_hazard_wb = wb_ctrl_wxd & T_8105;
  assign T_8107 = io_fpu_dec_ren1 & T_8098;
  assign T_8109 = io_fpu_dec_ren2 & T_8100;
  assign T_8110 = id_raddr3 == wb_waddr;
  assign T_8111 = io_fpu_dec_ren3 & T_8110;
  assign T_8113 = io_fpu_dec_wen & T_8102;
  assign T_8114 = T_8107 | T_8109;
  assign T_8115 = T_8114 | T_8111;
  assign T_8116 = T_8115 | T_8113;
  assign fp_data_hazard_wb = wb_ctrl_wfd & T_8116;
  assign T_8117 = data_hazard_wb & wb_set_sboard;
  assign T_8118 = T_8117 | fp_data_hazard_wb;
  assign id_wb_hazard = wb_reg_valid & T_8118;
  assign T_8122 = wb_dcache_miss & wb_ctrl_wfd;
  assign T_8123 = T_8122 | io_fpu_sboard_set;
  assign T_8124 = T_8123 & wb_valid;
  assign T_8128 = T_8124 ? T_8038 : {{31'd0}, 1'h0};
  assign T_8129 = T_8120 | T_8128;
  assign GEN_170 = T_8124 ? T_8129 : T_8120;
  assign T_8131 = dmem_resp_replay & T_7937;
  assign T_8133 = GEN_214 << dmem_resp_waddr;
  assign T_8135 = T_8131 ? T_8133 : {{255'd0}, 1'h0};
  assign T_8136 = ~ T_8135;
  assign GEN_220 = {{224'd0}, T_8129};
  assign T_8137 = GEN_220 & T_8136;
  assign T_8138 = T_8124 | T_8131;
  assign GEN_171 = T_8138 ? T_8137 : {{224'd0}, GEN_170};
  assign T_8140 = GEN_216 << io_fpu_sboard_clra;
  assign T_8142 = io_fpu_sboard_clr ? T_8140 : {{31'd0}, 1'h0};
  assign T_8143 = ~ T_8142;
  assign GEN_222 = {{224'd0}, T_8143};
  assign T_8144 = T_8137 & GEN_222;
  assign T_8145 = T_8138 | io_fpu_sboard_clr;
  assign GEN_172 = T_8145 ? T_8144 : GEN_171;
  assign T_8147 = io_fpu_fcsr_rdy == 1'h0;
  assign T_8148 = id_csr_en & T_8147;
  assign T_8149 = T_8120 >> id_raddr1;
  assign T_8150 = T_8149[0];
  assign T_8151 = io_fpu_dec_ren1 & T_8150;
  assign T_8152 = T_8120 >> id_raddr2;
  assign T_8153 = T_8152[0];
  assign T_8154 = io_fpu_dec_ren2 & T_8153;
  assign T_8155 = T_8120 >> id_raddr3;
  assign T_8156 = T_8155[0];
  assign T_8157 = io_fpu_dec_ren3 & T_8156;
  assign T_8158 = T_8120 >> id_waddr;
  assign T_8159 = T_8158[0];
  assign T_8160 = io_fpu_dec_wen & T_8159;
  assign T_8161 = T_8151 | T_8154;
  assign T_8162 = T_8161 | T_8157;
  assign T_8163 = T_8162 | T_8160;
  assign id_stall_fpu = T_8148 | T_8163;
  assign T_8167 = io_dmem_req_valid | dcache_blocked;
  assign T_8168 = T_7621 & T_8167;
  assign T_8169 = id_ex_hazard | id_mem_hazard;
  assign T_8170 = T_8169 | id_wb_hazard;
  assign T_8171 = T_8170 | id_sboard_hazard;
  assign T_8172 = id_ctrl_fp & id_stall_fpu;
  assign T_8173 = T_8171 | T_8172;
  assign T_8174 = id_ctrl_mem & dcache_blocked;
  assign T_8175 = T_8173 | T_8174;
  assign T_8183 = T_8175 | T_7423;
  assign ctrl_stalld = T_8183 | csr_io_csr_stall;
  assign T_8185 = io_imem_resp_valid == 1'h0;
  assign T_8186 = T_8185 | take_pc_mem_wb;
  assign T_8187 = T_8186 | ctrl_stalld;
  assign T_8188 = T_8187 | csr_io_interrupt;
  assign T_8189 = wb_xcpt | csr_io_eret;
  assign T_8190 = replay_wb ? wb_reg_pc : mem_npc;
  assign T_8191 = T_8189 ? csr_io_evec : T_8190;
  assign T_8192 = wb_reg_valid & wb_ctrl_fence_i;
  assign T_8194 = io_dmem_s2_nack == 1'h0;
  assign T_8195 = T_8192 & T_8194;
  assign T_8197 = ctrl_stalld == 1'h0;
  assign T_8198 = T_8197 | csr_io_interrupt;
  assign T_8199 = T_8198 | take_pc_mem;
  assign T_8202 = mem_reg_valid & T_7836;
  assign T_8203 = T_8202 & mem_wrong_npc;
  assign T_8204 = T_8203 & mem_cfi_taken;
  assign T_8207 = T_8204 & T_7910;
  assign T_8208 = mem_ctrl_jal | mem_ctrl_jalr;
  assign T_8209 = mem_reg_inst[19:15];
  assign T_8212 = T_8209 & 5'h19;
  assign GEN_223 = {{4'd0}, 1'h1};
  assign T_8213 = GEN_223 == T_8212;
  assign T_8214 = mem_ctrl_jalr & T_8213;
  assign T_8215 = mem_reg_valid & mem_ctrl_branch;
  assign T_8218 = T_8215 & T_7910;
  assign T_8219 = mem_reg_valid & io_imem_btb_update_bits_isJump;
  assign T_8222 = T_8219 & T_7836;
  assign T_8225 = T_8222 & T_7910;
  assign T_8226 = mem_waddr[0];
  assign T_8227 = mem_ctrl_wxd & T_8226;
  assign T_8230 = T_7574 & id_ctrl_fp;
  assign T_8231 = dmem_resp_valid & T_7937;
  assign T_8232 = ex_reg_valid & ex_ctrl_mem;
  assign ex_dcache_tag = {ex_waddr,ex_ctrl_fp};
  assign T_8234 = T_7484[63:38];
  assign T_8235 = alu_io_adder_out[39:38];
  assign T_8236 = $signed(T_8235);
  assign T_8238 = T_8234 == GEN_186;
  assign T_8240 = T_8234 == GEN_187;
  assign T_8241 = T_8238 | T_8240;
  assign T_8243 = $signed(T_8236) != $signed(GEN_189);
  assign T_8244 = $signed(T_8234);
  assign T_8246 = $signed(T_8244) == $signed(GEN_191);
  assign T_8249 = $signed(T_8244) == $signed(GEN_193);
  assign T_8250 = T_8246 | T_8249;
  assign T_8252 = $signed(T_8236) == $signed(GEN_195);
  assign T_8253 = T_8236[0];
  assign T_8254 = T_8250 ? T_8252 : T_8253;
  assign T_8255 = T_8241 ? T_8243 : T_8254;
  assign T_8256 = alu_io_adder_out[38:0];
  assign T_8257 = {T_8255,T_8256};
  assign T_8259 = mem_ctrl_fp ? io_fpu_store_data : mem_reg_rs2;
  assign T_8262 = wb_xcpt & T_7400;
  assign T_8281_funct = T_8299;
  assign T_8281_rs2 = T_8298;
  assign T_8281_rs1 = T_8297;
  assign T_8281_xd = T_8296;
  assign T_8281_xs1 = T_8295;
  assign T_8281_xs2 = T_8294;
  assign T_8281_rd = T_8293;
  assign T_8281_opcode = T_8292;
  assign T_8291 = wb_reg_inst;
  assign T_8292 = T_8291[6:0];
  assign T_8293 = T_8291[11:7];
  assign T_8294 = T_8291[12];
  assign T_8295 = T_8291[13];
  assign T_8296 = T_8291[14];
  assign T_8297 = T_8291[19:15];
  assign T_8298 = T_8291[24:20];
  assign T_8299 = T_8291[31:25];
  assign T_8300 = csr_io_time[31:0];
  assign T_8302 = rf_wen ? rf_waddr : {{7'd0}, 1'h0};
  assign T_8303 = wb_reg_inst[19:15];
  assign T_8306 = wb_reg_inst[24:20];
  assign T_8310 = reset == 1'h0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_295 = {1{$random}};
  ex_ctrl_legal = GEN_295[0:0];
  GEN_296 = {1{$random}};
  ex_ctrl_fp = GEN_296[0:0];
  GEN_297 = {1{$random}};
  ex_ctrl_rocc = GEN_297[0:0];
  GEN_298 = {1{$random}};
  ex_ctrl_branch = GEN_298[0:0];
  GEN_299 = {1{$random}};
  ex_ctrl_jal = GEN_299[0:0];
  GEN_300 = {1{$random}};
  ex_ctrl_jalr = GEN_300[0:0];
  GEN_301 = {1{$random}};
  ex_ctrl_rxs2 = GEN_301[0:0];
  GEN_302 = {1{$random}};
  ex_ctrl_rxs1 = GEN_302[0:0];
  GEN_303 = {1{$random}};
  ex_ctrl_sel_alu2 = GEN_303[1:0];
  GEN_304 = {1{$random}};
  ex_ctrl_sel_alu1 = GEN_304[1:0];
  GEN_305 = {1{$random}};
  ex_ctrl_sel_imm = GEN_305[2:0];
  GEN_306 = {1{$random}};
  ex_ctrl_alu_dw = GEN_306[0:0];
  GEN_307 = {1{$random}};
  ex_ctrl_alu_fn = GEN_307[3:0];
  GEN_308 = {1{$random}};
  ex_ctrl_mem = GEN_308[0:0];
  GEN_309 = {1{$random}};
  ex_ctrl_mem_cmd = GEN_309[4:0];
  GEN_310 = {1{$random}};
  ex_ctrl_mem_type = GEN_310[2:0];
  GEN_311 = {1{$random}};
  ex_ctrl_rfs1 = GEN_311[0:0];
  GEN_312 = {1{$random}};
  ex_ctrl_rfs2 = GEN_312[0:0];
  GEN_313 = {1{$random}};
  ex_ctrl_rfs3 = GEN_313[0:0];
  GEN_314 = {1{$random}};
  ex_ctrl_wfd = GEN_314[0:0];
  GEN_315 = {1{$random}};
  ex_ctrl_div = GEN_315[0:0];
  GEN_316 = {1{$random}};
  ex_ctrl_wxd = GEN_316[0:0];
  GEN_317 = {1{$random}};
  ex_ctrl_csr = GEN_317[2:0];
  GEN_318 = {1{$random}};
  ex_ctrl_fence_i = GEN_318[0:0];
  GEN_319 = {1{$random}};
  ex_ctrl_fence = GEN_319[0:0];
  GEN_320 = {1{$random}};
  ex_ctrl_amo = GEN_320[0:0];
  GEN_321 = {1{$random}};
  mem_ctrl_legal = GEN_321[0:0];
  GEN_322 = {1{$random}};
  mem_ctrl_fp = GEN_322[0:0];
  GEN_323 = {1{$random}};
  mem_ctrl_rocc = GEN_323[0:0];
  GEN_324 = {1{$random}};
  mem_ctrl_branch = GEN_324[0:0];
  GEN_325 = {1{$random}};
  mem_ctrl_jal = GEN_325[0:0];
  GEN_326 = {1{$random}};
  mem_ctrl_jalr = GEN_326[0:0];
  GEN_327 = {1{$random}};
  mem_ctrl_rxs2 = GEN_327[0:0];
  GEN_328 = {1{$random}};
  mem_ctrl_rxs1 = GEN_328[0:0];
  GEN_329 = {1{$random}};
  mem_ctrl_sel_alu2 = GEN_329[1:0];
  GEN_330 = {1{$random}};
  mem_ctrl_sel_alu1 = GEN_330[1:0];
  GEN_331 = {1{$random}};
  mem_ctrl_sel_imm = GEN_331[2:0];
  GEN_332 = {1{$random}};
  mem_ctrl_alu_dw = GEN_332[0:0];
  GEN_333 = {1{$random}};
  mem_ctrl_alu_fn = GEN_333[3:0];
  GEN_334 = {1{$random}};
  mem_ctrl_mem = GEN_334[0:0];
  GEN_335 = {1{$random}};
  mem_ctrl_mem_cmd = GEN_335[4:0];
  GEN_336 = {1{$random}};
  mem_ctrl_mem_type = GEN_336[2:0];
  GEN_337 = {1{$random}};
  mem_ctrl_rfs1 = GEN_337[0:0];
  GEN_338 = {1{$random}};
  mem_ctrl_rfs2 = GEN_338[0:0];
  GEN_339 = {1{$random}};
  mem_ctrl_rfs3 = GEN_339[0:0];
  GEN_340 = {1{$random}};
  mem_ctrl_wfd = GEN_340[0:0];
  GEN_341 = {1{$random}};
  mem_ctrl_div = GEN_341[0:0];
  GEN_342 = {1{$random}};
  mem_ctrl_wxd = GEN_342[0:0];
  GEN_343 = {1{$random}};
  mem_ctrl_csr = GEN_343[2:0];
  GEN_344 = {1{$random}};
  mem_ctrl_fence_i = GEN_344[0:0];
  GEN_345 = {1{$random}};
  mem_ctrl_fence = GEN_345[0:0];
  GEN_346 = {1{$random}};
  mem_ctrl_amo = GEN_346[0:0];
  GEN_347 = {1{$random}};
  wb_ctrl_legal = GEN_347[0:0];
  GEN_348 = {1{$random}};
  wb_ctrl_fp = GEN_348[0:0];
  GEN_349 = {1{$random}};
  wb_ctrl_rocc = GEN_349[0:0];
  GEN_350 = {1{$random}};
  wb_ctrl_branch = GEN_350[0:0];
  GEN_351 = {1{$random}};
  wb_ctrl_jal = GEN_351[0:0];
  GEN_352 = {1{$random}};
  wb_ctrl_jalr = GEN_352[0:0];
  GEN_353 = {1{$random}};
  wb_ctrl_rxs2 = GEN_353[0:0];
  GEN_354 = {1{$random}};
  wb_ctrl_rxs1 = GEN_354[0:0];
  GEN_355 = {1{$random}};
  wb_ctrl_sel_alu2 = GEN_355[1:0];
  GEN_356 = {1{$random}};
  wb_ctrl_sel_alu1 = GEN_356[1:0];
  GEN_357 = {1{$random}};
  wb_ctrl_sel_imm = GEN_357[2:0];
  GEN_358 = {1{$random}};
  wb_ctrl_alu_dw = GEN_358[0:0];
  GEN_359 = {1{$random}};
  wb_ctrl_alu_fn = GEN_359[3:0];
  GEN_360 = {1{$random}};
  wb_ctrl_mem = GEN_360[0:0];
  GEN_361 = {1{$random}};
  wb_ctrl_mem_cmd = GEN_361[4:0];
  GEN_362 = {1{$random}};
  wb_ctrl_mem_type = GEN_362[2:0];
  GEN_363 = {1{$random}};
  wb_ctrl_rfs1 = GEN_363[0:0];
  GEN_364 = {1{$random}};
  wb_ctrl_rfs2 = GEN_364[0:0];
  GEN_365 = {1{$random}};
  wb_ctrl_rfs3 = GEN_365[0:0];
  GEN_366 = {1{$random}};
  wb_ctrl_wfd = GEN_366[0:0];
  GEN_367 = {1{$random}};
  wb_ctrl_div = GEN_367[0:0];
  GEN_368 = {1{$random}};
  wb_ctrl_wxd = GEN_368[0:0];
  GEN_369 = {1{$random}};
  wb_ctrl_csr = GEN_369[2:0];
  GEN_370 = {1{$random}};
  wb_ctrl_fence_i = GEN_370[0:0];
  GEN_371 = {1{$random}};
  wb_ctrl_fence = GEN_371[0:0];
  GEN_372 = {1{$random}};
  wb_ctrl_amo = GEN_372[0:0];
  GEN_373 = {1{$random}};
  ex_reg_xcpt_interrupt = GEN_373[0:0];
  GEN_374 = {1{$random}};
  ex_reg_valid = GEN_374[0:0];
  GEN_375 = {1{$random}};
  ex_reg_btb_hit = GEN_375[0:0];
  GEN_376 = {1{$random}};
  ex_reg_btb_resp_taken = GEN_376[0:0];
  GEN_377 = {1{$random}};
  ex_reg_btb_resp_mask = GEN_377[0:0];
  GEN_378 = {1{$random}};
  ex_reg_btb_resp_bridx = GEN_378[0:0];
  GEN_379 = {2{$random}};
  ex_reg_btb_resp_target = GEN_379[38:0];
  GEN_380 = {1{$random}};
  ex_reg_btb_resp_entry = GEN_380[5:0];
  GEN_381 = {1{$random}};
  ex_reg_btb_resp_bht_history = GEN_381[6:0];
  GEN_382 = {1{$random}};
  ex_reg_btb_resp_bht_value = GEN_382[1:0];
  GEN_383 = {1{$random}};
  ex_reg_xcpt = GEN_383[0:0];
  GEN_384 = {1{$random}};
  ex_reg_flush_pipe = GEN_384[0:0];
  GEN_385 = {1{$random}};
  ex_reg_load_use = GEN_385[0:0];
  GEN_386 = {2{$random}};
  ex_reg_cause = GEN_386[63:0];
  GEN_387 = {2{$random}};
  ex_reg_pc = GEN_387[39:0];
  GEN_388 = {1{$random}};
  ex_reg_inst = GEN_388[31:0];
  GEN_389 = {1{$random}};
  mem_reg_xcpt_interrupt = GEN_389[0:0];
  GEN_390 = {1{$random}};
  mem_reg_valid = GEN_390[0:0];
  GEN_391 = {1{$random}};
  mem_reg_btb_hit = GEN_391[0:0];
  GEN_392 = {1{$random}};
  mem_reg_btb_resp_taken = GEN_392[0:0];
  GEN_393 = {1{$random}};
  mem_reg_btb_resp_mask = GEN_393[0:0];
  GEN_394 = {1{$random}};
  mem_reg_btb_resp_bridx = GEN_394[0:0];
  GEN_395 = {2{$random}};
  mem_reg_btb_resp_target = GEN_395[38:0];
  GEN_396 = {1{$random}};
  mem_reg_btb_resp_entry = GEN_396[5:0];
  GEN_397 = {1{$random}};
  mem_reg_btb_resp_bht_history = GEN_397[6:0];
  GEN_398 = {1{$random}};
  mem_reg_btb_resp_bht_value = GEN_398[1:0];
  GEN_399 = {1{$random}};
  mem_reg_xcpt = GEN_399[0:0];
  GEN_400 = {1{$random}};
  mem_reg_replay = GEN_400[0:0];
  GEN_401 = {1{$random}};
  mem_reg_flush_pipe = GEN_401[0:0];
  GEN_402 = {2{$random}};
  mem_reg_cause = GEN_402[63:0];
  GEN_403 = {1{$random}};
  mem_reg_slow_bypass = GEN_403[0:0];
  GEN_404 = {1{$random}};
  mem_reg_load = GEN_404[0:0];
  GEN_405 = {1{$random}};
  mem_reg_store = GEN_405[0:0];
  GEN_406 = {2{$random}};
  mem_reg_pc = GEN_406[39:0];
  GEN_407 = {1{$random}};
  mem_reg_inst = GEN_407[31:0];
  GEN_408 = {2{$random}};
  mem_reg_wdata = GEN_408[63:0];
  GEN_409 = {2{$random}};
  mem_reg_rs2 = GEN_409[63:0];
  GEN_410 = {1{$random}};
  wb_reg_valid = GEN_410[0:0];
  GEN_411 = {1{$random}};
  wb_reg_xcpt = GEN_411[0:0];
  GEN_412 = {1{$random}};
  wb_reg_mem_xcpt = GEN_412[0:0];
  GEN_413 = {1{$random}};
  wb_reg_replay = GEN_413[0:0];
  GEN_414 = {2{$random}};
  wb_reg_cause = GEN_414[63:0];
  GEN_415 = {1{$random}};
  wb_reg_rocc_pending = GEN_415[0:0];
  GEN_416 = {2{$random}};
  wb_reg_pc = GEN_416[39:0];
  GEN_417 = {1{$random}};
  wb_reg_inst = GEN_417[31:0];
  GEN_418 = {2{$random}};
  wb_reg_wdata = GEN_418[63:0];
  GEN_419 = {2{$random}};
  wb_reg_rs2 = GEN_419[63:0];
  GEN_420 = {1{$random}};
  id_reg_fence = GEN_420[0:0];
  GEN_421 = {2{$random}};
  for (initvar = 0; initvar < 31; initvar = initvar+1)
    T_7291[initvar] = GEN_421[63:0];
  GEN_422 = {1{$random}};
  ex_reg_rs_bypass_0 = GEN_422[0:0];
  GEN_423 = {1{$random}};
  ex_reg_rs_bypass_1 = GEN_423[0:0];
  GEN_424 = {1{$random}};
  ex_reg_rs_lsb_0 = GEN_424[1:0];
  GEN_425 = {1{$random}};
  ex_reg_rs_lsb_1 = GEN_425[1:0];
  GEN_426 = {2{$random}};
  ex_reg_rs_msb_0 = GEN_426[61:0];
  GEN_427 = {2{$random}};
  ex_reg_rs_msb_1 = GEN_427[61:0];
  GEN_428 = {1{$random}};
  T_7904 = GEN_428[0:0];
  GEN_429 = {1{$random}};
  T_8017 = GEN_429[31:0];
  GEN_430 = {1{$random}};
  T_8120 = GEN_430[31:0];
  GEN_431 = {1{$random}};
  dcache_blocked = GEN_431[0:0];
  GEN_432 = {2{$random}};
  T_8304 = GEN_432[63:0];
  GEN_433 = {2{$random}};
  T_8305 = GEN_433[63:0];
  GEN_434 = {2{$random}};
  T_8307 = GEN_434[63:0];
  GEN_435 = {2{$random}};
  T_8308 = GEN_435[63:0];
  GEN_436 = {1{$random}};
  GEN_154 = GEN_436[0:0];
  GEN_437 = {2{$random}};
  GEN_155 = GEN_437[63:0];
  GEN_438 = {1{$random}};
  GEN_156 = GEN_438[0:0];
  GEN_439 = {1{$random}};
  GEN_157 = GEN_439[4:0];
  GEN_440 = {1{$random}};
  GEN_158 = GEN_440[0:0];
  GEN_441 = {1{$random}};
  GEN_161 = GEN_441[0:0];
  GEN_442 = {1{$random}};
  GEN_162 = GEN_442[0:0];
  GEN_443 = {1{$random}};
  GEN_164 = GEN_443[0:0];
  GEN_444 = {1{$random}};
  GEN_165 = GEN_444[0:0];
  GEN_445 = {1{$random}};
  GEN_174 = GEN_445[0:0];
  GEN_446 = {1{$random}};
  GEN_175 = GEN_446[0:0];
  GEN_447 = {1{$random}};
  GEN_177 = GEN_447[0:0];
  GEN_448 = {1{$random}};
  GEN_178 = GEN_448[0:0];
  GEN_449 = {1{$random}};
  GEN_179 = GEN_449[0:0];
  GEN_450 = {1{$random}};
  GEN_181 = GEN_450[0:0];
  GEN_451 = {1{$random}};
  GEN_183 = GEN_451[0:0];
  GEN_452 = {1{$random}};
  GEN_188 = GEN_452[0:0];
  GEN_453 = {1{$random}};
  GEN_194 = GEN_453[0:0];
  GEN_454 = {1{$random}};
  GEN_196 = GEN_454[0:0];
  GEN_455 = {1{$random}};
  GEN_201 = GEN_455[0:0];
  GEN_456 = {1{$random}};
  GEN_202 = GEN_456[2:0];
  GEN_457 = {1{$random}};
  GEN_203 = GEN_457[1:0];
  GEN_458 = {3{$random}};
  GEN_204 = GEN_458[64:0];
  GEN_459 = {3{$random}};
  GEN_205 = GEN_459[64:0];
  GEN_460 = {3{$random}};
  GEN_206 = GEN_460[64:0];
  GEN_461 = {1{$random}};
  GEN_207 = GEN_461[0:0];
  GEN_462 = {1{$random}};
  GEN_208 = GEN_462[0:0];
  GEN_463 = {1{$random}};
  GEN_209 = GEN_463[0:0];
  GEN_464 = {1{$random}};
  GEN_210 = GEN_464[0:0];
  GEN_465 = {1{$random}};
  GEN_211 = GEN_465[0:0];
  GEN_466 = {2{$random}};
  GEN_212 = GEN_466[39:0];
  GEN_467 = {1{$random}};
  GEN_213 = GEN_467[8:0];
  GEN_468 = {1{$random}};
  GEN_218 = GEN_468[4:0];
  GEN_469 = {1{$random}};
  GEN_219 = GEN_469[2:0];
  GEN_470 = {2{$random}};
  GEN_221 = GEN_470[63:0];
  GEN_471 = {1{$random}};
  GEN_224 = GEN_471[0:0];
  GEN_472 = {1{$random}};
  GEN_225 = GEN_472[0:0];
  GEN_473 = {2{$random}};
  GEN_226 = GEN_473[63:0];
  GEN_474 = {2{$random}};
  GEN_227 = GEN_474[63:0];
  GEN_475 = {1{$random}};
  GEN_228 = GEN_475[0:0];
  GEN_476 = {1{$random}};
  GEN_229 = GEN_476[0:0];
  GEN_477 = {1{$random}};
  GEN_230 = GEN_477[0:0];
  GEN_478 = {1{$random}};
  GEN_231 = GEN_478[0:0];
  GEN_479 = {1{$random}};
  GEN_232 = GEN_479[0:0];
  GEN_480 = {1{$random}};
  GEN_233 = GEN_480[0:0];
  GEN_481 = {1{$random}};
  GEN_234 = GEN_481[0:0];
  GEN_482 = {1{$random}};
  GEN_235 = GEN_482[0:0];
  GEN_483 = {1{$random}};
  GEN_236 = GEN_483[2:0];
  GEN_484 = {1{$random}};
  GEN_237 = GEN_484[1:0];
  GEN_485 = {1{$random}};
  GEN_238 = GEN_485[2:0];
  GEN_486 = {1{$random}};
  GEN_239 = GEN_486[0:0];
  GEN_487 = {1{$random}};
  GEN_240 = GEN_487[3:0];
  GEN_488 = {2{$random}};
  GEN_241 = GEN_488[63:0];
  GEN_489 = {1{$random}};
  GEN_242 = GEN_489[0:0];
  GEN_490 = {1{$random}};
  GEN_243 = GEN_490[0:0];
  GEN_491 = {3{$random}};
  GEN_244 = GEN_491[64:0];
  GEN_492 = {1{$random}};
  GEN_245 = GEN_492[4:0];
  GEN_493 = {1{$random}};
  GEN_246 = GEN_493[0:0];
  GEN_494 = {1{$random}};
  GEN_247 = GEN_494[0:0];
  GEN_495 = {1{$random}};
  GEN_248 = GEN_495[0:0];
  GEN_496 = {1{$random}};
  GEN_249 = GEN_496[4:0];
  GEN_497 = {2{$random}};
  GEN_250 = GEN_497[63:0];
  GEN_498 = {1{$random}};
  GEN_251 = GEN_498[0:0];
  GEN_499 = {2{$random}};
  GEN_252 = GEN_499[39:0];
  GEN_500 = {1{$random}};
  GEN_253 = GEN_500[8:0];
  GEN_501 = {1{$random}};
  GEN_254 = GEN_501[4:0];
  GEN_502 = {1{$random}};
  GEN_255 = GEN_502[2:0];
  GEN_503 = {1{$random}};
  GEN_256 = GEN_503[0:0];
  GEN_504 = {2{$random}};
  GEN_257 = GEN_504[63:0];
  GEN_505 = {1{$random}};
  GEN_258 = GEN_505[0:0];
  GEN_506 = {2{$random}};
  GEN_259 = GEN_506[63:0];
  GEN_507 = {1{$random}};
  GEN_260 = GEN_507[0:0];
  GEN_508 = {1{$random}};
  GEN_261 = GEN_508[0:0];
  GEN_509 = {1{$random}};
  GEN_262 = GEN_509[0:0];
  GEN_510 = {1{$random}};
  GEN_263 = GEN_510[25:0];
  GEN_511 = {1{$random}};
  GEN_264 = GEN_511[1:0];
  GEN_512 = {1{$random}};
  GEN_265 = GEN_512[2:0];
  GEN_513 = {1{$random}};
  GEN_266 = GEN_513[0:0];
  GEN_514 = {1{$random}};
  GEN_267 = GEN_514[2:0];
  GEN_515 = {1{$random}};
  GEN_268 = GEN_515[11:0];
  GEN_516 = {2{$random}};
  GEN_269 = GEN_516[63:0];
  GEN_517 = {1{$random}};
  GEN_270 = GEN_517[0:0];
  GEN_518 = {1{$random}};
  GEN_271 = GEN_518[0:0];
  GEN_519 = {1{$random}};
  GEN_272 = GEN_519[4:0];
  GEN_520 = {1{$random}};
  GEN_273 = GEN_520[0:0];
  GEN_521 = {1{$random}};
  GEN_274 = GEN_521[0:0];
  GEN_522 = {1{$random}};
  GEN_275 = GEN_522[0:0];
  GEN_523 = {1{$random}};
  GEN_276 = GEN_523[0:0];
  GEN_524 = {1{$random}};
  GEN_277 = GEN_524[0:0];
  GEN_525 = {1{$random}};
  GEN_278 = GEN_525[0:0];
  GEN_526 = {1{$random}};
  GEN_279 = GEN_526[0:0];
  GEN_527 = {1{$random}};
  GEN_280 = GEN_527[0:0];
  GEN_528 = {1{$random}};
  GEN_281 = GEN_528[0:0];
  GEN_529 = {1{$random}};
  GEN_282 = GEN_529[0:0];
  GEN_530 = {1{$random}};
  GEN_283 = GEN_530[0:0];
  GEN_531 = {1{$random}};
  GEN_284 = GEN_531[0:0];
  GEN_532 = {1{$random}};
  GEN_285 = GEN_532[0:0];
  GEN_533 = {1{$random}};
  GEN_286 = GEN_533[0:0];
  GEN_534 = {1{$random}};
  GEN_287 = GEN_534[0:0];
  GEN_535 = {1{$random}};
  GEN_288 = GEN_535[0:0];
  GEN_536 = {1{$random}};
  GEN_289 = GEN_536[2:0];
  GEN_537 = {1{$random}};
  GEN_290 = GEN_537[1:0];
  GEN_538 = {3{$random}};
  GEN_291 = GEN_538[64:0];
  GEN_539 = {3{$random}};
  GEN_292 = GEN_539[64:0];
  GEN_540 = {3{$random}};
  GEN_293 = GEN_540[64:0];
  GEN_541 = {1{$random}};
  GEN_294 = GEN_541[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      ex_ctrl_legal <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_fp <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rocc <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_branch <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_jal <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_jalr <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rxs2 <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rxs1 <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_sel_alu2 <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_sel_alu1 <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_sel_imm <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_alu_dw <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_alu_fn <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_mem <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_mem_cmd <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_mem_type <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rfs1 <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rfs2 <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_rfs3 <= GEN_38;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_wfd <= GEN_39;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_div <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_wxd <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_csr <= GEN_42;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_fence_i <= GEN_43;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_fence <= GEN_44;
    end
    if(1'h0) begin
    end else begin
      ex_ctrl_amo <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_legal <= GEN_73;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fp <= GEN_74;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rocc <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_branch <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_jal <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_jalr <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rxs2 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rxs1 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_sel_alu2 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_sel_alu1 <= GEN_82;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_sel_imm <= GEN_83;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_alu_dw <= GEN_84;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_alu_fn <= GEN_85;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_mem <= GEN_86;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_mem_cmd <= GEN_87;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_mem_type <= GEN_88;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rfs1 <= GEN_89;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rfs2 <= GEN_90;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_rfs3 <= GEN_91;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_wfd <= GEN_92;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_div <= GEN_93;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_wxd <= GEN_94;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_csr <= GEN_95;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fence_i <= GEN_96;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fence <= GEN_97;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_amo <= GEN_98;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_legal <= GEN_117;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fp <= GEN_118;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rocc <= GEN_119;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_branch <= GEN_120;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_jal <= GEN_121;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_jalr <= GEN_122;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rxs2 <= GEN_123;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rxs1 <= GEN_124;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_sel_alu2 <= GEN_125;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_sel_alu1 <= GEN_126;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_sel_imm <= GEN_127;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_alu_dw <= GEN_128;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_alu_fn <= GEN_129;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_mem <= GEN_130;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_mem_cmd <= GEN_131;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_mem_type <= GEN_132;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rfs1 <= GEN_133;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rfs2 <= GEN_134;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_rfs3 <= GEN_135;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_wfd <= GEN_136;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_div <= GEN_137;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_wxd <= GEN_138;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_csr <= GEN_139;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fence_i <= GEN_140;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fence <= GEN_141;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_amo <= GEN_142;
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt_interrupt <= T_7581;
    end
    if(1'h0) begin
    end else begin
      ex_reg_valid <= T_7574;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_hit <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_taken <= GEN_47;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_mask <= GEN_48;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_bridx <= GEN_49;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_target <= GEN_50;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_entry <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_bht_history <= GEN_52;
    end
    if(1'h0) begin
    end else begin
      ex_reg_btb_resp_bht_value <= GEN_53;
    end
    if(1'h0) begin
    end else begin
      ex_reg_xcpt <= T_7577;
    end
    if(1'h0) begin
    end else begin
      ex_reg_flush_pipe <= GEN_54;
    end
    if(1'h0) begin
    end else begin
      ex_reg_load_use <= GEN_55;
    end
    if(1'h0) begin
    end else begin
      ex_reg_cause <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      ex_reg_pc <= GEN_63;
    end
    if(1'h0) begin
    end else begin
      ex_reg_inst <= GEN_62;
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt_interrupt <= T_7848;
    end
    if(1'h0) begin
    end else begin
      mem_reg_valid <= T_7839;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_hit <= GEN_101;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_taken <= GEN_102;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_mask <= GEN_103;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_bridx <= GEN_104;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_target <= GEN_105;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_entry <= GEN_106;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_bht_history <= GEN_107;
    end
    if(1'h0) begin
    end else begin
      mem_reg_btb_resp_bht_value <= GEN_108;
    end
    if(1'h0) begin
    end else begin
      mem_reg_xcpt <= T_7845;
    end
    if(1'h0) begin
    end else begin
      mem_reg_replay <= T_7842;
    end
    if(1'h0) begin
    end else begin
      mem_reg_flush_pipe <= GEN_109;
    end
    if(1'h0) begin
    end else begin
      mem_reg_cause <= GEN_64;
    end
    if(1'h0) begin
    end else begin
      mem_reg_slow_bypass <= GEN_110;
    end
    if(1'h0) begin
    end else begin
      mem_reg_load <= GEN_99;
    end
    if(1'h0) begin
    end else begin
      mem_reg_store <= GEN_100;
    end
    if(1'h0) begin
    end else begin
      mem_reg_pc <= GEN_112;
    end
    if(1'h0) begin
    end else begin
      mem_reg_inst <= GEN_111;
    end
    if(1'h0) begin
    end else begin
      mem_reg_wdata <= GEN_113;
    end
    if(1'h0) begin
    end else begin
      mem_reg_rs2 <= GEN_114;
    end
    if(1'h0) begin
    end else begin
      wb_reg_valid <= T_7908;
    end
    if(1'h0) begin
    end else begin
      wb_reg_xcpt <= T_7914;
    end
    if(1'h0) begin
    end else begin
      wb_reg_mem_xcpt <= T_7919;
    end
    if(1'h0) begin
    end else begin
      wb_reg_replay <= T_7911;
    end
    if(1'h0) begin
    end else begin
      wb_reg_cause <= GEN_115;
    end
    if(reset) begin
      wb_reg_rocc_pending <= 1'h0;
    end else begin
      wb_reg_rocc_pending <= GEN_148;
    end
    if(1'h0) begin
    end else begin
      wb_reg_pc <= GEN_146;
    end
    if(1'h0) begin
    end else begin
      wb_reg_inst <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      wb_reg_wdata <= GEN_143;
    end
    if(1'h0) begin
    end else begin
      wb_reg_rs2 <= GEN_144;
    end
    if(reset) begin
      id_reg_fence <= 1'h0;
    end else begin
      id_reg_fence <= T_7415;
    end
    if(T_7291_T_7961_en & T_7291_T_7961_mask) begin
      T_7291[T_7291_T_7961_addr] <= T_7291_T_7961_data;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_bypass_0 <= GEN_56;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_bypass_1 <= GEN_59;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_lsb_0 <= GEN_57;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_lsb_1 <= GEN_60;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_msb_0 <= GEN_58;
    end
    if(1'h0) begin
    end else begin
      ex_reg_rs_msb_1 <= GEN_61;
    end
    if(1'h0) begin
    end else begin
      T_7904 <= T_7903;
    end
    if(reset) begin
      T_8017 <= 32'h0;
    end else begin
      T_8017 <= GEN_169[31:0];
    end
    if(reset) begin
      T_8120 <= 32'h0;
    end else begin
      T_8120 <= GEN_172[31:0];
    end
    if(1'h0) begin
    end else begin
      dcache_blocked <= T_8168;
    end
    if(1'h0) begin
    end else begin
      T_8304 <= T_7484;
    end
    if(1'h0) begin
    end else begin
      T_8305 <= T_8304;
    end
    if(1'h0) begin
    end else begin
      T_8307 <= T_7486;
    end
    if(1'h0) begin
    end else begin
      T_8308 <= T_8307;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_8310) begin
          $fwrite(32'h80000002,"C%d: %d [%d] pc=[%h] W[r%d=%h][%d] R[r%d=%h] R[r%d=%h] inst=[%h] DASM(%h)\n",io_prci_id,T_8300,wb_valid,wb_reg_pc,T_8302,rf_wdata,rf_wen,T_8303,T_8305,T_8306,T_8308,wb_reg_inst,wb_reg_inst);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FlowThroughSerializer(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module ICache(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  input  [19:0] io_s1_ppn,
  input   io_s1_kill,
  input   io_resp_ready,
  output  io_resp_valid,
  output [31:0] io_resp_bits_data,
  output [63:0] io_resp_bits_datablock,
  input   io_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  reg [1:0] state;
  reg [31:0] GEN_5;
  reg  invalidated;
  reg [31:0] GEN_6;
  wire  stall;
  wire  rdy;
  reg [31:0] refill_addr;
  reg [31:0] GEN_7;
  wire  s1_any_tag_hit;
  reg  s1_valid;
  reg [31:0] GEN_8;
  reg [38:0] s1_vaddr;
  reg [63:0] GEN_9;
  wire [11:0] T_934;
  wire [31:0] s1_paddr;
  wire [19:0] s1_tag;
  wire  T_935;
  wire [38:0] s0_vaddr;
  wire  T_937;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire [38:0] GEN_0;
  wire  T_946;
  wire  T_947;
  wire  out_valid;
  wire [5:0] s1_idx;
  wire  s1_hit;
  wire  T_949;
  wire  s1_miss;
  wire  T_952;
  wire  T_953;
  wire  T_955;
  wire  T_956;
  wire [31:0] GEN_1;
  wire [19:0] refill_tag;
  wire  FlowThroughSerializer_957_clk;
  wire  FlowThroughSerializer_957_reset;
  wire  FlowThroughSerializer_957_io_in_ready;
  wire  FlowThroughSerializer_957_io_in_valid;
  wire [2:0] FlowThroughSerializer_957_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_957_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_957_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_957_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_957_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_957_io_in_bits_data;
  wire  FlowThroughSerializer_957_io_out_ready;
  wire  FlowThroughSerializer_957_io_out_valid;
  wire [2:0] FlowThroughSerializer_957_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_957_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_957_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_957_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_957_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_957_io_out_bits_data;
  wire  FlowThroughSerializer_957_io_cnt;
  wire  FlowThroughSerializer_957_io_done;
  wire  T_958;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_10;
  wire  T_961;
  wire [2:0] GEN_72;
  wire [3:0] T_963;
  wire [2:0] T_964;
  wire [2:0] GEN_2;
  wire  refill_wrap;
  wire  T_965;
  wire  refill_done;
  reg [15:0] T_968;
  reg [31:0] GEN_11;
  wire  T_969;
  wire  T_970;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  wire  T_974;
  wire  T_975;
  wire [14:0] T_976;
  wire [15:0] T_977;
  wire [15:0] GEN_3;
  wire [1:0] repl_way;
  reg [19:0] tag_array_0 [0:63];
  reg [31:0] GEN_12;
  wire [19:0] tag_array_0_tag_rdata_data;
  wire [5:0] tag_array_0_tag_rdata_addr;
  wire  tag_array_0_tag_rdata_en;
  reg [5:0] GEN_13;
  reg  GEN_14;
  wire [19:0] tag_array_0_T_1019_data;
  wire [5:0] tag_array_0_T_1019_addr;
  wire  tag_array_0_T_1019_mask;
  wire  tag_array_0_T_1019_en;
  reg [19:0] tag_array_1 [0:63];
  reg [31:0] GEN_15;
  wire [19:0] tag_array_1_tag_rdata_data;
  wire [5:0] tag_array_1_tag_rdata_addr;
  wire  tag_array_1_tag_rdata_en;
  reg [5:0] GEN_16;
  reg  GEN_17;
  wire [19:0] tag_array_1_T_1019_data;
  wire [5:0] tag_array_1_T_1019_addr;
  wire  tag_array_1_T_1019_mask;
  wire  tag_array_1_T_1019_en;
  reg [19:0] tag_array_2 [0:63];
  reg [31:0] GEN_18;
  wire [19:0] tag_array_2_tag_rdata_data;
  wire [5:0] tag_array_2_tag_rdata_addr;
  wire  tag_array_2_tag_rdata_en;
  reg [5:0] GEN_19;
  reg  GEN_20;
  wire [19:0] tag_array_2_T_1019_data;
  wire [5:0] tag_array_2_T_1019_addr;
  wire  tag_array_2_T_1019_mask;
  wire  tag_array_2_T_1019_en;
  reg [19:0] tag_array_3 [0:63];
  reg [31:0] GEN_21;
  wire [19:0] tag_array_3_tag_rdata_data;
  wire [5:0] tag_array_3_tag_rdata_addr;
  wire  tag_array_3_tag_rdata_en;
  reg [5:0] GEN_22;
  reg  GEN_23;
  wire [19:0] tag_array_3_T_1019_data;
  wire [5:0] tag_array_3_T_1019_addr;
  wire  tag_array_3_T_1019_mask;
  wire  tag_array_3_T_1019_en;
  wire [5:0] T_986;
  wire [5:0] T_991;
  wire [19:0] T_1000_0;
  wire [19:0] T_1000_1;
  wire [19:0] T_1000_2;
  wire [19:0] T_1000_3;
  wire [1:0] GEN_73;
  wire  T_1003;
  wire [1:0] GEN_74;
  wire  T_1005;
  wire  T_1007;
  wire  T_1009;
  wire  T_1015_0;
  wire  T_1015_1;
  wire  T_1015_2;
  wire  T_1015_3;
  wire  GEN_25;
  wire  GEN_27;
  wire  GEN_29;
  wire  GEN_31;
  reg [255:0] vb_array;
  reg [255:0] GEN_24;
  wire  T_1023;
  wire  T_1024;
  wire [7:0] T_1025;
  wire [255:0] GEN_75;
  wire [255:0] T_1028;
  wire [255:0] T_1029;
  wire [255:0] T_1030;
  wire [255:0] GEN_32;
  wire [255:0] GEN_33;
  wire  GEN_34;
  wire  s1_disparity_0;
  wire  s1_disparity_1;
  wire  s1_disparity_2;
  wire  s1_disparity_3;
  wire  T_1043;
  wire [6:0] T_1045;
  wire [127:0] GEN_76;
  wire [127:0] T_1048;
  wire [255:0] GEN_77;
  wire [255:0] T_1051;
  wire [255:0] T_1052;
  wire [255:0] GEN_35;
  wire  T_1054;
  wire [6:0] T_1056;
  wire [127:0] T_1059;
  wire [255:0] GEN_80;
  wire [255:0] T_1062;
  wire [255:0] T_1063;
  wire [255:0] GEN_36;
  wire  T_1065;
  wire [7:0] T_1067;
  wire [255:0] T_1070;
  wire [255:0] T_1073;
  wire [255:0] T_1074;
  wire [255:0] GEN_37;
  wire  T_1076;
  wire [7:0] T_1078;
  wire [255:0] T_1081;
  wire [255:0] T_1084;
  wire [255:0] T_1085;
  wire [255:0] GEN_38;
  wire  s1_tag_match_0;
  wire  s1_tag_match_1;
  wire  s1_tag_match_2;
  wire  s1_tag_match_3;
  wire  s1_tag_hit_0;
  wire  s1_tag_hit_1;
  wire  s1_tag_hit_2;
  wire  s1_tag_hit_3;
  wire [63:0] s1_dout_0;
  wire [63:0] s1_dout_1;
  wire [63:0] s1_dout_2;
  wire [63:0] s1_dout_3;
  wire  T_1109;
  wire [255:0] T_1113;
  wire  T_1114;
  wire  T_1116;
  wire [19:0] T_1120;
  wire  T_1121;
  wire  T_1122;
  wire [255:0] T_1133;
  wire  T_1134;
  wire  T_1136;
  wire [19:0] T_1140;
  wire  T_1141;
  wire  T_1142;
  wire [255:0] T_1153;
  wire  T_1154;
  wire  T_1156;
  wire [19:0] T_1160;
  wire  T_1161;
  wire  T_1162;
  wire [255:0] T_1173;
  wire  T_1174;
  wire  T_1176;
  wire [19:0] T_1180;
  wire  T_1181;
  wire  T_1182;
  wire  T_1188;
  wire  T_1189;
  wire  T_1190;
  wire  T_1191;
  wire  T_1192;
  wire  T_1193;
  wire  T_1195;
  wire  T_1196;
  reg [63:0] T_1199 [0:511];
  reg [63:0] GEN_26;
  wire [63:0] T_1199_T_1211_data;
  wire [8:0] T_1199_T_1211_addr;
  wire  T_1199_T_1211_en;
  reg [8:0] GEN_28;
  reg  GEN_30;
  wire [63:0] T_1199_T_1204_data;
  wire [8:0] T_1199_T_1204_addr;
  wire  T_1199_T_1204_mask;
  wire  T_1199_T_1204_en;
  wire  T_1202;
  wire [8:0] T_1203;
  wire [63:0] GEN_42;
  wire [8:0] T_1205;
  wire [8:0] T_1210;
  reg [63:0] T_1214 [0:511];
  reg [63:0] GEN_39;
  wire [63:0] T_1214_T_1226_data;
  wire [8:0] T_1214_T_1226_addr;
  wire  T_1214_T_1226_en;
  reg [8:0] GEN_40;
  reg  GEN_41;
  wire [63:0] T_1214_T_1219_data;
  wire [8:0] T_1214_T_1219_addr;
  wire  T_1214_T_1219_mask;
  wire  T_1214_T_1219_en;
  wire  T_1217;
  wire [8:0] T_1225;
  reg [63:0] T_1229 [0:511];
  reg [63:0] GEN_43;
  wire [63:0] T_1229_T_1241_data;
  wire [8:0] T_1229_T_1241_addr;
  wire  T_1229_T_1241_en;
  reg [8:0] GEN_44;
  reg  GEN_45;
  wire [63:0] T_1229_T_1234_data;
  wire [8:0] T_1229_T_1234_addr;
  wire  T_1229_T_1234_mask;
  wire  T_1229_T_1234_en;
  wire  T_1232;
  wire [8:0] T_1240;
  reg [63:0] T_1244 [0:511];
  reg [63:0] GEN_46;
  wire [63:0] T_1244_T_1256_data;
  wire [8:0] T_1244_T_1256_addr;
  wire  T_1244_T_1256_en;
  reg [8:0] GEN_47;
  reg  GEN_48;
  wire [63:0] T_1244_T_1249_data;
  wire [8:0] T_1244_T_1249_addr;
  wire  T_1244_T_1249_mask;
  wire  T_1244_T_1249_en;
  wire  T_1247;
  wire [8:0] T_1255;
  wire [63:0] T_1258;
  wire [63:0] T_1260;
  wire [63:0] T_1262;
  wire [63:0] T_1264;
  wire [63:0] T_1266;
  wire [63:0] T_1267;
  wire [63:0] T_1268;
  wire [63:0] T_1269;
  wire  T_1270;
  wire [25:0] T_1271;
  wire [25:0] T_1380_addr_block;
  wire [1:0] T_1380_client_xact_id;
  wire [2:0] T_1380_addr_beat;
  wire  T_1380_is_builtin_type;
  wire [2:0] T_1380_a_type;
  wire [11:0] T_1380_union;
  wire [63:0] T_1380_data;
  wire  T_1411;
  wire [1:0] GEN_63;
  wire [1:0] GEN_64;
  wire  GEN_65;
  wire  T_1413;
  wire [1:0] GEN_66;
  wire [1:0] GEN_67;
  wire  T_1414;
  wire [1:0] GEN_68;
  wire [1:0] GEN_69;
  wire  T_1415;
  wire [1:0] GEN_70;
  wire [1:0] GEN_71;
  reg [31:0] GEN_4;
  reg [31:0] GEN_49;
  FlowThroughSerializer FlowThroughSerializer_957 (
    .clk(FlowThroughSerializer_957_clk),
    .reset(FlowThroughSerializer_957_reset),
    .io_in_ready(FlowThroughSerializer_957_io_in_ready),
    .io_in_valid(FlowThroughSerializer_957_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_957_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_957_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_957_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_957_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_957_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_957_io_in_bits_data),
    .io_out_ready(FlowThroughSerializer_957_io_out_ready),
    .io_out_valid(FlowThroughSerializer_957_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_957_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_957_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_957_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_957_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_957_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_957_io_out_bits_data),
    .io_cnt(FlowThroughSerializer_957_io_cnt),
    .io_done(FlowThroughSerializer_957_io_done)
  );
  assign io_resp_valid = s1_hit;
  assign io_resp_bits_data = GEN_4;
  assign io_resp_bits_datablock = T_1269;
  assign io_mem_acquire_valid = T_1270;
  assign io_mem_acquire_bits_addr_block = T_1380_addr_block;
  assign io_mem_acquire_bits_client_xact_id = T_1380_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = T_1380_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = T_1380_is_builtin_type;
  assign io_mem_acquire_bits_a_type = T_1380_a_type;
  assign io_mem_acquire_bits_union = T_1380_union;
  assign io_mem_acquire_bits_data = T_1380_data;
  assign io_mem_grant_ready = FlowThroughSerializer_957_io_in_ready;
  assign stall = io_resp_ready == 1'h0;
  assign rdy = T_953;
  assign s1_any_tag_hit = T_1196;
  assign T_934 = s1_vaddr[11:0];
  assign s1_paddr = {io_s1_ppn,T_934};
  assign s1_tag = s1_paddr[31:12];
  assign T_935 = s1_valid & stall;
  assign s0_vaddr = T_935 ? s1_vaddr : io_req_bits_addr;
  assign T_937 = io_req_valid & rdy;
  assign T_940 = io_s1_kill == 1'h0;
  assign T_941 = T_935 & T_940;
  assign T_942 = T_937 | T_941;
  assign GEN_0 = T_937 ? io_req_bits_addr : s1_vaddr;
  assign T_946 = s1_valid & T_940;
  assign T_947 = state == 2'h0;
  assign out_valid = T_946 & T_947;
  assign s1_idx = s1_vaddr[11:6];
  assign s1_hit = out_valid & s1_any_tag_hit;
  assign T_949 = s1_any_tag_hit == 1'h0;
  assign s1_miss = out_valid & T_949;
  assign T_952 = s1_miss == 1'h0;
  assign T_953 = T_947 & T_952;
  assign T_955 = s1_valid & T_947;
  assign T_956 = T_955 & s1_miss;
  assign GEN_1 = T_956 ? s1_paddr : refill_addr;
  assign refill_tag = refill_addr[31:12];
  assign FlowThroughSerializer_957_clk = clk;
  assign FlowThroughSerializer_957_reset = reset;
  assign FlowThroughSerializer_957_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_957_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_957_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_957_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_957_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_957_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_957_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_957_io_out_ready = 1'h1;
  assign T_958 = FlowThroughSerializer_957_io_out_ready & FlowThroughSerializer_957_io_out_valid;
  assign T_961 = refill_cnt == 3'h7;
  assign GEN_72 = {{2'd0}, 1'h1};
  assign T_963 = refill_cnt + GEN_72;
  assign T_964 = T_963[2:0];
  assign GEN_2 = T_958 ? T_964 : refill_cnt;
  assign refill_wrap = T_958 & T_961;
  assign T_965 = state == 2'h3;
  assign refill_done = T_965 & refill_wrap;
  assign T_969 = T_968[0];
  assign T_970 = T_968[2];
  assign T_971 = T_969 ^ T_970;
  assign T_972 = T_968[3];
  assign T_973 = T_971 ^ T_972;
  assign T_974 = T_968[5];
  assign T_975 = T_973 ^ T_974;
  assign T_976 = T_968[15:1];
  assign T_977 = {T_975,T_976};
  assign GEN_3 = s1_miss ? T_977 : T_968;
  assign repl_way = T_968[1:0];
  assign tag_array_0_tag_rdata_addr = T_991;
  assign tag_array_0_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_0_tag_rdata_data = tag_array_0[GEN_13];
  `else
  assign tag_array_0_tag_rdata_data = GEN_13 >= 7'h40 ? $random : tag_array_0[GEN_13];
  `endif
  assign tag_array_0_T_1019_data = T_1000_0;
  assign tag_array_0_T_1019_addr = s1_idx;
  assign tag_array_0_T_1019_mask = GEN_25;
  assign tag_array_0_T_1019_en = refill_done;
  assign tag_array_1_tag_rdata_addr = T_991;
  assign tag_array_1_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_1_tag_rdata_data = tag_array_1[GEN_16];
  `else
  assign tag_array_1_tag_rdata_data = GEN_16 >= 7'h40 ? $random : tag_array_1[GEN_16];
  `endif
  assign tag_array_1_T_1019_data = T_1000_1;
  assign tag_array_1_T_1019_addr = s1_idx;
  assign tag_array_1_T_1019_mask = GEN_27;
  assign tag_array_1_T_1019_en = refill_done;
  assign tag_array_2_tag_rdata_addr = T_991;
  assign tag_array_2_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_2_tag_rdata_data = tag_array_2[GEN_19];
  `else
  assign tag_array_2_tag_rdata_data = GEN_19 >= 7'h40 ? $random : tag_array_2[GEN_19];
  `endif
  assign tag_array_2_T_1019_data = T_1000_2;
  assign tag_array_2_T_1019_addr = s1_idx;
  assign tag_array_2_T_1019_mask = GEN_29;
  assign tag_array_2_T_1019_en = refill_done;
  assign tag_array_3_tag_rdata_addr = T_991;
  assign tag_array_3_tag_rdata_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_array_3_tag_rdata_data = tag_array_3[GEN_22];
  `else
  assign tag_array_3_tag_rdata_data = GEN_22 >= 7'h40 ? $random : tag_array_3[GEN_22];
  `endif
  assign tag_array_3_T_1019_data = T_1000_3;
  assign tag_array_3_T_1019_addr = s1_idx;
  assign tag_array_3_T_1019_mask = GEN_31;
  assign tag_array_3_T_1019_en = refill_done;
  assign T_986 = s0_vaddr[11:6];
  assign T_991 = T_986;
  assign T_1000_0 = refill_tag;
  assign T_1000_1 = refill_tag;
  assign T_1000_2 = refill_tag;
  assign T_1000_3 = refill_tag;
  assign GEN_73 = {{1'd0}, 1'h0};
  assign T_1003 = repl_way == GEN_73;
  assign GEN_74 = {{1'd0}, 1'h1};
  assign T_1005 = repl_way == GEN_74;
  assign T_1007 = repl_way == 2'h2;
  assign T_1009 = repl_way == 2'h3;
  assign T_1015_0 = T_1003;
  assign T_1015_1 = T_1005;
  assign T_1015_2 = T_1007;
  assign T_1015_3 = T_1009;
  assign GEN_25 = refill_done ? T_1015_0 : 1'h0;
  assign GEN_27 = refill_done ? T_1015_1 : 1'h0;
  assign GEN_29 = refill_done ? T_1015_2 : 1'h0;
  assign GEN_31 = refill_done ? T_1015_3 : 1'h0;
  assign T_1023 = invalidated == 1'h0;
  assign T_1024 = refill_done & T_1023;
  assign T_1025 = {repl_way,s1_idx};
  assign GEN_75 = {{255'd0}, 1'h1};
  assign T_1028 = GEN_75 << T_1025;
  assign T_1029 = vb_array | T_1028;
  assign T_1030 = ~ vb_array;
  assign GEN_32 = T_1024 ? T_1029 : vb_array;
  assign GEN_33 = io_invalidate ? {{255'd0}, 1'h0} : GEN_32;
  assign GEN_34 = io_invalidate ? 1'h1 : invalidated;
  assign s1_disparity_0 = 1'h0;
  assign s1_disparity_1 = 1'h0;
  assign s1_disparity_2 = 1'h0;
  assign s1_disparity_3 = 1'h0;
  assign T_1043 = s1_valid & s1_disparity_0;
  assign T_1045 = {1'h0,s1_idx};
  assign GEN_76 = {{127'd0}, 1'h1};
  assign T_1048 = GEN_76 << T_1045;
  assign GEN_77 = {{128'd0}, T_1048};
  assign T_1051 = T_1030 | GEN_77;
  assign T_1052 = ~ T_1051;
  assign GEN_35 = T_1043 ? T_1052 : GEN_33;
  assign T_1054 = s1_valid & s1_disparity_1;
  assign T_1056 = {1'h1,s1_idx};
  assign T_1059 = GEN_76 << T_1056;
  assign GEN_80 = {{128'd0}, T_1059};
  assign T_1062 = T_1030 | GEN_80;
  assign T_1063 = ~ T_1062;
  assign GEN_36 = T_1054 ? T_1063 : GEN_35;
  assign T_1065 = s1_valid & s1_disparity_2;
  assign T_1067 = {2'h2,s1_idx};
  assign T_1070 = GEN_75 << T_1067;
  assign T_1073 = T_1030 | T_1070;
  assign T_1074 = ~ T_1073;
  assign GEN_37 = T_1065 ? T_1074 : GEN_36;
  assign T_1076 = s1_valid & s1_disparity_3;
  assign T_1078 = {2'h3,s1_idx};
  assign T_1081 = GEN_75 << T_1078;
  assign T_1084 = T_1030 | T_1081;
  assign T_1085 = ~ T_1084;
  assign GEN_38 = T_1076 ? T_1085 : GEN_37;
  assign s1_tag_match_0 = T_1121;
  assign s1_tag_match_1 = T_1141;
  assign s1_tag_match_2 = T_1161;
  assign s1_tag_match_3 = T_1181;
  assign s1_tag_hit_0 = T_1122;
  assign s1_tag_hit_1 = T_1142;
  assign s1_tag_hit_2 = T_1162;
  assign s1_tag_hit_3 = T_1182;
  assign s1_dout_0 = T_1199_T_1211_data;
  assign s1_dout_1 = T_1214_T_1226_data;
  assign s1_dout_2 = T_1229_T_1241_data;
  assign s1_dout_3 = T_1244_T_1256_data;
  assign T_1109 = io_invalidate == 1'h0;
  assign T_1113 = vb_array >> T_1045;
  assign T_1114 = T_1113[0];
  assign T_1116 = T_1109 & T_1114;
  assign T_1120 = tag_array_0_tag_rdata_data;
  assign T_1121 = T_1120 == s1_tag;
  assign T_1122 = T_1116 & s1_tag_match_0;
  assign T_1133 = vb_array >> T_1056;
  assign T_1134 = T_1133[0];
  assign T_1136 = T_1109 & T_1134;
  assign T_1140 = tag_array_1_tag_rdata_data;
  assign T_1141 = T_1140 == s1_tag;
  assign T_1142 = T_1136 & s1_tag_match_1;
  assign T_1153 = vb_array >> T_1067;
  assign T_1154 = T_1153[0];
  assign T_1156 = T_1109 & T_1154;
  assign T_1160 = tag_array_2_tag_rdata_data;
  assign T_1161 = T_1160 == s1_tag;
  assign T_1162 = T_1156 & s1_tag_match_2;
  assign T_1173 = vb_array >> T_1078;
  assign T_1174 = T_1173[0];
  assign T_1176 = T_1109 & T_1174;
  assign T_1180 = tag_array_3_tag_rdata_data;
  assign T_1181 = T_1180 == s1_tag;
  assign T_1182 = T_1176 & s1_tag_match_3;
  assign T_1188 = s1_tag_hit_0 | s1_tag_hit_1;
  assign T_1189 = T_1188 | s1_tag_hit_2;
  assign T_1190 = T_1189 | s1_tag_hit_3;
  assign T_1191 = s1_disparity_0 | s1_disparity_1;
  assign T_1192 = T_1191 | s1_disparity_2;
  assign T_1193 = T_1192 | s1_disparity_3;
  assign T_1195 = T_1193 == 1'h0;
  assign T_1196 = T_1190 & T_1195;
  assign T_1199_T_1211_addr = T_1210;
  assign T_1199_T_1211_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1199_T_1211_data = T_1199[GEN_28];
  `else
  assign T_1199_T_1211_data = GEN_28 >= 10'h200 ? $random : T_1199[GEN_28];
  `endif
  assign T_1199_T_1204_data = GEN_42;
  assign T_1199_T_1204_addr = T_1203;
  assign T_1199_T_1204_mask = T_1202;
  assign T_1199_T_1204_en = T_1202;
  assign T_1202 = FlowThroughSerializer_957_io_out_valid & T_1003;
  assign T_1203 = {s1_idx,refill_cnt};
  assign GEN_42 = FlowThroughSerializer_957_io_out_bits_data;
  assign T_1205 = s0_vaddr[11:3];
  assign T_1210 = T_1205;
  assign T_1214_T_1226_addr = T_1225;
  assign T_1214_T_1226_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1214_T_1226_data = T_1214[GEN_40];
  `else
  assign T_1214_T_1226_data = GEN_40 >= 10'h200 ? $random : T_1214[GEN_40];
  `endif
  assign T_1214_T_1219_data = GEN_42;
  assign T_1214_T_1219_addr = T_1203;
  assign T_1214_T_1219_mask = T_1217;
  assign T_1214_T_1219_en = T_1217;
  assign T_1217 = FlowThroughSerializer_957_io_out_valid & T_1005;
  assign T_1225 = T_1205;
  assign T_1229_T_1241_addr = T_1240;
  assign T_1229_T_1241_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1229_T_1241_data = T_1229[GEN_44];
  `else
  assign T_1229_T_1241_data = GEN_44 >= 10'h200 ? $random : T_1229[GEN_44];
  `endif
  assign T_1229_T_1234_data = GEN_42;
  assign T_1229_T_1234_addr = T_1203;
  assign T_1229_T_1234_mask = T_1232;
  assign T_1229_T_1234_en = T_1232;
  assign T_1232 = FlowThroughSerializer_957_io_out_valid & T_1007;
  assign T_1240 = T_1205;
  assign T_1244_T_1256_addr = T_1255;
  assign T_1244_T_1256_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1244_T_1256_data = T_1244[GEN_47];
  `else
  assign T_1244_T_1256_data = GEN_47 >= 10'h200 ? $random : T_1244[GEN_47];
  `endif
  assign T_1244_T_1249_data = GEN_42;
  assign T_1244_T_1249_addr = T_1203;
  assign T_1244_T_1249_mask = T_1247;
  assign T_1244_T_1249_en = T_1247;
  assign T_1247 = FlowThroughSerializer_957_io_out_valid & T_1009;
  assign T_1255 = T_1205;
  assign T_1258 = s1_tag_hit_0 ? s1_dout_0 : {{63'd0}, 1'h0};
  assign T_1260 = s1_tag_hit_1 ? s1_dout_1 : {{63'd0}, 1'h0};
  assign T_1262 = s1_tag_hit_2 ? s1_dout_2 : {{63'd0}, 1'h0};
  assign T_1264 = s1_tag_hit_3 ? s1_dout_3 : {{63'd0}, 1'h0};
  assign T_1266 = T_1258 | T_1260;
  assign T_1267 = T_1266 | T_1262;
  assign T_1268 = T_1267 | T_1264;
  assign T_1269 = T_1268;
  assign T_1270 = state == 2'h1;
  assign T_1271 = refill_addr[31:6];
  assign T_1380_addr_block = T_1271;
  assign T_1380_client_xact_id = {{1'd0}, 1'h0};
  assign T_1380_addr_beat = {{2'd0}, 1'h0};
  assign T_1380_is_builtin_type = 1'h1;
  assign T_1380_a_type = 3'h1;
  assign T_1380_union = 12'h1c1;
  assign T_1380_data = {{63'd0}, 1'h0};
  assign T_1411 = 2'h0 == state;
  assign GEN_63 = s1_miss ? 2'h1 : state;
  assign GEN_64 = T_1411 ? GEN_63 : state;
  assign GEN_65 = T_1411 ? 1'h0 : GEN_34;
  assign T_1413 = 2'h1 == state;
  assign GEN_66 = io_mem_acquire_ready ? 2'h2 : GEN_64;
  assign GEN_67 = T_1413 ? GEN_66 : GEN_64;
  assign T_1414 = 2'h2 == state;
  assign GEN_68 = io_mem_grant_valid ? 2'h3 : GEN_67;
  assign GEN_69 = T_1414 ? GEN_68 : GEN_67;
  assign T_1415 = 2'h3 == state;
  assign GEN_70 = refill_done ? 2'h0 : GEN_69;
  assign GEN_71 = T_1415 ? GEN_70 : GEN_69;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_5 = {1{$random}};
  state = GEN_5[1:0];
  GEN_6 = {1{$random}};
  invalidated = GEN_6[0:0];
  GEN_7 = {1{$random}};
  refill_addr = GEN_7[31:0];
  GEN_8 = {1{$random}};
  s1_valid = GEN_8[0:0];
  GEN_9 = {2{$random}};
  s1_vaddr = GEN_9[38:0];
  GEN_10 = {1{$random}};
  refill_cnt = GEN_10[2:0];
  GEN_11 = {1{$random}};
  T_968 = GEN_11[15:0];
  GEN_12 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_0[initvar] = GEN_12[19:0];
  GEN_15 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_1[initvar] = GEN_15[19:0];
  GEN_18 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_2[initvar] = GEN_18[19:0];
  GEN_21 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_array_3[initvar] = GEN_21[19:0];
  GEN_24 = {8{$random}};
  vb_array = GEN_24[255:0];
  GEN_26 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1199[initvar] = GEN_26[63:0];
  GEN_39 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1214[initvar] = GEN_39[63:0];
  GEN_43 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1229[initvar] = GEN_43[63:0];
  GEN_46 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_1244[initvar] = GEN_46[63:0];
  GEN_49 = {1{$random}};
  GEN_4 = GEN_49[31:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 2'h0;
    end else begin
      state <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      invalidated <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      refill_addr <= GEN_1;
    end
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_942;
    end
    if(1'h0) begin
    end else begin
      s1_vaddr <= GEN_0;
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      refill_cnt <= GEN_2;
    end
    if(reset) begin
      T_968 <= 16'h1;
    end else begin
      T_968 <= GEN_3;
    end
    GEN_13 <= tag_array_0_tag_rdata_addr;
    GEN_14 <= tag_array_0_tag_rdata_en;
    if(tag_array_0_T_1019_en & tag_array_0_T_1019_mask) begin
      tag_array_0[tag_array_0_T_1019_addr] <= tag_array_0_T_1019_data;
    end
    GEN_16 <= tag_array_1_tag_rdata_addr;
    GEN_17 <= tag_array_1_tag_rdata_en;
    if(tag_array_1_T_1019_en & tag_array_1_T_1019_mask) begin
      tag_array_1[tag_array_1_T_1019_addr] <= tag_array_1_T_1019_data;
    end
    GEN_19 <= tag_array_2_tag_rdata_addr;
    GEN_20 <= tag_array_2_tag_rdata_en;
    if(tag_array_2_T_1019_en & tag_array_2_T_1019_mask) begin
      tag_array_2[tag_array_2_T_1019_addr] <= tag_array_2_T_1019_data;
    end
    GEN_22 <= tag_array_3_tag_rdata_addr;
    GEN_23 <= tag_array_3_tag_rdata_en;
    if(tag_array_3_T_1019_en & tag_array_3_T_1019_mask) begin
      tag_array_3[tag_array_3_T_1019_addr] <= tag_array_3_T_1019_data;
    end
    if(reset) begin
      vb_array <= 256'h0;
    end else begin
      vb_array <= GEN_38;
    end
    GEN_28 <= T_1199_T_1211_addr;
    GEN_30 <= T_1199_T_1211_en;
    if(T_1199_T_1204_en & T_1199_T_1204_mask) begin
      T_1199[T_1199_T_1204_addr] <= T_1199_T_1204_data;
    end
    GEN_40 <= T_1214_T_1226_addr;
    GEN_41 <= T_1214_T_1226_en;
    if(T_1214_T_1219_en & T_1214_T_1219_mask) begin
      T_1214[T_1214_T_1219_addr] <= T_1214_T_1219_data;
    end
    GEN_44 <= T_1229_T_1241_addr;
    GEN_45 <= T_1229_T_1241_en;
    if(T_1229_T_1234_en & T_1229_T_1234_mask) begin
      T_1229[T_1229_T_1234_addr] <= T_1229_T_1234_data;
    end
    GEN_47 <= T_1244_T_1256_addr;
    GEN_48 <= T_1244_T_1256_en;
    if(T_1244_T_1249_en & T_1244_T_1249_mask) begin
      T_1244[T_1244_T_1249_addr] <= T_1244_T_1249_data;
    end
  end
endmodule
module RocketCAM(
  input   clk,
  input   reset,
  input   io_clear,
  input  [7:0] io_clear_mask,
  input  [33:0] io_tag,
  output  io_hit,
  output [7:0] io_hits,
  output [7:0] io_valid_bits,
  input   io_write,
  input  [33:0] io_write_tag,
  input  [2:0] io_write_addr
);
  reg [33:0] cam_tags [0:7];
  reg [63:0] GEN_1;
  wire [33:0] cam_tags_T_25_data;
  wire [2:0] cam_tags_T_25_addr;
  wire  cam_tags_T_25_en;
  wire [33:0] cam_tags_T_30_data;
  wire [2:0] cam_tags_T_30_addr;
  wire  cam_tags_T_30_en;
  wire [33:0] cam_tags_T_35_data;
  wire [2:0] cam_tags_T_35_addr;
  wire  cam_tags_T_35_en;
  wire [33:0] cam_tags_T_40_data;
  wire [2:0] cam_tags_T_40_addr;
  wire  cam_tags_T_40_en;
  wire [33:0] cam_tags_T_45_data;
  wire [2:0] cam_tags_T_45_addr;
  wire  cam_tags_T_45_en;
  wire [33:0] cam_tags_T_50_data;
  wire [2:0] cam_tags_T_50_addr;
  wire  cam_tags_T_50_en;
  wire [33:0] cam_tags_T_55_data;
  wire [2:0] cam_tags_T_55_addr;
  wire  cam_tags_T_55_en;
  wire [33:0] cam_tags_T_60_data;
  wire [2:0] cam_tags_T_60_addr;
  wire  cam_tags_T_60_en;
  wire [33:0] cam_tags_T_20_data;
  wire [2:0] cam_tags_T_20_addr;
  wire  cam_tags_T_20_mask;
  wire  cam_tags_T_20_en;
  reg [7:0] vb_array;
  reg [31:0] GEN_2;
  wire [7:0] GEN_7;
  wire [7:0] T_14;
  wire [7:0] T_15;
  wire [7:0] GEN_0;
  wire [7:0] T_21;
  wire [7:0] T_22;
  wire [7:0] GEN_6;
  wire  T_23;
  wire  T_26;
  wire  T_27;
  wire  T_28;
  wire  T_31;
  wire  T_32;
  wire  T_33;
  wire  T_36;
  wire  T_37;
  wire  T_38;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_46;
  wire  T_47;
  wire  T_48;
  wire  T_51;
  wire  T_52;
  wire  T_53;
  wire  T_56;
  wire  T_57;
  wire  T_58;
  wire  T_61;
  wire  T_62;
  wire  T_68_0;
  wire  T_68_1;
  wire  T_68_2;
  wire  T_68_3;
  wire  T_68_4;
  wire  T_68_5;
  wire  T_68_6;
  wire  T_68_7;
  wire [1:0] T_70;
  wire [1:0] T_71;
  wire [3:0] T_72;
  wire [1:0] T_73;
  wire [1:0] T_74;
  wire [3:0] T_75;
  wire [7:0] T_76;
  wire [7:0] GEN_8;
  wire  T_78;
  assign io_hit = T_78;
  assign io_hits = T_76;
  assign io_valid_bits = vb_array;
  assign cam_tags_T_25_addr = {{2'd0}, 1'h0};
  assign cam_tags_T_25_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_25_data = cam_tags[cam_tags_T_25_addr];
  `else
  assign cam_tags_T_25_data = cam_tags_T_25_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_25_addr];
  `endif
  assign cam_tags_T_30_addr = {{2'd0}, 1'h1};
  assign cam_tags_T_30_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_30_data = cam_tags[cam_tags_T_30_addr];
  `else
  assign cam_tags_T_30_data = cam_tags_T_30_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_30_addr];
  `endif
  assign cam_tags_T_35_addr = {{1'd0}, 2'h2};
  assign cam_tags_T_35_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_35_data = cam_tags[cam_tags_T_35_addr];
  `else
  assign cam_tags_T_35_data = cam_tags_T_35_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_35_addr];
  `endif
  assign cam_tags_T_40_addr = {{1'd0}, 2'h3};
  assign cam_tags_T_40_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_40_data = cam_tags[cam_tags_T_40_addr];
  `else
  assign cam_tags_T_40_data = cam_tags_T_40_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_40_addr];
  `endif
  assign cam_tags_T_45_addr = 3'h4;
  assign cam_tags_T_45_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_45_data = cam_tags[cam_tags_T_45_addr];
  `else
  assign cam_tags_T_45_data = cam_tags_T_45_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_45_addr];
  `endif
  assign cam_tags_T_50_addr = 3'h5;
  assign cam_tags_T_50_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_50_data = cam_tags[cam_tags_T_50_addr];
  `else
  assign cam_tags_T_50_data = cam_tags_T_50_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_50_addr];
  `endif
  assign cam_tags_T_55_addr = 3'h6;
  assign cam_tags_T_55_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_55_data = cam_tags[cam_tags_T_55_addr];
  `else
  assign cam_tags_T_55_data = cam_tags_T_55_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_55_addr];
  `endif
  assign cam_tags_T_60_addr = 3'h7;
  assign cam_tags_T_60_en = 1'h1;
  `ifdef SYNTHESIS
  assign cam_tags_T_60_data = cam_tags[cam_tags_T_60_addr];
  `else
  assign cam_tags_T_60_data = cam_tags_T_60_addr >= 4'h8 ? $random : cam_tags[cam_tags_T_60_addr];
  `endif
  assign cam_tags_T_20_data = io_write_tag;
  assign cam_tags_T_20_addr = io_write_addr;
  assign cam_tags_T_20_mask = io_write;
  assign cam_tags_T_20_en = io_write;
  assign GEN_7 = {{7'd0}, 1'h1};
  assign T_14 = GEN_7 << io_write_addr;
  assign T_15 = vb_array | T_14;
  assign GEN_0 = io_write ? T_15 : vb_array;
  assign T_21 = ~ io_clear_mask;
  assign T_22 = vb_array & T_21;
  assign GEN_6 = io_clear ? T_22 : GEN_0;
  assign T_23 = vb_array[0];
  assign T_26 = cam_tags_T_25_data == io_tag;
  assign T_27 = T_23 & T_26;
  assign T_28 = vb_array[1];
  assign T_31 = cam_tags_T_30_data == io_tag;
  assign T_32 = T_28 & T_31;
  assign T_33 = vb_array[2];
  assign T_36 = cam_tags_T_35_data == io_tag;
  assign T_37 = T_33 & T_36;
  assign T_38 = vb_array[3];
  assign T_41 = cam_tags_T_40_data == io_tag;
  assign T_42 = T_38 & T_41;
  assign T_43 = vb_array[4];
  assign T_46 = cam_tags_T_45_data == io_tag;
  assign T_47 = T_43 & T_46;
  assign T_48 = vb_array[5];
  assign T_51 = cam_tags_T_50_data == io_tag;
  assign T_52 = T_48 & T_51;
  assign T_53 = vb_array[6];
  assign T_56 = cam_tags_T_55_data == io_tag;
  assign T_57 = T_53 & T_56;
  assign T_58 = vb_array[7];
  assign T_61 = cam_tags_T_60_data == io_tag;
  assign T_62 = T_58 & T_61;
  assign T_68_0 = T_27;
  assign T_68_1 = T_32;
  assign T_68_2 = T_37;
  assign T_68_3 = T_42;
  assign T_68_4 = T_47;
  assign T_68_5 = T_52;
  assign T_68_6 = T_57;
  assign T_68_7 = T_62;
  assign T_70 = {T_68_1,T_68_0};
  assign T_71 = {T_68_3,T_68_2};
  assign T_72 = {T_71,T_70};
  assign T_73 = {T_68_5,T_68_4};
  assign T_74 = {T_68_7,T_68_6};
  assign T_75 = {T_74,T_73};
  assign T_76 = {T_75,T_72};
  assign GEN_8 = {{7'd0}, 1'h0};
  assign T_78 = io_hits != GEN_8;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    cam_tags[initvar] = GEN_1[33:0];
  GEN_2 = {1{$random}};
  vb_array = GEN_2[7:0];
  end
`endif
  always @(posedge clk) begin
    if(cam_tags_T_20_en & cam_tags_T_20_mask) begin
      cam_tags[cam_tags_T_20_addr] <= cam_tags_T_20_data;
    end
    if(reset) begin
      vb_array <= 8'h0;
    end else begin
      vb_array <= GEN_6;
    end
  end
endmodule
module TLB(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [6:0] io_req_bits_asid,
  input  [27:0] io_req_bits_vpn,
  input   io_req_bits_passthrough,
  input   io_req_bits_instruction,
  input   io_req_bits_store,
  output  io_resp_miss,
  output [19:0] io_resp_ppn,
  output  io_resp_xcpt_ld,
  output  io_resp_xcpt_st,
  output  io_resp_xcpt_if,
  output [7:0] io_resp_hit_idx,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_ptw_invalidate
);
  wire  tag_cam_clk;
  wire  tag_cam_reset;
  wire  tag_cam_io_clear;
  wire [7:0] tag_cam_io_clear_mask;
  wire [33:0] tag_cam_io_tag;
  wire  tag_cam_io_hit;
  wire [7:0] tag_cam_io_hits;
  wire [7:0] tag_cam_io_valid_bits;
  wire  tag_cam_io_write;
  wire [33:0] tag_cam_io_write_tag;
  wire [2:0] tag_cam_io_write_addr;
  reg [19:0] tag_ram [0:7];
  reg [31:0] GEN_63;
  wire [19:0] tag_ram_T_562_data;
  wire [2:0] tag_ram_T_562_addr;
  wire  tag_ram_T_562_en;
  wire [19:0] tag_ram_T_564_data;
  wire [2:0] tag_ram_T_564_addr;
  wire  tag_ram_T_564_en;
  wire [19:0] tag_ram_T_566_data;
  wire [2:0] tag_ram_T_566_addr;
  wire  tag_ram_T_566_en;
  wire [19:0] tag_ram_T_568_data;
  wire [2:0] tag_ram_T_568_addr;
  wire  tag_ram_T_568_en;
  wire [19:0] tag_ram_T_570_data;
  wire [2:0] tag_ram_T_570_addr;
  wire  tag_ram_T_570_en;
  wire [19:0] tag_ram_T_572_data;
  wire [2:0] tag_ram_T_572_addr;
  wire  tag_ram_T_572_en;
  wire [19:0] tag_ram_T_574_data;
  wire [2:0] tag_ram_T_574_addr;
  wire  tag_ram_T_574_en;
  wire [19:0] tag_ram_T_576_data;
  wire [2:0] tag_ram_T_576_addr;
  wire  tag_ram_T_576_en;
  wire [19:0] tag_ram_T_232_data;
  wire [2:0] tag_ram_T_232_addr;
  wire  tag_ram_T_232_mask;
  wire  tag_ram_T_232_en;
  reg [1:0] state;
  reg [31:0] GEN_64;
  reg [33:0] r_refill_tag;
  reg [63:0] GEN_65;
  reg [2:0] r_refill_waddr;
  reg [31:0] GEN_66;
  reg [6:0] r_req_asid;
  reg [31:0] GEN_67;
  reg [27:0] r_req_vpn;
  reg [31:0] GEN_68;
  reg  r_req_passthrough;
  reg [31:0] GEN_77;
  reg  r_req_instruction;
  reg [31:0] GEN_86;
  reg  r_req_store;
  reg [31:0] GEN_95;
  wire [26:0] T_168;
  wire [33:0] lookup_tag;
  wire  T_169;
  wire  T_170;
  wire [3:0] T_171;
  wire [3:0] T_172;
  wire [3:0] GEN_146;
  wire  T_174;
  wire [3:0] T_175;
  wire [1:0] T_176;
  wire [1:0] T_177;
  wire [1:0] GEN_147;
  wire  T_179;
  wire [1:0] T_180;
  wire  T_181;
  wire [1:0] T_182;
  wire [2:0] tag_hit_addr;
  reg  ur_array_0;
  reg [31:0] GEN_104;
  reg  ur_array_1;
  reg [31:0] GEN_113;
  reg  ur_array_2;
  reg [31:0] GEN_122;
  reg  ur_array_3;
  reg [31:0] GEN_153;
  reg  ur_array_4;
  reg [31:0] GEN_154;
  reg  ur_array_5;
  reg [31:0] GEN_155;
  reg  ur_array_6;
  reg [31:0] GEN_156;
  reg  ur_array_7;
  reg [31:0] GEN_157;
  reg  uw_array_0;
  reg [31:0] GEN_158;
  reg  uw_array_1;
  reg [31:0] GEN_159;
  reg  uw_array_2;
  reg [31:0] GEN_160;
  reg  uw_array_3;
  reg [31:0] GEN_161;
  reg  uw_array_4;
  reg [31:0] GEN_162;
  reg  uw_array_5;
  reg [31:0] GEN_163;
  reg  uw_array_6;
  reg [31:0] GEN_164;
  reg  uw_array_7;
  reg [31:0] GEN_165;
  reg  ux_array_0;
  reg [31:0] GEN_166;
  reg  ux_array_1;
  reg [31:0] GEN_167;
  reg  ux_array_2;
  reg [31:0] GEN_168;
  reg  ux_array_3;
  reg [31:0] GEN_169;
  reg  ux_array_4;
  reg [31:0] GEN_170;
  reg  ux_array_5;
  reg [31:0] GEN_171;
  reg  ux_array_6;
  reg [31:0] GEN_172;
  reg  ux_array_7;
  reg [31:0] GEN_174;
  reg  sr_array_0;
  reg [31:0] GEN_175;
  reg  sr_array_1;
  reg [31:0] GEN_176;
  reg  sr_array_2;
  reg [31:0] GEN_177;
  reg  sr_array_3;
  reg [31:0] GEN_178;
  reg  sr_array_4;
  reg [31:0] GEN_179;
  reg  sr_array_5;
  reg [31:0] GEN_180;
  reg  sr_array_6;
  reg [31:0] GEN_181;
  reg  sr_array_7;
  reg [31:0] GEN_184;
  reg  sw_array_0;
  reg [31:0] GEN_185;
  reg  sw_array_1;
  reg [31:0] GEN_186;
  reg  sw_array_2;
  reg [31:0] GEN_187;
  reg  sw_array_3;
  reg [31:0] GEN_192;
  reg  sw_array_4;
  reg [31:0] GEN_194;
  reg  sw_array_5;
  reg [31:0] GEN_198;
  reg  sw_array_6;
  reg [31:0] GEN_201;
  reg  sw_array_7;
  reg [31:0] GEN_202;
  reg  sx_array_0;
  reg [31:0] GEN_203;
  reg  sx_array_1;
  reg [31:0] GEN_204;
  reg  sx_array_2;
  reg [31:0] GEN_205;
  reg  sx_array_3;
  reg [31:0] GEN_206;
  reg  sx_array_4;
  reg [31:0] GEN_207;
  reg  sx_array_5;
  reg [31:0] GEN_208;
  reg  sx_array_6;
  reg [31:0] GEN_209;
  reg  sx_array_7;
  reg [31:0] GEN_210;
  reg  dirty_array_0;
  reg [31:0] GEN_211;
  reg  dirty_array_1;
  reg [31:0] GEN_212;
  reg  dirty_array_2;
  reg [31:0] GEN_213;
  reg  dirty_array_3;
  reg [31:0] GEN_214;
  reg  dirty_array_4;
  reg [31:0] GEN_215;
  reg  dirty_array_5;
  reg [31:0] GEN_216;
  reg  dirty_array_6;
  reg [31:0] GEN_217;
  reg  dirty_array_7;
  reg [31:0] GEN_218;
  wire [3:0] GEN_148;
  wire  T_234;
  wire  T_235;
  wire  T_237;
  wire  T_238;
  wire  GEN_0;
  wire [2:0] GEN_149;
  wire  GEN_7;
  wire [2:0] GEN_150;
  wire  GEN_8;
  wire [2:0] GEN_151;
  wire  GEN_9;
  wire [2:0] GEN_152;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  T_245;
  wire  T_246;
  wire  GEN_1;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire  GEN_21;
  wire  GEN_22;
  wire  T_253;
  wire  T_254;
  wire  GEN_2;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_3;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  wire  GEN_38;
  wire  T_262;
  wire  GEN_4;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire [3:0] GEN_173;
  wire  T_264;
  wire  T_265;
  wire  T_267;
  wire  GEN_5;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_6;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire [7:0] T_268;
  wire [7:0] GEN_182;
  wire  T_270;
  wire  has_invalid_entry;
  wire  T_273;
  wire  T_274;
  wire  T_275;
  wire  T_276;
  wire  T_277;
  wire  T_278;
  wire  T_279;
  wire [2:0] T_289;
  wire [2:0] T_290;
  wire [2:0] T_291;
  wire [2:0] T_292;
  wire [2:0] T_293;
  wire [2:0] T_294;
  wire [2:0] invalid_entry;
  reg [7:0] T_296;
  reg [31:0] GEN_219;
  wire [7:0] T_298;
  wire  T_299;
  wire [1:0] T_300;
  wire [7:0] T_301;
  wire  T_302;
  wire [2:0] T_303;
  wire [7:0] T_304;
  wire  T_305;
  wire [3:0] T_306;
  wire [2:0] T_307;
  wire [2:0] repl_waddr;
  wire  T_309;
  wire  do_mprv;
  wire [1:0] priv;
  wire [1:0] GEN_183;
  wire  priv_s;
  wire  T_312;
  wire  T_314;
  wire  priv_uses_vm;
  wire [1:0] T_321;
  wire [1:0] T_322;
  wire [3:0] T_323;
  wire [1:0] T_324;
  wire [1:0] T_325;
  wire [3:0] T_326;
  wire [7:0] ur_bits;
  wire [7:0] T_328;
  wire [7:0] pum_ok;
  wire [1:0] T_329;
  wire [1:0] T_330;
  wire [3:0] T_331;
  wire [1:0] T_332;
  wire [1:0] T_333;
  wire [3:0] T_334;
  wire [7:0] T_335;
  wire [7:0] T_336;
  wire [7:0] r_array;
  wire [1:0] T_337;
  wire [1:0] T_338;
  wire [3:0] T_339;
  wire [1:0] T_340;
  wire [1:0] T_341;
  wire [3:0] T_342;
  wire [7:0] T_343;
  wire [7:0] T_344;
  wire [1:0] T_345;
  wire [1:0] T_346;
  wire [3:0] T_347;
  wire [1:0] T_348;
  wire [1:0] T_349;
  wire [3:0] T_350;
  wire [7:0] T_351;
  wire [7:0] w_array;
  wire [1:0] T_352;
  wire [1:0] T_353;
  wire [3:0] T_354;
  wire [1:0] T_355;
  wire [1:0] T_356;
  wire [3:0] T_357;
  wire [7:0] T_358;
  wire [1:0] T_359;
  wire [1:0] T_360;
  wire [3:0] T_361;
  wire [1:0] T_362;
  wire [1:0] T_363;
  wire [3:0] T_364;
  wire [7:0] T_365;
  wire [7:0] x_array;
  wire  T_367;
  wire  T_369;
  wire  T_371;
  wire  vm_enabled;
  wire  T_372;
  wire  T_373;
  wire  bad_va;
  wire [1:0] T_374;
  wire [1:0] T_375;
  wire [3:0] T_376;
  wire [1:0] T_377;
  wire [1:0] T_378;
  wire [3:0] T_379;
  wire [7:0] T_380;
  wire [7:0] T_382;
  wire [7:0] T_383;
  wire [7:0] T_384;
  wire [7:0] tag_hits;
  wire  tag_hit;
  wire  tlb_hit;
  wire  T_387;
  wire  T_388;
  wire  T_390;
  wire  tlb_miss;
  wire  T_391;
  wire  T_406;
  wire [8:0] GEN_188;
  wire [8:0] T_408;
  wire [7:0] T_409;
  wire [7:0] T_410;
  wire [7:0] T_411;
  wire [7:0] T_413;
  wire [7:0] T_414;
  wire [1:0] T_415;
  wire  T_416;
  wire [10:0] GEN_189;
  wire [10:0] T_418;
  wire [7:0] T_419;
  wire [7:0] T_420;
  wire [7:0] T_421;
  wire [7:0] T_423;
  wire [7:0] T_424;
  wire [2:0] T_425;
  wire  T_426;
  wire [14:0] GEN_190;
  wire [14:0] T_428;
  wire [7:0] T_429;
  wire [7:0] T_430;
  wire [7:0] T_431;
  wire [7:0] T_433;
  wire [7:0] T_434;
  wire [7:0] GEN_131;
  wire [31:0] paddr;
  wire [31:0] GEN_191;
  wire  T_440;
  wire [2:0] T_444;
  wire  T_446;
  wire [31:0] GEN_193;
  wire  T_448;
  wire  T_449;
  wire [2:0] T_452;
  wire  T_454;
  wire [31:0] GEN_195;
  wire  T_456;
  wire  T_457;
  wire [2:0] T_460;
  wire [31:0] GEN_196;
  wire  T_462;
  wire [31:0] GEN_197;
  wire  T_464;
  wire  T_465;
  wire [2:0] T_468;
  wire  T_470;
  wire [31:0] GEN_199;
  wire  T_472;
  wire  T_473;
  wire [2:0] T_476;
  wire [31:0] GEN_200;
  wire  T_478;
  wire  T_480;
  wire  T_481;
  wire [2:0] T_484;
  wire  T_486;
  wire [2:0] T_492;
  wire [2:0] T_497;
  wire [2:0] T_498;
  wire [2:0] T_499;
  wire [2:0] T_500;
  wire [2:0] T_501;
  wire [2:0] T_502;
  wire  addr_prot_x;
  wire  addr_prot_w;
  wire  addr_prot_r;
  wire  T_510;
  wire  T_511;
  wire  T_512;
  wire  T_513;
  wire  T_515;
  wire  T_517;
  wire  T_518;
  wire  T_519;
  wire [7:0] T_520;
  wire  T_522;
  wire  T_524;
  wire  T_525;
  wire  T_526;
  wire  T_530;
  wire  T_531;
  wire  T_532;
  wire [7:0] T_533;
  wire  T_535;
  wire  T_537;
  wire  T_538;
  wire  T_539;
  wire  T_543;
  wire  T_544;
  wire  T_545;
  wire [7:0] T_546;
  wire  T_548;
  wire  T_550;
  wire  T_551;
  wire  T_552;
  wire  T_553;
  wire  T_554;
  wire  T_555;
  wire  T_556;
  wire  T_557;
  wire  T_558;
  wire  T_559;
  wire  T_560;
  wire [19:0] T_578;
  wire [19:0] T_580;
  wire [19:0] T_582;
  wire [19:0] T_584;
  wire [19:0] T_586;
  wire [19:0] T_588;
  wire [19:0] T_590;
  wire [19:0] T_592;
  wire [19:0] T_594;
  wire [19:0] T_595;
  wire [19:0] T_596;
  wire [19:0] T_597;
  wire [19:0] T_598;
  wire [19:0] T_599;
  wire [19:0] T_600;
  wire [19:0] T_601;
  wire [19:0] T_602;
  wire [19:0] T_603;
  wire  T_606;
  wire  T_607;
  wire  T_608;
  wire [1:0] GEN_132;
  wire [33:0] GEN_133;
  wire [2:0] GEN_134;
  wire [6:0] GEN_135;
  wire [27:0] GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire [1:0] GEN_140;
  wire [1:0] GEN_141;
  wire [1:0] GEN_142;
  wire [1:0] GEN_143;
  wire  T_611;
  wire [1:0] GEN_144;
  wire [1:0] GEN_145;
  RocketCAM tag_cam (
    .clk(tag_cam_clk),
    .reset(tag_cam_reset),
    .io_clear(tag_cam_io_clear),
    .io_clear_mask(tag_cam_io_clear_mask),
    .io_tag(tag_cam_io_tag),
    .io_hit(tag_cam_io_hit),
    .io_hits(tag_cam_io_hits),
    .io_valid_bits(tag_cam_io_valid_bits),
    .io_write(tag_cam_io_write),
    .io_write_tag(tag_cam_io_write_tag),
    .io_write_addr(tag_cam_io_write_addr)
  );
  assign io_req_ready = T_513;
  assign io_resp_miss = tlb_miss;
  assign io_resp_ppn = T_603;
  assign io_resp_xcpt_ld = T_526;
  assign io_resp_xcpt_st = T_539;
  assign io_resp_xcpt_if = T_552;
  assign io_resp_hit_idx = tag_cam_io_hits;
  assign io_ptw_req_valid = T_606;
  assign io_ptw_req_bits_addr = r_refill_tag[26:0];
  assign io_ptw_req_bits_prv = io_ptw_status_prv;
  assign io_ptw_req_bits_store = r_req_store;
  assign io_ptw_req_bits_fetch = r_req_instruction;
  assign tag_cam_clk = clk;
  assign tag_cam_reset = reset;
  assign tag_cam_io_clear = io_ptw_invalidate;
  assign tag_cam_io_clear_mask = 8'hff;
  assign tag_cam_io_tag = lookup_tag;
  assign tag_cam_io_write = T_170;
  assign tag_cam_io_write_tag = r_refill_tag;
  assign tag_cam_io_write_addr = r_refill_waddr;
  assign tag_ram_T_562_addr = {{2'd0}, 1'h0};
  assign tag_ram_T_562_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_562_data = tag_ram[tag_ram_T_562_addr];
  `else
  assign tag_ram_T_562_data = tag_ram_T_562_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_562_addr];
  `endif
  assign tag_ram_T_564_addr = {{2'd0}, 1'h1};
  assign tag_ram_T_564_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_564_data = tag_ram[tag_ram_T_564_addr];
  `else
  assign tag_ram_T_564_data = tag_ram_T_564_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_564_addr];
  `endif
  assign tag_ram_T_566_addr = {{1'd0}, 2'h2};
  assign tag_ram_T_566_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_566_data = tag_ram[tag_ram_T_566_addr];
  `else
  assign tag_ram_T_566_data = tag_ram_T_566_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_566_addr];
  `endif
  assign tag_ram_T_568_addr = {{1'd0}, 2'h3};
  assign tag_ram_T_568_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_568_data = tag_ram[tag_ram_T_568_addr];
  `else
  assign tag_ram_T_568_data = tag_ram_T_568_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_568_addr];
  `endif
  assign tag_ram_T_570_addr = 3'h4;
  assign tag_ram_T_570_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_570_data = tag_ram[tag_ram_T_570_addr];
  `else
  assign tag_ram_T_570_data = tag_ram_T_570_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_570_addr];
  `endif
  assign tag_ram_T_572_addr = 3'h5;
  assign tag_ram_T_572_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_572_data = tag_ram[tag_ram_T_572_addr];
  `else
  assign tag_ram_T_572_data = tag_ram_T_572_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_572_addr];
  `endif
  assign tag_ram_T_574_addr = 3'h6;
  assign tag_ram_T_574_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_574_data = tag_ram[tag_ram_T_574_addr];
  `else
  assign tag_ram_T_574_data = tag_ram_T_574_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_574_addr];
  `endif
  assign tag_ram_T_576_addr = 3'h7;
  assign tag_ram_T_576_en = 1'h1;
  `ifdef SYNTHESIS
  assign tag_ram_T_576_data = tag_ram[tag_ram_T_576_addr];
  `else
  assign tag_ram_T_576_data = tag_ram_T_576_addr >= 4'h8 ? $random : tag_ram[tag_ram_T_576_addr];
  `endif
  assign tag_ram_T_232_data = io_ptw_resp_bits_pte_ppn;
  assign tag_ram_T_232_addr = r_refill_waddr;
  assign tag_ram_T_232_mask = io_ptw_resp_valid;
  assign tag_ram_T_232_en = io_ptw_resp_valid;
  assign T_168 = io_req_bits_vpn[26:0];
  assign lookup_tag = {io_req_bits_asid,T_168};
  assign T_169 = state == 2'h2;
  assign T_170 = T_169 & io_ptw_resp_valid;
  assign T_171 = tag_cam_io_hits[7:4];
  assign T_172 = tag_cam_io_hits[3:0];
  assign GEN_146 = {{3'd0}, 1'h0};
  assign T_174 = T_171 != GEN_146;
  assign T_175 = T_171 | T_172;
  assign T_176 = T_175[3:2];
  assign T_177 = T_175[1:0];
  assign GEN_147 = {{1'd0}, 1'h0};
  assign T_179 = T_176 != GEN_147;
  assign T_180 = T_176 | T_177;
  assign T_181 = T_180[1];
  assign T_182 = {T_179,T_181};
  assign tag_hit_addr = {T_174,T_182};
  assign GEN_148 = {{2'd0}, 2'h2};
  assign T_234 = io_ptw_resp_bits_pte_typ >= GEN_148;
  assign T_235 = io_ptw_resp_bits_pte_v & T_234;
  assign T_237 = io_ptw_resp_bits_pte_typ < 4'h8;
  assign T_238 = T_235 & T_237;
  assign GEN_0 = T_238;
  assign GEN_149 = {{2'd0}, 1'h0};
  assign GEN_7 = GEN_149 == r_refill_waddr ? GEN_0 : ur_array_0;
  assign GEN_150 = {{2'd0}, 1'h1};
  assign GEN_8 = GEN_150 == r_refill_waddr ? GEN_0 : ur_array_1;
  assign GEN_151 = {{1'd0}, 2'h2};
  assign GEN_9 = GEN_151 == r_refill_waddr ? GEN_0 : ur_array_2;
  assign GEN_152 = {{1'd0}, 2'h3};
  assign GEN_10 = GEN_152 == r_refill_waddr ? GEN_0 : ur_array_3;
  assign GEN_11 = 3'h4 == r_refill_waddr ? GEN_0 : ur_array_4;
  assign GEN_12 = 3'h5 == r_refill_waddr ? GEN_0 : ur_array_5;
  assign GEN_13 = 3'h6 == r_refill_waddr ? GEN_0 : ur_array_6;
  assign GEN_14 = 3'h7 == r_refill_waddr ? GEN_0 : ur_array_7;
  assign T_245 = io_ptw_resp_bits_pte_typ[0];
  assign T_246 = T_238 & T_245;
  assign GEN_1 = T_246;
  assign GEN_15 = GEN_149 == r_refill_waddr ? GEN_1 : uw_array_0;
  assign GEN_16 = GEN_150 == r_refill_waddr ? GEN_1 : uw_array_1;
  assign GEN_17 = GEN_151 == r_refill_waddr ? GEN_1 : uw_array_2;
  assign GEN_18 = GEN_152 == r_refill_waddr ? GEN_1 : uw_array_3;
  assign GEN_19 = 3'h4 == r_refill_waddr ? GEN_1 : uw_array_4;
  assign GEN_20 = 3'h5 == r_refill_waddr ? GEN_1 : uw_array_5;
  assign GEN_21 = 3'h6 == r_refill_waddr ? GEN_1 : uw_array_6;
  assign GEN_22 = 3'h7 == r_refill_waddr ? GEN_1 : uw_array_7;
  assign T_253 = io_ptw_resp_bits_pte_typ[1];
  assign T_254 = T_238 & T_253;
  assign GEN_2 = T_254;
  assign GEN_23 = GEN_149 == r_refill_waddr ? GEN_2 : ux_array_0;
  assign GEN_24 = GEN_150 == r_refill_waddr ? GEN_2 : ux_array_1;
  assign GEN_25 = GEN_151 == r_refill_waddr ? GEN_2 : ux_array_2;
  assign GEN_26 = GEN_152 == r_refill_waddr ? GEN_2 : ux_array_3;
  assign GEN_27 = 3'h4 == r_refill_waddr ? GEN_2 : ux_array_4;
  assign GEN_28 = 3'h5 == r_refill_waddr ? GEN_2 : ux_array_5;
  assign GEN_29 = 3'h6 == r_refill_waddr ? GEN_2 : ux_array_6;
  assign GEN_30 = 3'h7 == r_refill_waddr ? GEN_2 : ux_array_7;
  assign GEN_3 = T_235;
  assign GEN_31 = GEN_149 == r_refill_waddr ? GEN_3 : sr_array_0;
  assign GEN_32 = GEN_150 == r_refill_waddr ? GEN_3 : sr_array_1;
  assign GEN_33 = GEN_151 == r_refill_waddr ? GEN_3 : sr_array_2;
  assign GEN_34 = GEN_152 == r_refill_waddr ? GEN_3 : sr_array_3;
  assign GEN_35 = 3'h4 == r_refill_waddr ? GEN_3 : sr_array_4;
  assign GEN_36 = 3'h5 == r_refill_waddr ? GEN_3 : sr_array_5;
  assign GEN_37 = 3'h6 == r_refill_waddr ? GEN_3 : sr_array_6;
  assign GEN_38 = 3'h7 == r_refill_waddr ? GEN_3 : sr_array_7;
  assign T_262 = T_235 & T_245;
  assign GEN_4 = T_262;
  assign GEN_39 = GEN_149 == r_refill_waddr ? GEN_4 : sw_array_0;
  assign GEN_40 = GEN_150 == r_refill_waddr ? GEN_4 : sw_array_1;
  assign GEN_41 = GEN_151 == r_refill_waddr ? GEN_4 : sw_array_2;
  assign GEN_42 = GEN_152 == r_refill_waddr ? GEN_4 : sw_array_3;
  assign GEN_43 = 3'h4 == r_refill_waddr ? GEN_4 : sw_array_4;
  assign GEN_44 = 3'h5 == r_refill_waddr ? GEN_4 : sw_array_5;
  assign GEN_45 = 3'h6 == r_refill_waddr ? GEN_4 : sw_array_6;
  assign GEN_46 = 3'h7 == r_refill_waddr ? GEN_4 : sw_array_7;
  assign GEN_173 = {{1'd0}, 3'h4};
  assign T_264 = io_ptw_resp_bits_pte_typ >= GEN_173;
  assign T_265 = io_ptw_resp_bits_pte_v & T_264;
  assign T_267 = T_265 & T_253;
  assign GEN_5 = T_267;
  assign GEN_47 = GEN_149 == r_refill_waddr ? GEN_5 : sx_array_0;
  assign GEN_48 = GEN_150 == r_refill_waddr ? GEN_5 : sx_array_1;
  assign GEN_49 = GEN_151 == r_refill_waddr ? GEN_5 : sx_array_2;
  assign GEN_50 = GEN_152 == r_refill_waddr ? GEN_5 : sx_array_3;
  assign GEN_51 = 3'h4 == r_refill_waddr ? GEN_5 : sx_array_4;
  assign GEN_52 = 3'h5 == r_refill_waddr ? GEN_5 : sx_array_5;
  assign GEN_53 = 3'h6 == r_refill_waddr ? GEN_5 : sx_array_6;
  assign GEN_54 = 3'h7 == r_refill_waddr ? GEN_5 : sx_array_7;
  assign GEN_6 = io_ptw_resp_bits_pte_d;
  assign GEN_55 = GEN_149 == r_refill_waddr ? GEN_6 : dirty_array_0;
  assign GEN_56 = GEN_150 == r_refill_waddr ? GEN_6 : dirty_array_1;
  assign GEN_57 = GEN_151 == r_refill_waddr ? GEN_6 : dirty_array_2;
  assign GEN_58 = GEN_152 == r_refill_waddr ? GEN_6 : dirty_array_3;
  assign GEN_59 = 3'h4 == r_refill_waddr ? GEN_6 : dirty_array_4;
  assign GEN_60 = 3'h5 == r_refill_waddr ? GEN_6 : dirty_array_5;
  assign GEN_61 = 3'h6 == r_refill_waddr ? GEN_6 : dirty_array_6;
  assign GEN_62 = 3'h7 == r_refill_waddr ? GEN_6 : dirty_array_7;
  assign GEN_69 = io_ptw_resp_valid ? GEN_7 : ur_array_0;
  assign GEN_70 = io_ptw_resp_valid ? GEN_8 : ur_array_1;
  assign GEN_71 = io_ptw_resp_valid ? GEN_9 : ur_array_2;
  assign GEN_72 = io_ptw_resp_valid ? GEN_10 : ur_array_3;
  assign GEN_73 = io_ptw_resp_valid ? GEN_11 : ur_array_4;
  assign GEN_74 = io_ptw_resp_valid ? GEN_12 : ur_array_5;
  assign GEN_75 = io_ptw_resp_valid ? GEN_13 : ur_array_6;
  assign GEN_76 = io_ptw_resp_valid ? GEN_14 : ur_array_7;
  assign GEN_78 = io_ptw_resp_valid ? GEN_15 : uw_array_0;
  assign GEN_79 = io_ptw_resp_valid ? GEN_16 : uw_array_1;
  assign GEN_80 = io_ptw_resp_valid ? GEN_17 : uw_array_2;
  assign GEN_81 = io_ptw_resp_valid ? GEN_18 : uw_array_3;
  assign GEN_82 = io_ptw_resp_valid ? GEN_19 : uw_array_4;
  assign GEN_83 = io_ptw_resp_valid ? GEN_20 : uw_array_5;
  assign GEN_84 = io_ptw_resp_valid ? GEN_21 : uw_array_6;
  assign GEN_85 = io_ptw_resp_valid ? GEN_22 : uw_array_7;
  assign GEN_87 = io_ptw_resp_valid ? GEN_23 : ux_array_0;
  assign GEN_88 = io_ptw_resp_valid ? GEN_24 : ux_array_1;
  assign GEN_89 = io_ptw_resp_valid ? GEN_25 : ux_array_2;
  assign GEN_90 = io_ptw_resp_valid ? GEN_26 : ux_array_3;
  assign GEN_91 = io_ptw_resp_valid ? GEN_27 : ux_array_4;
  assign GEN_92 = io_ptw_resp_valid ? GEN_28 : ux_array_5;
  assign GEN_93 = io_ptw_resp_valid ? GEN_29 : ux_array_6;
  assign GEN_94 = io_ptw_resp_valid ? GEN_30 : ux_array_7;
  assign GEN_96 = io_ptw_resp_valid ? GEN_31 : sr_array_0;
  assign GEN_97 = io_ptw_resp_valid ? GEN_32 : sr_array_1;
  assign GEN_98 = io_ptw_resp_valid ? GEN_33 : sr_array_2;
  assign GEN_99 = io_ptw_resp_valid ? GEN_34 : sr_array_3;
  assign GEN_100 = io_ptw_resp_valid ? GEN_35 : sr_array_4;
  assign GEN_101 = io_ptw_resp_valid ? GEN_36 : sr_array_5;
  assign GEN_102 = io_ptw_resp_valid ? GEN_37 : sr_array_6;
  assign GEN_103 = io_ptw_resp_valid ? GEN_38 : sr_array_7;
  assign GEN_105 = io_ptw_resp_valid ? GEN_39 : sw_array_0;
  assign GEN_106 = io_ptw_resp_valid ? GEN_40 : sw_array_1;
  assign GEN_107 = io_ptw_resp_valid ? GEN_41 : sw_array_2;
  assign GEN_108 = io_ptw_resp_valid ? GEN_42 : sw_array_3;
  assign GEN_109 = io_ptw_resp_valid ? GEN_43 : sw_array_4;
  assign GEN_110 = io_ptw_resp_valid ? GEN_44 : sw_array_5;
  assign GEN_111 = io_ptw_resp_valid ? GEN_45 : sw_array_6;
  assign GEN_112 = io_ptw_resp_valid ? GEN_46 : sw_array_7;
  assign GEN_114 = io_ptw_resp_valid ? GEN_47 : sx_array_0;
  assign GEN_115 = io_ptw_resp_valid ? GEN_48 : sx_array_1;
  assign GEN_116 = io_ptw_resp_valid ? GEN_49 : sx_array_2;
  assign GEN_117 = io_ptw_resp_valid ? GEN_50 : sx_array_3;
  assign GEN_118 = io_ptw_resp_valid ? GEN_51 : sx_array_4;
  assign GEN_119 = io_ptw_resp_valid ? GEN_52 : sx_array_5;
  assign GEN_120 = io_ptw_resp_valid ? GEN_53 : sx_array_6;
  assign GEN_121 = io_ptw_resp_valid ? GEN_54 : sx_array_7;
  assign GEN_123 = io_ptw_resp_valid ? GEN_55 : dirty_array_0;
  assign GEN_124 = io_ptw_resp_valid ? GEN_56 : dirty_array_1;
  assign GEN_125 = io_ptw_resp_valid ? GEN_57 : dirty_array_2;
  assign GEN_126 = io_ptw_resp_valid ? GEN_58 : dirty_array_3;
  assign GEN_127 = io_ptw_resp_valid ? GEN_59 : dirty_array_4;
  assign GEN_128 = io_ptw_resp_valid ? GEN_60 : dirty_array_5;
  assign GEN_129 = io_ptw_resp_valid ? GEN_61 : dirty_array_6;
  assign GEN_130 = io_ptw_resp_valid ? GEN_62 : dirty_array_7;
  assign T_268 = ~ tag_cam_io_valid_bits;
  assign GEN_182 = {{7'd0}, 1'h0};
  assign T_270 = T_268 == GEN_182;
  assign has_invalid_entry = T_270 == 1'h0;
  assign T_273 = T_268[0];
  assign T_274 = T_268[1];
  assign T_275 = T_268[2];
  assign T_276 = T_268[3];
  assign T_277 = T_268[4];
  assign T_278 = T_268[5];
  assign T_279 = T_268[6];
  assign T_289 = T_279 ? 3'h6 : 3'h7;
  assign T_290 = T_278 ? 3'h5 : T_289;
  assign T_291 = T_277 ? 3'h4 : T_290;
  assign T_292 = T_276 ? {{1'd0}, 2'h3} : T_291;
  assign T_293 = T_275 ? {{1'd0}, 2'h2} : T_292;
  assign T_294 = T_274 ? {{2'd0}, 1'h1} : T_293;
  assign invalid_entry = T_273 ? {{2'd0}, 1'h0} : T_294;
  assign T_298 = T_296 >> 1'h1;
  assign T_299 = T_298[0];
  assign T_300 = {1'h1,T_299};
  assign T_301 = T_296 >> T_300;
  assign T_302 = T_301[0];
  assign T_303 = {T_300,T_302};
  assign T_304 = T_296 >> T_303;
  assign T_305 = T_304[0];
  assign T_306 = {T_303,T_305};
  assign T_307 = T_306[2:0];
  assign repl_waddr = has_invalid_entry ? invalid_entry : T_307;
  assign T_309 = io_req_bits_instruction == 1'h0;
  assign do_mprv = io_ptw_status_mprv & T_309;
  assign priv = do_mprv ? io_ptw_status_mpp : io_ptw_status_prv;
  assign GEN_183 = {{1'd0}, 1'h1};
  assign priv_s = priv == GEN_183;
  assign T_312 = priv <= GEN_183;
  assign T_314 = io_ptw_status_debug == 1'h0;
  assign priv_uses_vm = T_312 & T_314;
  assign T_321 = {ur_array_1,ur_array_0};
  assign T_322 = {ur_array_3,ur_array_2};
  assign T_323 = {T_322,T_321};
  assign T_324 = {ur_array_5,ur_array_4};
  assign T_325 = {ur_array_7,ur_array_6};
  assign T_326 = {T_325,T_324};
  assign ur_bits = {T_326,T_323};
  assign T_328 = io_ptw_status_pum ? ur_bits : {{7'd0}, 1'h0};
  assign pum_ok = ~ T_328;
  assign T_329 = {sr_array_1,sr_array_0};
  assign T_330 = {sr_array_3,sr_array_2};
  assign T_331 = {T_330,T_329};
  assign T_332 = {sr_array_5,sr_array_4};
  assign T_333 = {sr_array_7,sr_array_6};
  assign T_334 = {T_333,T_332};
  assign T_335 = {T_334,T_331};
  assign T_336 = T_335 & pum_ok;
  assign r_array = priv_s ? T_336 : ur_bits;
  assign T_337 = {sw_array_1,sw_array_0};
  assign T_338 = {sw_array_3,sw_array_2};
  assign T_339 = {T_338,T_337};
  assign T_340 = {sw_array_5,sw_array_4};
  assign T_341 = {sw_array_7,sw_array_6};
  assign T_342 = {T_341,T_340};
  assign T_343 = {T_342,T_339};
  assign T_344 = T_343 & pum_ok;
  assign T_345 = {uw_array_1,uw_array_0};
  assign T_346 = {uw_array_3,uw_array_2};
  assign T_347 = {T_346,T_345};
  assign T_348 = {uw_array_5,uw_array_4};
  assign T_349 = {uw_array_7,uw_array_6};
  assign T_350 = {T_349,T_348};
  assign T_351 = {T_350,T_347};
  assign w_array = priv_s ? T_344 : T_351;
  assign T_352 = {sx_array_1,sx_array_0};
  assign T_353 = {sx_array_3,sx_array_2};
  assign T_354 = {T_353,T_352};
  assign T_355 = {sx_array_5,sx_array_4};
  assign T_356 = {sx_array_7,sx_array_6};
  assign T_357 = {T_356,T_355};
  assign T_358 = {T_357,T_354};
  assign T_359 = {ux_array_1,ux_array_0};
  assign T_360 = {ux_array_3,ux_array_2};
  assign T_361 = {T_360,T_359};
  assign T_362 = {ux_array_5,ux_array_4};
  assign T_363 = {ux_array_7,ux_array_6};
  assign T_364 = {T_363,T_362};
  assign T_365 = {T_364,T_361};
  assign x_array = priv_s ? T_358 : T_365;
  assign T_367 = io_ptw_status_vm[3];
  assign T_369 = T_367 & priv_uses_vm;
  assign T_371 = io_req_bits_passthrough == 1'h0;
  assign vm_enabled = T_369 & T_371;
  assign T_372 = io_req_bits_vpn[27];
  assign T_373 = io_req_bits_vpn[26];
  assign bad_va = T_372 != T_373;
  assign T_374 = {dirty_array_1,dirty_array_0};
  assign T_375 = {dirty_array_3,dirty_array_2};
  assign T_376 = {T_375,T_374};
  assign T_377 = {dirty_array_5,dirty_array_4};
  assign T_378 = {dirty_array_7,dirty_array_6};
  assign T_379 = {T_378,T_377};
  assign T_380 = {T_379,T_376};
  assign T_382 = io_req_bits_store ? w_array : {{7'd0}, 1'h0};
  assign T_383 = ~ T_382;
  assign T_384 = T_380 | T_383;
  assign tag_hits = tag_cam_io_hits & T_384;
  assign tag_hit = tag_hits != GEN_182;
  assign tlb_hit = vm_enabled & tag_hit;
  assign T_387 = tag_hit == 1'h0;
  assign T_388 = vm_enabled & T_387;
  assign T_390 = bad_va == 1'h0;
  assign tlb_miss = T_388 & T_390;
  assign T_391 = io_req_valid & tlb_hit;
  assign T_406 = tag_hit_addr[2];
  assign GEN_188 = {{1'd0}, 8'h1};
  assign T_408 = GEN_188 << 1'h1;
  assign T_409 = T_408[7:0];
  assign T_410 = ~ T_409;
  assign T_411 = T_296 & T_410;
  assign T_413 = T_406 ? {{7'd0}, 1'h0} : T_409;
  assign T_414 = T_411 | T_413;
  assign T_415 = {1'h1,T_406};
  assign T_416 = tag_hit_addr[1];
  assign GEN_189 = {{3'd0}, 8'h1};
  assign T_418 = GEN_189 << T_415;
  assign T_419 = T_418[7:0];
  assign T_420 = ~ T_419;
  assign T_421 = T_414 & T_420;
  assign T_423 = T_416 ? {{7'd0}, 1'h0} : T_419;
  assign T_424 = T_421 | T_423;
  assign T_425 = {T_415,T_416};
  assign T_426 = tag_hit_addr[0];
  assign GEN_190 = {{7'd0}, 8'h1};
  assign T_428 = GEN_190 << T_425;
  assign T_429 = T_428[7:0];
  assign T_430 = ~ T_429;
  assign T_431 = T_424 & T_430;
  assign T_433 = T_426 ? {{7'd0}, 1'h0} : T_429;
  assign T_434 = T_431 | T_433;
  assign GEN_131 = T_391 ? T_434 : T_296;
  assign paddr = {io_resp_ppn,12'h0};
  assign GEN_191 = {{19'd0}, 13'h1000};
  assign T_440 = paddr < GEN_191;
  assign T_444 = T_440 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_446 = GEN_191 <= paddr;
  assign GEN_193 = {{18'd0}, 14'h2000};
  assign T_448 = paddr < GEN_193;
  assign T_449 = T_446 & T_448;
  assign T_452 = T_449 ? 3'h5 : {{2'd0}, 1'h0};
  assign T_454 = GEN_193 <= paddr;
  assign GEN_195 = {{18'd0}, 14'h3000};
  assign T_456 = paddr < GEN_195;
  assign T_457 = T_454 & T_456;
  assign T_460 = T_457 ? 3'h3 : {{2'd0}, 1'h0};
  assign GEN_196 = {{1'd0}, 31'h40000000};
  assign T_462 = GEN_196 <= paddr;
  assign GEN_197 = {{1'd0}, 31'h44000000};
  assign T_464 = paddr < GEN_197;
  assign T_465 = T_462 & T_464;
  assign T_468 = T_465 ? 3'h3 : {{2'd0}, 1'h0};
  assign T_470 = GEN_197 <= paddr;
  assign GEN_199 = {{1'd0}, 31'h48000000};
  assign T_472 = paddr < GEN_199;
  assign T_473 = T_470 & T_472;
  assign T_476 = T_473 ? 3'h3 : {{2'd0}, 1'h0};
  assign GEN_200 = {{1'd0}, 31'h60000000};
  assign T_478 = GEN_200 <= paddr;
  assign T_480 = paddr < 32'h80000000;
  assign T_481 = T_478 & T_480;
  assign T_484 = T_481 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_486 = 32'h80000000 <= paddr;
  assign T_492 = T_486 ? 3'h7 : {{2'd0}, 1'h0};
  assign T_497 = T_444 | T_452;
  assign T_498 = T_497 | T_460;
  assign T_499 = T_498 | T_468;
  assign T_500 = T_499 | T_476;
  assign T_501 = T_500 | T_484;
  assign T_502 = T_501 | T_492;
  assign addr_prot_x = T_512;
  assign addr_prot_w = T_511;
  assign addr_prot_r = T_510;
  assign T_510 = T_502[0];
  assign T_511 = T_502[1];
  assign T_512 = T_502[2];
  assign T_513 = state == 2'h0;
  assign T_515 = tlb_miss == 1'h0;
  assign T_517 = addr_prot_r == 1'h0;
  assign T_518 = T_515 & T_517;
  assign T_519 = bad_va | T_518;
  assign T_520 = r_array & tag_cam_io_hits;
  assign T_522 = T_520 != GEN_182;
  assign T_524 = T_522 == 1'h0;
  assign T_525 = tlb_hit & T_524;
  assign T_526 = T_519 | T_525;
  assign T_530 = addr_prot_w == 1'h0;
  assign T_531 = T_515 & T_530;
  assign T_532 = bad_va | T_531;
  assign T_533 = w_array & tag_cam_io_hits;
  assign T_535 = T_533 != GEN_182;
  assign T_537 = T_535 == 1'h0;
  assign T_538 = tlb_hit & T_537;
  assign T_539 = T_532 | T_538;
  assign T_543 = addr_prot_x == 1'h0;
  assign T_544 = T_515 & T_543;
  assign T_545 = bad_va | T_544;
  assign T_546 = x_array & tag_cam_io_hits;
  assign T_548 = T_546 != GEN_182;
  assign T_550 = T_548 == 1'h0;
  assign T_551 = tlb_hit & T_550;
  assign T_552 = T_545 | T_551;
  assign T_553 = tag_cam_io_hits[0];
  assign T_554 = tag_cam_io_hits[1];
  assign T_555 = tag_cam_io_hits[2];
  assign T_556 = tag_cam_io_hits[3];
  assign T_557 = tag_cam_io_hits[4];
  assign T_558 = tag_cam_io_hits[5];
  assign T_559 = tag_cam_io_hits[6];
  assign T_560 = tag_cam_io_hits[7];
  assign T_578 = T_553 ? tag_ram_T_562_data : {{19'd0}, 1'h0};
  assign T_580 = T_554 ? tag_ram_T_564_data : {{19'd0}, 1'h0};
  assign T_582 = T_555 ? tag_ram_T_566_data : {{19'd0}, 1'h0};
  assign T_584 = T_556 ? tag_ram_T_568_data : {{19'd0}, 1'h0};
  assign T_586 = T_557 ? tag_ram_T_570_data : {{19'd0}, 1'h0};
  assign T_588 = T_558 ? tag_ram_T_572_data : {{19'd0}, 1'h0};
  assign T_590 = T_559 ? tag_ram_T_574_data : {{19'd0}, 1'h0};
  assign T_592 = T_560 ? tag_ram_T_576_data : {{19'd0}, 1'h0};
  assign T_594 = T_578 | T_580;
  assign T_595 = T_594 | T_582;
  assign T_596 = T_595 | T_584;
  assign T_597 = T_596 | T_586;
  assign T_598 = T_597 | T_588;
  assign T_599 = T_598 | T_590;
  assign T_600 = T_599 | T_592;
  assign T_601 = T_600;
  assign T_602 = io_req_bits_vpn[19:0];
  assign T_603 = vm_enabled ? T_601 : T_602;
  assign T_606 = state == 2'h1;
  assign T_607 = io_req_ready & io_req_valid;
  assign T_608 = T_607 & tlb_miss;
  assign GEN_132 = T_608 ? 2'h1 : state;
  assign GEN_133 = T_608 ? lookup_tag : r_refill_tag;
  assign GEN_134 = T_608 ? repl_waddr : r_refill_waddr;
  assign GEN_135 = T_608 ? io_req_bits_asid : r_req_asid;
  assign GEN_136 = T_608 ? io_req_bits_vpn : r_req_vpn;
  assign GEN_137 = T_608 ? io_req_bits_passthrough : r_req_passthrough;
  assign GEN_138 = T_608 ? io_req_bits_instruction : r_req_instruction;
  assign GEN_139 = T_608 ? io_req_bits_store : r_req_store;
  assign GEN_140 = io_ptw_invalidate ? 2'h0 : GEN_132;
  assign GEN_141 = io_ptw_invalidate ? 2'h3 : 2'h2;
  assign GEN_142 = io_ptw_req_ready ? GEN_141 : GEN_140;
  assign GEN_143 = T_606 ? GEN_142 : GEN_132;
  assign T_611 = T_169 & io_ptw_invalidate;
  assign GEN_144 = T_611 ? 2'h3 : GEN_143;
  assign GEN_145 = io_ptw_resp_valid ? 2'h0 : GEN_144;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_63 = {1{$random}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    tag_ram[initvar] = GEN_63[19:0];
  GEN_64 = {1{$random}};
  state = GEN_64[1:0];
  GEN_65 = {2{$random}};
  r_refill_tag = GEN_65[33:0];
  GEN_66 = {1{$random}};
  r_refill_waddr = GEN_66[2:0];
  GEN_67 = {1{$random}};
  r_req_asid = GEN_67[6:0];
  GEN_68 = {1{$random}};
  r_req_vpn = GEN_68[27:0];
  GEN_77 = {1{$random}};
  r_req_passthrough = GEN_77[0:0];
  GEN_86 = {1{$random}};
  r_req_instruction = GEN_86[0:0];
  GEN_95 = {1{$random}};
  r_req_store = GEN_95[0:0];
  GEN_104 = {1{$random}};
  ur_array_0 = GEN_104[0:0];
  GEN_113 = {1{$random}};
  ur_array_1 = GEN_113[0:0];
  GEN_122 = {1{$random}};
  ur_array_2 = GEN_122[0:0];
  GEN_153 = {1{$random}};
  ur_array_3 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  ur_array_4 = GEN_154[0:0];
  GEN_155 = {1{$random}};
  ur_array_5 = GEN_155[0:0];
  GEN_156 = {1{$random}};
  ur_array_6 = GEN_156[0:0];
  GEN_157 = {1{$random}};
  ur_array_7 = GEN_157[0:0];
  GEN_158 = {1{$random}};
  uw_array_0 = GEN_158[0:0];
  GEN_159 = {1{$random}};
  uw_array_1 = GEN_159[0:0];
  GEN_160 = {1{$random}};
  uw_array_2 = GEN_160[0:0];
  GEN_161 = {1{$random}};
  uw_array_3 = GEN_161[0:0];
  GEN_162 = {1{$random}};
  uw_array_4 = GEN_162[0:0];
  GEN_163 = {1{$random}};
  uw_array_5 = GEN_163[0:0];
  GEN_164 = {1{$random}};
  uw_array_6 = GEN_164[0:0];
  GEN_165 = {1{$random}};
  uw_array_7 = GEN_165[0:0];
  GEN_166 = {1{$random}};
  ux_array_0 = GEN_166[0:0];
  GEN_167 = {1{$random}};
  ux_array_1 = GEN_167[0:0];
  GEN_168 = {1{$random}};
  ux_array_2 = GEN_168[0:0];
  GEN_169 = {1{$random}};
  ux_array_3 = GEN_169[0:0];
  GEN_170 = {1{$random}};
  ux_array_4 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  ux_array_5 = GEN_171[0:0];
  GEN_172 = {1{$random}};
  ux_array_6 = GEN_172[0:0];
  GEN_174 = {1{$random}};
  ux_array_7 = GEN_174[0:0];
  GEN_175 = {1{$random}};
  sr_array_0 = GEN_175[0:0];
  GEN_176 = {1{$random}};
  sr_array_1 = GEN_176[0:0];
  GEN_177 = {1{$random}};
  sr_array_2 = GEN_177[0:0];
  GEN_178 = {1{$random}};
  sr_array_3 = GEN_178[0:0];
  GEN_179 = {1{$random}};
  sr_array_4 = GEN_179[0:0];
  GEN_180 = {1{$random}};
  sr_array_5 = GEN_180[0:0];
  GEN_181 = {1{$random}};
  sr_array_6 = GEN_181[0:0];
  GEN_184 = {1{$random}};
  sr_array_7 = GEN_184[0:0];
  GEN_185 = {1{$random}};
  sw_array_0 = GEN_185[0:0];
  GEN_186 = {1{$random}};
  sw_array_1 = GEN_186[0:0];
  GEN_187 = {1{$random}};
  sw_array_2 = GEN_187[0:0];
  GEN_192 = {1{$random}};
  sw_array_3 = GEN_192[0:0];
  GEN_194 = {1{$random}};
  sw_array_4 = GEN_194[0:0];
  GEN_198 = {1{$random}};
  sw_array_5 = GEN_198[0:0];
  GEN_201 = {1{$random}};
  sw_array_6 = GEN_201[0:0];
  GEN_202 = {1{$random}};
  sw_array_7 = GEN_202[0:0];
  GEN_203 = {1{$random}};
  sx_array_0 = GEN_203[0:0];
  GEN_204 = {1{$random}};
  sx_array_1 = GEN_204[0:0];
  GEN_205 = {1{$random}};
  sx_array_2 = GEN_205[0:0];
  GEN_206 = {1{$random}};
  sx_array_3 = GEN_206[0:0];
  GEN_207 = {1{$random}};
  sx_array_4 = GEN_207[0:0];
  GEN_208 = {1{$random}};
  sx_array_5 = GEN_208[0:0];
  GEN_209 = {1{$random}};
  sx_array_6 = GEN_209[0:0];
  GEN_210 = {1{$random}};
  sx_array_7 = GEN_210[0:0];
  GEN_211 = {1{$random}};
  dirty_array_0 = GEN_211[0:0];
  GEN_212 = {1{$random}};
  dirty_array_1 = GEN_212[0:0];
  GEN_213 = {1{$random}};
  dirty_array_2 = GEN_213[0:0];
  GEN_214 = {1{$random}};
  dirty_array_3 = GEN_214[0:0];
  GEN_215 = {1{$random}};
  dirty_array_4 = GEN_215[0:0];
  GEN_216 = {1{$random}};
  dirty_array_5 = GEN_216[0:0];
  GEN_217 = {1{$random}};
  dirty_array_6 = GEN_217[0:0];
  GEN_218 = {1{$random}};
  dirty_array_7 = GEN_218[0:0];
  GEN_219 = {1{$random}};
  T_296 = GEN_219[7:0];
  end
`endif
  always @(posedge clk) begin
    if(tag_ram_T_232_en & tag_ram_T_232_mask) begin
      tag_ram[tag_ram_T_232_addr] <= tag_ram_T_232_data;
    end
    if(reset) begin
      state <= 2'h0;
    end else begin
      state <= GEN_145;
    end
    if(1'h0) begin
    end else begin
      r_refill_tag <= GEN_133;
    end
    if(1'h0) begin
    end else begin
      r_refill_waddr <= GEN_134;
    end
    if(1'h0) begin
    end else begin
      r_req_asid <= GEN_135;
    end
    if(1'h0) begin
    end else begin
      r_req_vpn <= GEN_136;
    end
    if(1'h0) begin
    end else begin
      r_req_passthrough <= GEN_137;
    end
    if(1'h0) begin
    end else begin
      r_req_instruction <= GEN_138;
    end
    if(1'h0) begin
    end else begin
      r_req_store <= GEN_139;
    end
    if(1'h0) begin
    end else begin
      ur_array_0 <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      ur_array_1 <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      ur_array_2 <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      ur_array_3 <= GEN_72;
    end
    if(1'h0) begin
    end else begin
      ur_array_4 <= GEN_73;
    end
    if(1'h0) begin
    end else begin
      ur_array_5 <= GEN_74;
    end
    if(1'h0) begin
    end else begin
      ur_array_6 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      ur_array_7 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      uw_array_0 <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      uw_array_1 <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      uw_array_2 <= GEN_80;
    end
    if(1'h0) begin
    end else begin
      uw_array_3 <= GEN_81;
    end
    if(1'h0) begin
    end else begin
      uw_array_4 <= GEN_82;
    end
    if(1'h0) begin
    end else begin
      uw_array_5 <= GEN_83;
    end
    if(1'h0) begin
    end else begin
      uw_array_6 <= GEN_84;
    end
    if(1'h0) begin
    end else begin
      uw_array_7 <= GEN_85;
    end
    if(1'h0) begin
    end else begin
      ux_array_0 <= GEN_87;
    end
    if(1'h0) begin
    end else begin
      ux_array_1 <= GEN_88;
    end
    if(1'h0) begin
    end else begin
      ux_array_2 <= GEN_89;
    end
    if(1'h0) begin
    end else begin
      ux_array_3 <= GEN_90;
    end
    if(1'h0) begin
    end else begin
      ux_array_4 <= GEN_91;
    end
    if(1'h0) begin
    end else begin
      ux_array_5 <= GEN_92;
    end
    if(1'h0) begin
    end else begin
      ux_array_6 <= GEN_93;
    end
    if(1'h0) begin
    end else begin
      ux_array_7 <= GEN_94;
    end
    if(1'h0) begin
    end else begin
      sr_array_0 <= GEN_96;
    end
    if(1'h0) begin
    end else begin
      sr_array_1 <= GEN_97;
    end
    if(1'h0) begin
    end else begin
      sr_array_2 <= GEN_98;
    end
    if(1'h0) begin
    end else begin
      sr_array_3 <= GEN_99;
    end
    if(1'h0) begin
    end else begin
      sr_array_4 <= GEN_100;
    end
    if(1'h0) begin
    end else begin
      sr_array_5 <= GEN_101;
    end
    if(1'h0) begin
    end else begin
      sr_array_6 <= GEN_102;
    end
    if(1'h0) begin
    end else begin
      sr_array_7 <= GEN_103;
    end
    if(1'h0) begin
    end else begin
      sw_array_0 <= GEN_105;
    end
    if(1'h0) begin
    end else begin
      sw_array_1 <= GEN_106;
    end
    if(1'h0) begin
    end else begin
      sw_array_2 <= GEN_107;
    end
    if(1'h0) begin
    end else begin
      sw_array_3 <= GEN_108;
    end
    if(1'h0) begin
    end else begin
      sw_array_4 <= GEN_109;
    end
    if(1'h0) begin
    end else begin
      sw_array_5 <= GEN_110;
    end
    if(1'h0) begin
    end else begin
      sw_array_6 <= GEN_111;
    end
    if(1'h0) begin
    end else begin
      sw_array_7 <= GEN_112;
    end
    if(1'h0) begin
    end else begin
      sx_array_0 <= GEN_114;
    end
    if(1'h0) begin
    end else begin
      sx_array_1 <= GEN_115;
    end
    if(1'h0) begin
    end else begin
      sx_array_2 <= GEN_116;
    end
    if(1'h0) begin
    end else begin
      sx_array_3 <= GEN_117;
    end
    if(1'h0) begin
    end else begin
      sx_array_4 <= GEN_118;
    end
    if(1'h0) begin
    end else begin
      sx_array_5 <= GEN_119;
    end
    if(1'h0) begin
    end else begin
      sx_array_6 <= GEN_120;
    end
    if(1'h0) begin
    end else begin
      sx_array_7 <= GEN_121;
    end
    if(1'h0) begin
    end else begin
      dirty_array_0 <= GEN_123;
    end
    if(1'h0) begin
    end else begin
      dirty_array_1 <= GEN_124;
    end
    if(1'h0) begin
    end else begin
      dirty_array_2 <= GEN_125;
    end
    if(1'h0) begin
    end else begin
      dirty_array_3 <= GEN_126;
    end
    if(1'h0) begin
    end else begin
      dirty_array_4 <= GEN_127;
    end
    if(1'h0) begin
    end else begin
      dirty_array_5 <= GEN_128;
    end
    if(1'h0) begin
    end else begin
      dirty_array_6 <= GEN_129;
    end
    if(1'h0) begin
    end else begin
      dirty_array_7 <= GEN_130;
    end
    if(1'h0) begin
    end else begin
      T_296 <= GEN_131;
    end
  end
endmodule
module BTB(
  input   clk,
  input   reset,
  input   io_req_valid,
  input  [38:0] io_req_bits_addr,
  output  io_resp_valid,
  output  io_resp_bits_taken,
  output  io_resp_bits_mask,
  output  io_resp_bits_bridx,
  output [38:0] io_resp_bits_target,
  output [5:0] io_resp_bits_entry,
  output [6:0] io_resp_bits_bht_history,
  output [1:0] io_resp_bits_bht_value,
  input   io_btb_update_valid,
  input   io_btb_update_bits_prediction_valid,
  input   io_btb_update_bits_prediction_bits_taken,
  input   io_btb_update_bits_prediction_bits_mask,
  input   io_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_btb_update_bits_prediction_bits_target,
  input  [5:0] io_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_btb_update_bits_pc,
  input  [38:0] io_btb_update_bits_target,
  input   io_btb_update_bits_taken,
  input   io_btb_update_bits_isJump,
  input   io_btb_update_bits_isReturn,
  input  [38:0] io_btb_update_bits_br_pc,
  input   io_bht_update_valid,
  input   io_bht_update_bits_prediction_valid,
  input   io_bht_update_bits_prediction_bits_taken,
  input   io_bht_update_bits_prediction_bits_mask,
  input   io_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_bht_update_bits_prediction_bits_target,
  input  [5:0] io_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_bht_update_bits_pc,
  input   io_bht_update_bits_taken,
  input   io_bht_update_bits_mispredict,
  input   io_ras_update_valid,
  input   io_ras_update_bits_isCall,
  input   io_ras_update_bits_isReturn,
  input  [38:0] io_ras_update_bits_returnAddr,
  input   io_ras_update_bits_prediction_valid,
  input   io_ras_update_bits_prediction_bits_taken,
  input   io_ras_update_bits_prediction_bits_mask,
  input   io_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_ras_update_bits_prediction_bits_target,
  input  [5:0] io_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_ras_update_bits_prediction_bits_bht_value,
  input   io_invalidate
);
  reg [61:0] idxValid;
  reg [63:0] GEN_146;
  reg [11:0] idxs [0:61];
  reg [31:0] GEN_147;
  wire [11:0] idxs_T_1431_data;
  wire [5:0] idxs_T_1431_addr;
  wire  idxs_T_1431_en;
  wire [11:0] idxs_T_1434_data;
  wire [5:0] idxs_T_1434_addr;
  wire  idxs_T_1434_en;
  wire [11:0] idxs_T_1437_data;
  wire [5:0] idxs_T_1437_addr;
  wire  idxs_T_1437_en;
  wire [11:0] idxs_T_1440_data;
  wire [5:0] idxs_T_1440_addr;
  wire  idxs_T_1440_en;
  wire [11:0] idxs_T_1443_data;
  wire [5:0] idxs_T_1443_addr;
  wire  idxs_T_1443_en;
  wire [11:0] idxs_T_1446_data;
  wire [5:0] idxs_T_1446_addr;
  wire  idxs_T_1446_en;
  wire [11:0] idxs_T_1449_data;
  wire [5:0] idxs_T_1449_addr;
  wire  idxs_T_1449_en;
  wire [11:0] idxs_T_1452_data;
  wire [5:0] idxs_T_1452_addr;
  wire  idxs_T_1452_en;
  wire [11:0] idxs_T_1455_data;
  wire [5:0] idxs_T_1455_addr;
  wire  idxs_T_1455_en;
  wire [11:0] idxs_T_1458_data;
  wire [5:0] idxs_T_1458_addr;
  wire  idxs_T_1458_en;
  wire [11:0] idxs_T_1461_data;
  wire [5:0] idxs_T_1461_addr;
  wire  idxs_T_1461_en;
  wire [11:0] idxs_T_1464_data;
  wire [5:0] idxs_T_1464_addr;
  wire  idxs_T_1464_en;
  wire [11:0] idxs_T_1467_data;
  wire [5:0] idxs_T_1467_addr;
  wire  idxs_T_1467_en;
  wire [11:0] idxs_T_1470_data;
  wire [5:0] idxs_T_1470_addr;
  wire  idxs_T_1470_en;
  wire [11:0] idxs_T_1473_data;
  wire [5:0] idxs_T_1473_addr;
  wire  idxs_T_1473_en;
  wire [11:0] idxs_T_1476_data;
  wire [5:0] idxs_T_1476_addr;
  wire  idxs_T_1476_en;
  wire [11:0] idxs_T_1479_data;
  wire [5:0] idxs_T_1479_addr;
  wire  idxs_T_1479_en;
  wire [11:0] idxs_T_1482_data;
  wire [5:0] idxs_T_1482_addr;
  wire  idxs_T_1482_en;
  wire [11:0] idxs_T_1485_data;
  wire [5:0] idxs_T_1485_addr;
  wire  idxs_T_1485_en;
  wire [11:0] idxs_T_1488_data;
  wire [5:0] idxs_T_1488_addr;
  wire  idxs_T_1488_en;
  wire [11:0] idxs_T_1491_data;
  wire [5:0] idxs_T_1491_addr;
  wire  idxs_T_1491_en;
  wire [11:0] idxs_T_1494_data;
  wire [5:0] idxs_T_1494_addr;
  wire  idxs_T_1494_en;
  wire [11:0] idxs_T_1497_data;
  wire [5:0] idxs_T_1497_addr;
  wire  idxs_T_1497_en;
  wire [11:0] idxs_T_1500_data;
  wire [5:0] idxs_T_1500_addr;
  wire  idxs_T_1500_en;
  wire [11:0] idxs_T_1503_data;
  wire [5:0] idxs_T_1503_addr;
  wire  idxs_T_1503_en;
  wire [11:0] idxs_T_1506_data;
  wire [5:0] idxs_T_1506_addr;
  wire  idxs_T_1506_en;
  wire [11:0] idxs_T_1509_data;
  wire [5:0] idxs_T_1509_addr;
  wire  idxs_T_1509_en;
  wire [11:0] idxs_T_1512_data;
  wire [5:0] idxs_T_1512_addr;
  wire  idxs_T_1512_en;
  wire [11:0] idxs_T_1515_data;
  wire [5:0] idxs_T_1515_addr;
  wire  idxs_T_1515_en;
  wire [11:0] idxs_T_1518_data;
  wire [5:0] idxs_T_1518_addr;
  wire  idxs_T_1518_en;
  wire [11:0] idxs_T_1521_data;
  wire [5:0] idxs_T_1521_addr;
  wire  idxs_T_1521_en;
  wire [11:0] idxs_T_1524_data;
  wire [5:0] idxs_T_1524_addr;
  wire  idxs_T_1524_en;
  wire [11:0] idxs_T_1527_data;
  wire [5:0] idxs_T_1527_addr;
  wire  idxs_T_1527_en;
  wire [11:0] idxs_T_1530_data;
  wire [5:0] idxs_T_1530_addr;
  wire  idxs_T_1530_en;
  wire [11:0] idxs_T_1533_data;
  wire [5:0] idxs_T_1533_addr;
  wire  idxs_T_1533_en;
  wire [11:0] idxs_T_1536_data;
  wire [5:0] idxs_T_1536_addr;
  wire  idxs_T_1536_en;
  wire [11:0] idxs_T_1539_data;
  wire [5:0] idxs_T_1539_addr;
  wire  idxs_T_1539_en;
  wire [11:0] idxs_T_1542_data;
  wire [5:0] idxs_T_1542_addr;
  wire  idxs_T_1542_en;
  wire [11:0] idxs_T_1545_data;
  wire [5:0] idxs_T_1545_addr;
  wire  idxs_T_1545_en;
  wire [11:0] idxs_T_1548_data;
  wire [5:0] idxs_T_1548_addr;
  wire  idxs_T_1548_en;
  wire [11:0] idxs_T_1551_data;
  wire [5:0] idxs_T_1551_addr;
  wire  idxs_T_1551_en;
  wire [11:0] idxs_T_1554_data;
  wire [5:0] idxs_T_1554_addr;
  wire  idxs_T_1554_en;
  wire [11:0] idxs_T_1557_data;
  wire [5:0] idxs_T_1557_addr;
  wire  idxs_T_1557_en;
  wire [11:0] idxs_T_1560_data;
  wire [5:0] idxs_T_1560_addr;
  wire  idxs_T_1560_en;
  wire [11:0] idxs_T_1563_data;
  wire [5:0] idxs_T_1563_addr;
  wire  idxs_T_1563_en;
  wire [11:0] idxs_T_1566_data;
  wire [5:0] idxs_T_1566_addr;
  wire  idxs_T_1566_en;
  wire [11:0] idxs_T_1569_data;
  wire [5:0] idxs_T_1569_addr;
  wire  idxs_T_1569_en;
  wire [11:0] idxs_T_1572_data;
  wire [5:0] idxs_T_1572_addr;
  wire  idxs_T_1572_en;
  wire [11:0] idxs_T_1575_data;
  wire [5:0] idxs_T_1575_addr;
  wire  idxs_T_1575_en;
  wire [11:0] idxs_T_1578_data;
  wire [5:0] idxs_T_1578_addr;
  wire  idxs_T_1578_en;
  wire [11:0] idxs_T_1581_data;
  wire [5:0] idxs_T_1581_addr;
  wire  idxs_T_1581_en;
  wire [11:0] idxs_T_1584_data;
  wire [5:0] idxs_T_1584_addr;
  wire  idxs_T_1584_en;
  wire [11:0] idxs_T_1587_data;
  wire [5:0] idxs_T_1587_addr;
  wire  idxs_T_1587_en;
  wire [11:0] idxs_T_1590_data;
  wire [5:0] idxs_T_1590_addr;
  wire  idxs_T_1590_en;
  wire [11:0] idxs_T_1593_data;
  wire [5:0] idxs_T_1593_addr;
  wire  idxs_T_1593_en;
  wire [11:0] idxs_T_1596_data;
  wire [5:0] idxs_T_1596_addr;
  wire  idxs_T_1596_en;
  wire [11:0] idxs_T_1599_data;
  wire [5:0] idxs_T_1599_addr;
  wire  idxs_T_1599_en;
  wire [11:0] idxs_T_1602_data;
  wire [5:0] idxs_T_1602_addr;
  wire  idxs_T_1602_en;
  wire [11:0] idxs_T_1605_data;
  wire [5:0] idxs_T_1605_addr;
  wire  idxs_T_1605_en;
  wire [11:0] idxs_T_1608_data;
  wire [5:0] idxs_T_1608_addr;
  wire  idxs_T_1608_en;
  wire [11:0] idxs_T_1611_data;
  wire [5:0] idxs_T_1611_addr;
  wire  idxs_T_1611_en;
  wire [11:0] idxs_T_1614_data;
  wire [5:0] idxs_T_1614_addr;
  wire  idxs_T_1614_en;
  wire [11:0] idxs_T_1972_data;
  wire [5:0] idxs_T_1972_addr;
  wire  idxs_T_1972_en;
  wire [11:0] idxs_T_1975_data;
  wire [5:0] idxs_T_1975_addr;
  wire  idxs_T_1975_en;
  wire [11:0] idxs_T_1978_data;
  wire [5:0] idxs_T_1978_addr;
  wire  idxs_T_1978_en;
  wire [11:0] idxs_T_1981_data;
  wire [5:0] idxs_T_1981_addr;
  wire  idxs_T_1981_en;
  wire [11:0] idxs_T_1984_data;
  wire [5:0] idxs_T_1984_addr;
  wire  idxs_T_1984_en;
  wire [11:0] idxs_T_1987_data;
  wire [5:0] idxs_T_1987_addr;
  wire  idxs_T_1987_en;
  wire [11:0] idxs_T_1990_data;
  wire [5:0] idxs_T_1990_addr;
  wire  idxs_T_1990_en;
  wire [11:0] idxs_T_1993_data;
  wire [5:0] idxs_T_1993_addr;
  wire  idxs_T_1993_en;
  wire [11:0] idxs_T_1996_data;
  wire [5:0] idxs_T_1996_addr;
  wire  idxs_T_1996_en;
  wire [11:0] idxs_T_1999_data;
  wire [5:0] idxs_T_1999_addr;
  wire  idxs_T_1999_en;
  wire [11:0] idxs_T_2002_data;
  wire [5:0] idxs_T_2002_addr;
  wire  idxs_T_2002_en;
  wire [11:0] idxs_T_2005_data;
  wire [5:0] idxs_T_2005_addr;
  wire  idxs_T_2005_en;
  wire [11:0] idxs_T_2008_data;
  wire [5:0] idxs_T_2008_addr;
  wire  idxs_T_2008_en;
  wire [11:0] idxs_T_2011_data;
  wire [5:0] idxs_T_2011_addr;
  wire  idxs_T_2011_en;
  wire [11:0] idxs_T_2014_data;
  wire [5:0] idxs_T_2014_addr;
  wire  idxs_T_2014_en;
  wire [11:0] idxs_T_2017_data;
  wire [5:0] idxs_T_2017_addr;
  wire  idxs_T_2017_en;
  wire [11:0] idxs_T_2020_data;
  wire [5:0] idxs_T_2020_addr;
  wire  idxs_T_2020_en;
  wire [11:0] idxs_T_2023_data;
  wire [5:0] idxs_T_2023_addr;
  wire  idxs_T_2023_en;
  wire [11:0] idxs_T_2026_data;
  wire [5:0] idxs_T_2026_addr;
  wire  idxs_T_2026_en;
  wire [11:0] idxs_T_2029_data;
  wire [5:0] idxs_T_2029_addr;
  wire  idxs_T_2029_en;
  wire [11:0] idxs_T_2032_data;
  wire [5:0] idxs_T_2032_addr;
  wire  idxs_T_2032_en;
  wire [11:0] idxs_T_2035_data;
  wire [5:0] idxs_T_2035_addr;
  wire  idxs_T_2035_en;
  wire [11:0] idxs_T_2038_data;
  wire [5:0] idxs_T_2038_addr;
  wire  idxs_T_2038_en;
  wire [11:0] idxs_T_2041_data;
  wire [5:0] idxs_T_2041_addr;
  wire  idxs_T_2041_en;
  wire [11:0] idxs_T_2044_data;
  wire [5:0] idxs_T_2044_addr;
  wire  idxs_T_2044_en;
  wire [11:0] idxs_T_2047_data;
  wire [5:0] idxs_T_2047_addr;
  wire  idxs_T_2047_en;
  wire [11:0] idxs_T_2050_data;
  wire [5:0] idxs_T_2050_addr;
  wire  idxs_T_2050_en;
  wire [11:0] idxs_T_2053_data;
  wire [5:0] idxs_T_2053_addr;
  wire  idxs_T_2053_en;
  wire [11:0] idxs_T_2056_data;
  wire [5:0] idxs_T_2056_addr;
  wire  idxs_T_2056_en;
  wire [11:0] idxs_T_2059_data;
  wire [5:0] idxs_T_2059_addr;
  wire  idxs_T_2059_en;
  wire [11:0] idxs_T_2062_data;
  wire [5:0] idxs_T_2062_addr;
  wire  idxs_T_2062_en;
  wire [11:0] idxs_T_2065_data;
  wire [5:0] idxs_T_2065_addr;
  wire  idxs_T_2065_en;
  wire [11:0] idxs_T_2068_data;
  wire [5:0] idxs_T_2068_addr;
  wire  idxs_T_2068_en;
  wire [11:0] idxs_T_2071_data;
  wire [5:0] idxs_T_2071_addr;
  wire  idxs_T_2071_en;
  wire [11:0] idxs_T_2074_data;
  wire [5:0] idxs_T_2074_addr;
  wire  idxs_T_2074_en;
  wire [11:0] idxs_T_2077_data;
  wire [5:0] idxs_T_2077_addr;
  wire  idxs_T_2077_en;
  wire [11:0] idxs_T_2080_data;
  wire [5:0] idxs_T_2080_addr;
  wire  idxs_T_2080_en;
  wire [11:0] idxs_T_2083_data;
  wire [5:0] idxs_T_2083_addr;
  wire  idxs_T_2083_en;
  wire [11:0] idxs_T_2086_data;
  wire [5:0] idxs_T_2086_addr;
  wire  idxs_T_2086_en;
  wire [11:0] idxs_T_2089_data;
  wire [5:0] idxs_T_2089_addr;
  wire  idxs_T_2089_en;
  wire [11:0] idxs_T_2092_data;
  wire [5:0] idxs_T_2092_addr;
  wire  idxs_T_2092_en;
  wire [11:0] idxs_T_2095_data;
  wire [5:0] idxs_T_2095_addr;
  wire  idxs_T_2095_en;
  wire [11:0] idxs_T_2098_data;
  wire [5:0] idxs_T_2098_addr;
  wire  idxs_T_2098_en;
  wire [11:0] idxs_T_2101_data;
  wire [5:0] idxs_T_2101_addr;
  wire  idxs_T_2101_en;
  wire [11:0] idxs_T_2104_data;
  wire [5:0] idxs_T_2104_addr;
  wire  idxs_T_2104_en;
  wire [11:0] idxs_T_2107_data;
  wire [5:0] idxs_T_2107_addr;
  wire  idxs_T_2107_en;
  wire [11:0] idxs_T_2110_data;
  wire [5:0] idxs_T_2110_addr;
  wire  idxs_T_2110_en;
  wire [11:0] idxs_T_2113_data;
  wire [5:0] idxs_T_2113_addr;
  wire  idxs_T_2113_en;
  wire [11:0] idxs_T_2116_data;
  wire [5:0] idxs_T_2116_addr;
  wire  idxs_T_2116_en;
  wire [11:0] idxs_T_2119_data;
  wire [5:0] idxs_T_2119_addr;
  wire  idxs_T_2119_en;
  wire [11:0] idxs_T_2122_data;
  wire [5:0] idxs_T_2122_addr;
  wire  idxs_T_2122_en;
  wire [11:0] idxs_T_2125_data;
  wire [5:0] idxs_T_2125_addr;
  wire  idxs_T_2125_en;
  wire [11:0] idxs_T_2128_data;
  wire [5:0] idxs_T_2128_addr;
  wire  idxs_T_2128_en;
  wire [11:0] idxs_T_2131_data;
  wire [5:0] idxs_T_2131_addr;
  wire  idxs_T_2131_en;
  wire [11:0] idxs_T_2134_data;
  wire [5:0] idxs_T_2134_addr;
  wire  idxs_T_2134_en;
  wire [11:0] idxs_T_2137_data;
  wire [5:0] idxs_T_2137_addr;
  wire  idxs_T_2137_en;
  wire [11:0] idxs_T_2140_data;
  wire [5:0] idxs_T_2140_addr;
  wire  idxs_T_2140_en;
  wire [11:0] idxs_T_2143_data;
  wire [5:0] idxs_T_2143_addr;
  wire  idxs_T_2143_en;
  wire [11:0] idxs_T_2146_data;
  wire [5:0] idxs_T_2146_addr;
  wire  idxs_T_2146_en;
  wire [11:0] idxs_T_2149_data;
  wire [5:0] idxs_T_2149_addr;
  wire  idxs_T_2149_en;
  wire [11:0] idxs_T_2152_data;
  wire [5:0] idxs_T_2152_addr;
  wire  idxs_T_2152_en;
  wire [11:0] idxs_T_2155_data;
  wire [5:0] idxs_T_2155_addr;
  wire  idxs_T_2155_en;
  wire [11:0] idxs_T_2872_data;
  wire [5:0] idxs_T_2872_addr;
  wire  idxs_T_2872_mask;
  wire  idxs_T_2872_en;
  reg [2:0] idxPages [0:61];
  reg [31:0] GEN_148;
  wire [2:0] idxPages_T_578_data;
  wire [5:0] idxPages_T_578_addr;
  wire  idxPages_T_578_en;
  wire [2:0] idxPages_T_583_data;
  wire [5:0] idxPages_T_583_addr;
  wire  idxPages_T_583_en;
  wire [2:0] idxPages_T_588_data;
  wire [5:0] idxPages_T_588_addr;
  wire  idxPages_T_588_en;
  wire [2:0] idxPages_T_593_data;
  wire [5:0] idxPages_T_593_addr;
  wire  idxPages_T_593_en;
  wire [2:0] idxPages_T_598_data;
  wire [5:0] idxPages_T_598_addr;
  wire  idxPages_T_598_en;
  wire [2:0] idxPages_T_603_data;
  wire [5:0] idxPages_T_603_addr;
  wire  idxPages_T_603_en;
  wire [2:0] idxPages_T_608_data;
  wire [5:0] idxPages_T_608_addr;
  wire  idxPages_T_608_en;
  wire [2:0] idxPages_T_613_data;
  wire [5:0] idxPages_T_613_addr;
  wire  idxPages_T_613_en;
  wire [2:0] idxPages_T_618_data;
  wire [5:0] idxPages_T_618_addr;
  wire  idxPages_T_618_en;
  wire [2:0] idxPages_T_623_data;
  wire [5:0] idxPages_T_623_addr;
  wire  idxPages_T_623_en;
  wire [2:0] idxPages_T_628_data;
  wire [5:0] idxPages_T_628_addr;
  wire  idxPages_T_628_en;
  wire [2:0] idxPages_T_633_data;
  wire [5:0] idxPages_T_633_addr;
  wire  idxPages_T_633_en;
  wire [2:0] idxPages_T_638_data;
  wire [5:0] idxPages_T_638_addr;
  wire  idxPages_T_638_en;
  wire [2:0] idxPages_T_643_data;
  wire [5:0] idxPages_T_643_addr;
  wire  idxPages_T_643_en;
  wire [2:0] idxPages_T_648_data;
  wire [5:0] idxPages_T_648_addr;
  wire  idxPages_T_648_en;
  wire [2:0] idxPages_T_653_data;
  wire [5:0] idxPages_T_653_addr;
  wire  idxPages_T_653_en;
  wire [2:0] idxPages_T_658_data;
  wire [5:0] idxPages_T_658_addr;
  wire  idxPages_T_658_en;
  wire [2:0] idxPages_T_663_data;
  wire [5:0] idxPages_T_663_addr;
  wire  idxPages_T_663_en;
  wire [2:0] idxPages_T_668_data;
  wire [5:0] idxPages_T_668_addr;
  wire  idxPages_T_668_en;
  wire [2:0] idxPages_T_673_data;
  wire [5:0] idxPages_T_673_addr;
  wire  idxPages_T_673_en;
  wire [2:0] idxPages_T_678_data;
  wire [5:0] idxPages_T_678_addr;
  wire  idxPages_T_678_en;
  wire [2:0] idxPages_T_683_data;
  wire [5:0] idxPages_T_683_addr;
  wire  idxPages_T_683_en;
  wire [2:0] idxPages_T_688_data;
  wire [5:0] idxPages_T_688_addr;
  wire  idxPages_T_688_en;
  wire [2:0] idxPages_T_693_data;
  wire [5:0] idxPages_T_693_addr;
  wire  idxPages_T_693_en;
  wire [2:0] idxPages_T_698_data;
  wire [5:0] idxPages_T_698_addr;
  wire  idxPages_T_698_en;
  wire [2:0] idxPages_T_703_data;
  wire [5:0] idxPages_T_703_addr;
  wire  idxPages_T_703_en;
  wire [2:0] idxPages_T_708_data;
  wire [5:0] idxPages_T_708_addr;
  wire  idxPages_T_708_en;
  wire [2:0] idxPages_T_713_data;
  wire [5:0] idxPages_T_713_addr;
  wire  idxPages_T_713_en;
  wire [2:0] idxPages_T_718_data;
  wire [5:0] idxPages_T_718_addr;
  wire  idxPages_T_718_en;
  wire [2:0] idxPages_T_723_data;
  wire [5:0] idxPages_T_723_addr;
  wire  idxPages_T_723_en;
  wire [2:0] idxPages_T_728_data;
  wire [5:0] idxPages_T_728_addr;
  wire  idxPages_T_728_en;
  wire [2:0] idxPages_T_733_data;
  wire [5:0] idxPages_T_733_addr;
  wire  idxPages_T_733_en;
  wire [2:0] idxPages_T_738_data;
  wire [5:0] idxPages_T_738_addr;
  wire  idxPages_T_738_en;
  wire [2:0] idxPages_T_743_data;
  wire [5:0] idxPages_T_743_addr;
  wire  idxPages_T_743_en;
  wire [2:0] idxPages_T_748_data;
  wire [5:0] idxPages_T_748_addr;
  wire  idxPages_T_748_en;
  wire [2:0] idxPages_T_753_data;
  wire [5:0] idxPages_T_753_addr;
  wire  idxPages_T_753_en;
  wire [2:0] idxPages_T_758_data;
  wire [5:0] idxPages_T_758_addr;
  wire  idxPages_T_758_en;
  wire [2:0] idxPages_T_763_data;
  wire [5:0] idxPages_T_763_addr;
  wire  idxPages_T_763_en;
  wire [2:0] idxPages_T_768_data;
  wire [5:0] idxPages_T_768_addr;
  wire  idxPages_T_768_en;
  wire [2:0] idxPages_T_773_data;
  wire [5:0] idxPages_T_773_addr;
  wire  idxPages_T_773_en;
  wire [2:0] idxPages_T_778_data;
  wire [5:0] idxPages_T_778_addr;
  wire  idxPages_T_778_en;
  wire [2:0] idxPages_T_783_data;
  wire [5:0] idxPages_T_783_addr;
  wire  idxPages_T_783_en;
  wire [2:0] idxPages_T_788_data;
  wire [5:0] idxPages_T_788_addr;
  wire  idxPages_T_788_en;
  wire [2:0] idxPages_T_793_data;
  wire [5:0] idxPages_T_793_addr;
  wire  idxPages_T_793_en;
  wire [2:0] idxPages_T_798_data;
  wire [5:0] idxPages_T_798_addr;
  wire  idxPages_T_798_en;
  wire [2:0] idxPages_T_803_data;
  wire [5:0] idxPages_T_803_addr;
  wire  idxPages_T_803_en;
  wire [2:0] idxPages_T_808_data;
  wire [5:0] idxPages_T_808_addr;
  wire  idxPages_T_808_en;
  wire [2:0] idxPages_T_813_data;
  wire [5:0] idxPages_T_813_addr;
  wire  idxPages_T_813_en;
  wire [2:0] idxPages_T_818_data;
  wire [5:0] idxPages_T_818_addr;
  wire  idxPages_T_818_en;
  wire [2:0] idxPages_T_823_data;
  wire [5:0] idxPages_T_823_addr;
  wire  idxPages_T_823_en;
  wire [2:0] idxPages_T_828_data;
  wire [5:0] idxPages_T_828_addr;
  wire  idxPages_T_828_en;
  wire [2:0] idxPages_T_833_data;
  wire [5:0] idxPages_T_833_addr;
  wire  idxPages_T_833_en;
  wire [2:0] idxPages_T_838_data;
  wire [5:0] idxPages_T_838_addr;
  wire  idxPages_T_838_en;
  wire [2:0] idxPages_T_843_data;
  wire [5:0] idxPages_T_843_addr;
  wire  idxPages_T_843_en;
  wire [2:0] idxPages_T_848_data;
  wire [5:0] idxPages_T_848_addr;
  wire  idxPages_T_848_en;
  wire [2:0] idxPages_T_853_data;
  wire [5:0] idxPages_T_853_addr;
  wire  idxPages_T_853_en;
  wire [2:0] idxPages_T_858_data;
  wire [5:0] idxPages_T_858_addr;
  wire  idxPages_T_858_en;
  wire [2:0] idxPages_T_863_data;
  wire [5:0] idxPages_T_863_addr;
  wire  idxPages_T_863_en;
  wire [2:0] idxPages_T_868_data;
  wire [5:0] idxPages_T_868_addr;
  wire  idxPages_T_868_en;
  wire [2:0] idxPages_T_873_data;
  wire [5:0] idxPages_T_873_addr;
  wire  idxPages_T_873_en;
  wire [2:0] idxPages_T_878_data;
  wire [5:0] idxPages_T_878_addr;
  wire  idxPages_T_878_en;
  wire [2:0] idxPages_T_883_data;
  wire [5:0] idxPages_T_883_addr;
  wire  idxPages_T_883_en;
  wire [2:0] idxPages_T_2874_data;
  wire [5:0] idxPages_T_2874_addr;
  wire  idxPages_T_2874_mask;
  wire  idxPages_T_2874_en;
  reg [11:0] tgts [0:61];
  reg [31:0] GEN_149;
  wire [11:0] tgts_T_3270_data;
  wire [5:0] tgts_T_3270_addr;
  wire  tgts_T_3270_en;
  wire [11:0] tgts_T_3272_data;
  wire [5:0] tgts_T_3272_addr;
  wire  tgts_T_3272_en;
  wire [11:0] tgts_T_3274_data;
  wire [5:0] tgts_T_3274_addr;
  wire  tgts_T_3274_en;
  wire [11:0] tgts_T_3276_data;
  wire [5:0] tgts_T_3276_addr;
  wire  tgts_T_3276_en;
  wire [11:0] tgts_T_3278_data;
  wire [5:0] tgts_T_3278_addr;
  wire  tgts_T_3278_en;
  wire [11:0] tgts_T_3280_data;
  wire [5:0] tgts_T_3280_addr;
  wire  tgts_T_3280_en;
  wire [11:0] tgts_T_3282_data;
  wire [5:0] tgts_T_3282_addr;
  wire  tgts_T_3282_en;
  wire [11:0] tgts_T_3284_data;
  wire [5:0] tgts_T_3284_addr;
  wire  tgts_T_3284_en;
  wire [11:0] tgts_T_3286_data;
  wire [5:0] tgts_T_3286_addr;
  wire  tgts_T_3286_en;
  wire [11:0] tgts_T_3288_data;
  wire [5:0] tgts_T_3288_addr;
  wire  tgts_T_3288_en;
  wire [11:0] tgts_T_3290_data;
  wire [5:0] tgts_T_3290_addr;
  wire  tgts_T_3290_en;
  wire [11:0] tgts_T_3292_data;
  wire [5:0] tgts_T_3292_addr;
  wire  tgts_T_3292_en;
  wire [11:0] tgts_T_3294_data;
  wire [5:0] tgts_T_3294_addr;
  wire  tgts_T_3294_en;
  wire [11:0] tgts_T_3296_data;
  wire [5:0] tgts_T_3296_addr;
  wire  tgts_T_3296_en;
  wire [11:0] tgts_T_3298_data;
  wire [5:0] tgts_T_3298_addr;
  wire  tgts_T_3298_en;
  wire [11:0] tgts_T_3300_data;
  wire [5:0] tgts_T_3300_addr;
  wire  tgts_T_3300_en;
  wire [11:0] tgts_T_3302_data;
  wire [5:0] tgts_T_3302_addr;
  wire  tgts_T_3302_en;
  wire [11:0] tgts_T_3304_data;
  wire [5:0] tgts_T_3304_addr;
  wire  tgts_T_3304_en;
  wire [11:0] tgts_T_3306_data;
  wire [5:0] tgts_T_3306_addr;
  wire  tgts_T_3306_en;
  wire [11:0] tgts_T_3308_data;
  wire [5:0] tgts_T_3308_addr;
  wire  tgts_T_3308_en;
  wire [11:0] tgts_T_3310_data;
  wire [5:0] tgts_T_3310_addr;
  wire  tgts_T_3310_en;
  wire [11:0] tgts_T_3312_data;
  wire [5:0] tgts_T_3312_addr;
  wire  tgts_T_3312_en;
  wire [11:0] tgts_T_3314_data;
  wire [5:0] tgts_T_3314_addr;
  wire  tgts_T_3314_en;
  wire [11:0] tgts_T_3316_data;
  wire [5:0] tgts_T_3316_addr;
  wire  tgts_T_3316_en;
  wire [11:0] tgts_T_3318_data;
  wire [5:0] tgts_T_3318_addr;
  wire  tgts_T_3318_en;
  wire [11:0] tgts_T_3320_data;
  wire [5:0] tgts_T_3320_addr;
  wire  tgts_T_3320_en;
  wire [11:0] tgts_T_3322_data;
  wire [5:0] tgts_T_3322_addr;
  wire  tgts_T_3322_en;
  wire [11:0] tgts_T_3324_data;
  wire [5:0] tgts_T_3324_addr;
  wire  tgts_T_3324_en;
  wire [11:0] tgts_T_3326_data;
  wire [5:0] tgts_T_3326_addr;
  wire  tgts_T_3326_en;
  wire [11:0] tgts_T_3328_data;
  wire [5:0] tgts_T_3328_addr;
  wire  tgts_T_3328_en;
  wire [11:0] tgts_T_3330_data;
  wire [5:0] tgts_T_3330_addr;
  wire  tgts_T_3330_en;
  wire [11:0] tgts_T_3332_data;
  wire [5:0] tgts_T_3332_addr;
  wire  tgts_T_3332_en;
  wire [11:0] tgts_T_3334_data;
  wire [5:0] tgts_T_3334_addr;
  wire  tgts_T_3334_en;
  wire [11:0] tgts_T_3336_data;
  wire [5:0] tgts_T_3336_addr;
  wire  tgts_T_3336_en;
  wire [11:0] tgts_T_3338_data;
  wire [5:0] tgts_T_3338_addr;
  wire  tgts_T_3338_en;
  wire [11:0] tgts_T_3340_data;
  wire [5:0] tgts_T_3340_addr;
  wire  tgts_T_3340_en;
  wire [11:0] tgts_T_3342_data;
  wire [5:0] tgts_T_3342_addr;
  wire  tgts_T_3342_en;
  wire [11:0] tgts_T_3344_data;
  wire [5:0] tgts_T_3344_addr;
  wire  tgts_T_3344_en;
  wire [11:0] tgts_T_3346_data;
  wire [5:0] tgts_T_3346_addr;
  wire  tgts_T_3346_en;
  wire [11:0] tgts_T_3348_data;
  wire [5:0] tgts_T_3348_addr;
  wire  tgts_T_3348_en;
  wire [11:0] tgts_T_3350_data;
  wire [5:0] tgts_T_3350_addr;
  wire  tgts_T_3350_en;
  wire [11:0] tgts_T_3352_data;
  wire [5:0] tgts_T_3352_addr;
  wire  tgts_T_3352_en;
  wire [11:0] tgts_T_3354_data;
  wire [5:0] tgts_T_3354_addr;
  wire  tgts_T_3354_en;
  wire [11:0] tgts_T_3356_data;
  wire [5:0] tgts_T_3356_addr;
  wire  tgts_T_3356_en;
  wire [11:0] tgts_T_3358_data;
  wire [5:0] tgts_T_3358_addr;
  wire  tgts_T_3358_en;
  wire [11:0] tgts_T_3360_data;
  wire [5:0] tgts_T_3360_addr;
  wire  tgts_T_3360_en;
  wire [11:0] tgts_T_3362_data;
  wire [5:0] tgts_T_3362_addr;
  wire  tgts_T_3362_en;
  wire [11:0] tgts_T_3364_data;
  wire [5:0] tgts_T_3364_addr;
  wire  tgts_T_3364_en;
  wire [11:0] tgts_T_3366_data;
  wire [5:0] tgts_T_3366_addr;
  wire  tgts_T_3366_en;
  wire [11:0] tgts_T_3368_data;
  wire [5:0] tgts_T_3368_addr;
  wire  tgts_T_3368_en;
  wire [11:0] tgts_T_3370_data;
  wire [5:0] tgts_T_3370_addr;
  wire  tgts_T_3370_en;
  wire [11:0] tgts_T_3372_data;
  wire [5:0] tgts_T_3372_addr;
  wire  tgts_T_3372_en;
  wire [11:0] tgts_T_3374_data;
  wire [5:0] tgts_T_3374_addr;
  wire  tgts_T_3374_en;
  wire [11:0] tgts_T_3376_data;
  wire [5:0] tgts_T_3376_addr;
  wire  tgts_T_3376_en;
  wire [11:0] tgts_T_3378_data;
  wire [5:0] tgts_T_3378_addr;
  wire  tgts_T_3378_en;
  wire [11:0] tgts_T_3380_data;
  wire [5:0] tgts_T_3380_addr;
  wire  tgts_T_3380_en;
  wire [11:0] tgts_T_3382_data;
  wire [5:0] tgts_T_3382_addr;
  wire  tgts_T_3382_en;
  wire [11:0] tgts_T_3384_data;
  wire [5:0] tgts_T_3384_addr;
  wire  tgts_T_3384_en;
  wire [11:0] tgts_T_3386_data;
  wire [5:0] tgts_T_3386_addr;
  wire  tgts_T_3386_en;
  wire [11:0] tgts_T_3388_data;
  wire [5:0] tgts_T_3388_addr;
  wire  tgts_T_3388_en;
  wire [11:0] tgts_T_3390_data;
  wire [5:0] tgts_T_3390_addr;
  wire  tgts_T_3390_en;
  wire [11:0] tgts_T_3392_data;
  wire [5:0] tgts_T_3392_addr;
  wire  tgts_T_3392_en;
  wire [11:0] tgts_T_2873_data;
  wire [5:0] tgts_T_2873_addr;
  wire  tgts_T_2873_mask;
  wire  tgts_T_2873_en;
  reg [2:0] tgtPages [0:61];
  reg [31:0] GEN_150;
  wire [2:0] tgtPages_T_888_data;
  wire [5:0] tgtPages_T_888_addr;
  wire  tgtPages_T_888_en;
  wire [2:0] tgtPages_T_893_data;
  wire [5:0] tgtPages_T_893_addr;
  wire  tgtPages_T_893_en;
  wire [2:0] tgtPages_T_898_data;
  wire [5:0] tgtPages_T_898_addr;
  wire  tgtPages_T_898_en;
  wire [2:0] tgtPages_T_903_data;
  wire [5:0] tgtPages_T_903_addr;
  wire  tgtPages_T_903_en;
  wire [2:0] tgtPages_T_908_data;
  wire [5:0] tgtPages_T_908_addr;
  wire  tgtPages_T_908_en;
  wire [2:0] tgtPages_T_913_data;
  wire [5:0] tgtPages_T_913_addr;
  wire  tgtPages_T_913_en;
  wire [2:0] tgtPages_T_918_data;
  wire [5:0] tgtPages_T_918_addr;
  wire  tgtPages_T_918_en;
  wire [2:0] tgtPages_T_923_data;
  wire [5:0] tgtPages_T_923_addr;
  wire  tgtPages_T_923_en;
  wire [2:0] tgtPages_T_928_data;
  wire [5:0] tgtPages_T_928_addr;
  wire  tgtPages_T_928_en;
  wire [2:0] tgtPages_T_933_data;
  wire [5:0] tgtPages_T_933_addr;
  wire  tgtPages_T_933_en;
  wire [2:0] tgtPages_T_938_data;
  wire [5:0] tgtPages_T_938_addr;
  wire  tgtPages_T_938_en;
  wire [2:0] tgtPages_T_943_data;
  wire [5:0] tgtPages_T_943_addr;
  wire  tgtPages_T_943_en;
  wire [2:0] tgtPages_T_948_data;
  wire [5:0] tgtPages_T_948_addr;
  wire  tgtPages_T_948_en;
  wire [2:0] tgtPages_T_953_data;
  wire [5:0] tgtPages_T_953_addr;
  wire  tgtPages_T_953_en;
  wire [2:0] tgtPages_T_958_data;
  wire [5:0] tgtPages_T_958_addr;
  wire  tgtPages_T_958_en;
  wire [2:0] tgtPages_T_963_data;
  wire [5:0] tgtPages_T_963_addr;
  wire  tgtPages_T_963_en;
  wire [2:0] tgtPages_T_968_data;
  wire [5:0] tgtPages_T_968_addr;
  wire  tgtPages_T_968_en;
  wire [2:0] tgtPages_T_973_data;
  wire [5:0] tgtPages_T_973_addr;
  wire  tgtPages_T_973_en;
  wire [2:0] tgtPages_T_978_data;
  wire [5:0] tgtPages_T_978_addr;
  wire  tgtPages_T_978_en;
  wire [2:0] tgtPages_T_983_data;
  wire [5:0] tgtPages_T_983_addr;
  wire  tgtPages_T_983_en;
  wire [2:0] tgtPages_T_988_data;
  wire [5:0] tgtPages_T_988_addr;
  wire  tgtPages_T_988_en;
  wire [2:0] tgtPages_T_993_data;
  wire [5:0] tgtPages_T_993_addr;
  wire  tgtPages_T_993_en;
  wire [2:0] tgtPages_T_998_data;
  wire [5:0] tgtPages_T_998_addr;
  wire  tgtPages_T_998_en;
  wire [2:0] tgtPages_T_1003_data;
  wire [5:0] tgtPages_T_1003_addr;
  wire  tgtPages_T_1003_en;
  wire [2:0] tgtPages_T_1008_data;
  wire [5:0] tgtPages_T_1008_addr;
  wire  tgtPages_T_1008_en;
  wire [2:0] tgtPages_T_1013_data;
  wire [5:0] tgtPages_T_1013_addr;
  wire  tgtPages_T_1013_en;
  wire [2:0] tgtPages_T_1018_data;
  wire [5:0] tgtPages_T_1018_addr;
  wire  tgtPages_T_1018_en;
  wire [2:0] tgtPages_T_1023_data;
  wire [5:0] tgtPages_T_1023_addr;
  wire  tgtPages_T_1023_en;
  wire [2:0] tgtPages_T_1028_data;
  wire [5:0] tgtPages_T_1028_addr;
  wire  tgtPages_T_1028_en;
  wire [2:0] tgtPages_T_1033_data;
  wire [5:0] tgtPages_T_1033_addr;
  wire  tgtPages_T_1033_en;
  wire [2:0] tgtPages_T_1038_data;
  wire [5:0] tgtPages_T_1038_addr;
  wire  tgtPages_T_1038_en;
  wire [2:0] tgtPages_T_1043_data;
  wire [5:0] tgtPages_T_1043_addr;
  wire  tgtPages_T_1043_en;
  wire [2:0] tgtPages_T_1048_data;
  wire [5:0] tgtPages_T_1048_addr;
  wire  tgtPages_T_1048_en;
  wire [2:0] tgtPages_T_1053_data;
  wire [5:0] tgtPages_T_1053_addr;
  wire  tgtPages_T_1053_en;
  wire [2:0] tgtPages_T_1058_data;
  wire [5:0] tgtPages_T_1058_addr;
  wire  tgtPages_T_1058_en;
  wire [2:0] tgtPages_T_1063_data;
  wire [5:0] tgtPages_T_1063_addr;
  wire  tgtPages_T_1063_en;
  wire [2:0] tgtPages_T_1068_data;
  wire [5:0] tgtPages_T_1068_addr;
  wire  tgtPages_T_1068_en;
  wire [2:0] tgtPages_T_1073_data;
  wire [5:0] tgtPages_T_1073_addr;
  wire  tgtPages_T_1073_en;
  wire [2:0] tgtPages_T_1078_data;
  wire [5:0] tgtPages_T_1078_addr;
  wire  tgtPages_T_1078_en;
  wire [2:0] tgtPages_T_1083_data;
  wire [5:0] tgtPages_T_1083_addr;
  wire  tgtPages_T_1083_en;
  wire [2:0] tgtPages_T_1088_data;
  wire [5:0] tgtPages_T_1088_addr;
  wire  tgtPages_T_1088_en;
  wire [2:0] tgtPages_T_1093_data;
  wire [5:0] tgtPages_T_1093_addr;
  wire  tgtPages_T_1093_en;
  wire [2:0] tgtPages_T_1098_data;
  wire [5:0] tgtPages_T_1098_addr;
  wire  tgtPages_T_1098_en;
  wire [2:0] tgtPages_T_1103_data;
  wire [5:0] tgtPages_T_1103_addr;
  wire  tgtPages_T_1103_en;
  wire [2:0] tgtPages_T_1108_data;
  wire [5:0] tgtPages_T_1108_addr;
  wire  tgtPages_T_1108_en;
  wire [2:0] tgtPages_T_1113_data;
  wire [5:0] tgtPages_T_1113_addr;
  wire  tgtPages_T_1113_en;
  wire [2:0] tgtPages_T_1118_data;
  wire [5:0] tgtPages_T_1118_addr;
  wire  tgtPages_T_1118_en;
  wire [2:0] tgtPages_T_1123_data;
  wire [5:0] tgtPages_T_1123_addr;
  wire  tgtPages_T_1123_en;
  wire [2:0] tgtPages_T_1128_data;
  wire [5:0] tgtPages_T_1128_addr;
  wire  tgtPages_T_1128_en;
  wire [2:0] tgtPages_T_1133_data;
  wire [5:0] tgtPages_T_1133_addr;
  wire  tgtPages_T_1133_en;
  wire [2:0] tgtPages_T_1138_data;
  wire [5:0] tgtPages_T_1138_addr;
  wire  tgtPages_T_1138_en;
  wire [2:0] tgtPages_T_1143_data;
  wire [5:0] tgtPages_T_1143_addr;
  wire  tgtPages_T_1143_en;
  wire [2:0] tgtPages_T_1148_data;
  wire [5:0] tgtPages_T_1148_addr;
  wire  tgtPages_T_1148_en;
  wire [2:0] tgtPages_T_1153_data;
  wire [5:0] tgtPages_T_1153_addr;
  wire  tgtPages_T_1153_en;
  wire [2:0] tgtPages_T_1158_data;
  wire [5:0] tgtPages_T_1158_addr;
  wire  tgtPages_T_1158_en;
  wire [2:0] tgtPages_T_1163_data;
  wire [5:0] tgtPages_T_1163_addr;
  wire  tgtPages_T_1163_en;
  wire [2:0] tgtPages_T_1168_data;
  wire [5:0] tgtPages_T_1168_addr;
  wire  tgtPages_T_1168_en;
  wire [2:0] tgtPages_T_1173_data;
  wire [5:0] tgtPages_T_1173_addr;
  wire  tgtPages_T_1173_en;
  wire [2:0] tgtPages_T_1178_data;
  wire [5:0] tgtPages_T_1178_addr;
  wire  tgtPages_T_1178_en;
  wire [2:0] tgtPages_T_1183_data;
  wire [5:0] tgtPages_T_1183_addr;
  wire  tgtPages_T_1183_en;
  wire [2:0] tgtPages_T_1188_data;
  wire [5:0] tgtPages_T_1188_addr;
  wire  tgtPages_T_1188_en;
  wire [2:0] tgtPages_T_1193_data;
  wire [5:0] tgtPages_T_1193_addr;
  wire  tgtPages_T_1193_en;
  wire [2:0] tgtPages_T_2875_data;
  wire [5:0] tgtPages_T_2875_addr;
  wire  tgtPages_T_2875_mask;
  wire  tgtPages_T_2875_en;
  reg [26:0] pages [0:5];
  reg [31:0] GEN_151;
  wire [26:0] pages_T_1400_data;
  wire [2:0] pages_T_1400_addr;
  wire  pages_T_1400_en;
  wire [26:0] pages_T_1403_data;
  wire [2:0] pages_T_1403_addr;
  wire  pages_T_1403_en;
  wire [26:0] pages_T_1406_data;
  wire [2:0] pages_T_1406_addr;
  wire  pages_T_1406_en;
  wire [26:0] pages_T_1409_data;
  wire [2:0] pages_T_1409_addr;
  wire  pages_T_1409_en;
  wire [26:0] pages_T_1412_data;
  wire [2:0] pages_T_1412_addr;
  wire  pages_T_1412_en;
  wire [26:0] pages_T_1415_data;
  wire [2:0] pages_T_1415_addr;
  wire  pages_T_1415_en;
  wire [26:0] pages_T_1941_data;
  wire [2:0] pages_T_1941_addr;
  wire  pages_T_1941_en;
  wire [26:0] pages_T_1944_data;
  wire [2:0] pages_T_1944_addr;
  wire  pages_T_1944_en;
  wire [26:0] pages_T_1947_data;
  wire [2:0] pages_T_1947_addr;
  wire  pages_T_1947_en;
  wire [26:0] pages_T_1950_data;
  wire [2:0] pages_T_1950_addr;
  wire  pages_T_1950_en;
  wire [26:0] pages_T_1953_data;
  wire [2:0] pages_T_1953_addr;
  wire  pages_T_1953_en;
  wire [26:0] pages_T_1956_data;
  wire [2:0] pages_T_1956_addr;
  wire  pages_T_1956_en;
  wire [26:0] pages_T_3177_data;
  wire [2:0] pages_T_3177_addr;
  wire  pages_T_3177_en;
  wire [26:0] pages_T_3179_data;
  wire [2:0] pages_T_3179_addr;
  wire  pages_T_3179_en;
  wire [26:0] pages_T_3181_data;
  wire [2:0] pages_T_3181_addr;
  wire  pages_T_3181_en;
  wire [26:0] pages_T_3183_data;
  wire [2:0] pages_T_3183_addr;
  wire  pages_T_3183_en;
  wire [26:0] pages_T_3185_data;
  wire [2:0] pages_T_3185_addr;
  wire  pages_T_3185_en;
  wire [26:0] pages_T_3187_data;
  wire [2:0] pages_T_3187_addr;
  wire  pages_T_3187_en;
  wire [26:0] pages_T_2891_data;
  wire [2:0] pages_T_2891_addr;
  wire  pages_T_2891_mask;
  wire  pages_T_2891_en;
  wire [26:0] pages_T_2895_data;
  wire [2:0] pages_T_2895_addr;
  wire  pages_T_2895_mask;
  wire  pages_T_2895_en;
  wire [26:0] pages_T_2899_data;
  wire [2:0] pages_T_2899_addr;
  wire  pages_T_2899_mask;
  wire  pages_T_2899_en;
  wire [26:0] pages_T_2907_data;
  wire [2:0] pages_T_2907_addr;
  wire  pages_T_2907_mask;
  wire  pages_T_2907_en;
  wire [26:0] pages_T_2911_data;
  wire [2:0] pages_T_2911_addr;
  wire  pages_T_2911_mask;
  wire  pages_T_2911_en;
  wire [26:0] pages_T_2915_data;
  wire [2:0] pages_T_2915_addr;
  wire  pages_T_2915_mask;
  wire  pages_T_2915_en;
  reg [5:0] pageValid;
  reg [31:0] GEN_152;
  wire [7:0] GEN_457;
  wire [7:0] T_580;
  wire [5:0] T_581;
  wire [7:0] T_585;
  wire [5:0] T_586;
  wire [7:0] T_590;
  wire [5:0] T_591;
  wire [7:0] T_595;
  wire [5:0] T_596;
  wire [7:0] T_600;
  wire [5:0] T_601;
  wire [7:0] T_605;
  wire [5:0] T_606;
  wire [7:0] T_610;
  wire [5:0] T_611;
  wire [7:0] T_615;
  wire [5:0] T_616;
  wire [7:0] T_620;
  wire [5:0] T_621;
  wire [7:0] T_625;
  wire [5:0] T_626;
  wire [7:0] T_630;
  wire [5:0] T_631;
  wire [7:0] T_635;
  wire [5:0] T_636;
  wire [7:0] T_640;
  wire [5:0] T_641;
  wire [7:0] T_645;
  wire [5:0] T_646;
  wire [7:0] T_650;
  wire [5:0] T_651;
  wire [7:0] T_655;
  wire [5:0] T_656;
  wire [7:0] T_660;
  wire [5:0] T_661;
  wire [7:0] T_665;
  wire [5:0] T_666;
  wire [7:0] T_670;
  wire [5:0] T_671;
  wire [7:0] T_675;
  wire [5:0] T_676;
  wire [7:0] T_680;
  wire [5:0] T_681;
  wire [7:0] T_685;
  wire [5:0] T_686;
  wire [7:0] T_690;
  wire [5:0] T_691;
  wire [7:0] T_695;
  wire [5:0] T_696;
  wire [7:0] T_700;
  wire [5:0] T_701;
  wire [7:0] T_705;
  wire [5:0] T_706;
  wire [7:0] T_710;
  wire [5:0] T_711;
  wire [7:0] T_715;
  wire [5:0] T_716;
  wire [7:0] T_720;
  wire [5:0] T_721;
  wire [7:0] T_725;
  wire [5:0] T_726;
  wire [7:0] T_730;
  wire [5:0] T_731;
  wire [7:0] T_735;
  wire [5:0] T_736;
  wire [7:0] T_740;
  wire [5:0] T_741;
  wire [7:0] T_745;
  wire [5:0] T_746;
  wire [7:0] T_750;
  wire [5:0] T_751;
  wire [7:0] T_755;
  wire [5:0] T_756;
  wire [7:0] T_760;
  wire [5:0] T_761;
  wire [7:0] T_765;
  wire [5:0] T_766;
  wire [7:0] T_770;
  wire [5:0] T_771;
  wire [7:0] T_775;
  wire [5:0] T_776;
  wire [7:0] T_780;
  wire [5:0] T_781;
  wire [7:0] T_785;
  wire [5:0] T_786;
  wire [7:0] T_790;
  wire [5:0] T_791;
  wire [7:0] T_795;
  wire [5:0] T_796;
  wire [7:0] T_800;
  wire [5:0] T_801;
  wire [7:0] T_805;
  wire [5:0] T_806;
  wire [7:0] T_810;
  wire [5:0] T_811;
  wire [7:0] T_815;
  wire [5:0] T_816;
  wire [7:0] T_820;
  wire [5:0] T_821;
  wire [7:0] T_825;
  wire [5:0] T_826;
  wire [7:0] T_830;
  wire [5:0] T_831;
  wire [7:0] T_835;
  wire [5:0] T_836;
  wire [7:0] T_840;
  wire [5:0] T_841;
  wire [7:0] T_845;
  wire [5:0] T_846;
  wire [7:0] T_850;
  wire [5:0] T_851;
  wire [7:0] T_855;
  wire [5:0] T_856;
  wire [7:0] T_860;
  wire [5:0] T_861;
  wire [7:0] T_865;
  wire [5:0] T_866;
  wire [7:0] T_870;
  wire [5:0] T_871;
  wire [7:0] T_875;
  wire [5:0] T_876;
  wire [7:0] T_880;
  wire [5:0] T_881;
  wire [7:0] T_885;
  wire [5:0] T_886;
  wire [7:0] T_890;
  wire [5:0] T_891;
  wire [7:0] T_895;
  wire [5:0] T_896;
  wire [7:0] T_900;
  wire [5:0] T_901;
  wire [7:0] T_905;
  wire [5:0] T_906;
  wire [7:0] T_910;
  wire [5:0] T_911;
  wire [7:0] T_915;
  wire [5:0] T_916;
  wire [7:0] T_920;
  wire [5:0] T_921;
  wire [7:0] T_925;
  wire [5:0] T_926;
  wire [7:0] T_930;
  wire [5:0] T_931;
  wire [7:0] T_935;
  wire [5:0] T_936;
  wire [7:0] T_940;
  wire [5:0] T_941;
  wire [7:0] T_945;
  wire [5:0] T_946;
  wire [7:0] T_950;
  wire [5:0] T_951;
  wire [7:0] T_955;
  wire [5:0] T_956;
  wire [7:0] T_960;
  wire [5:0] T_961;
  wire [7:0] T_965;
  wire [5:0] T_966;
  wire [7:0] T_970;
  wire [5:0] T_971;
  wire [7:0] T_975;
  wire [5:0] T_976;
  wire [7:0] T_980;
  wire [5:0] T_981;
  wire [7:0] T_985;
  wire [5:0] T_986;
  wire [7:0] T_990;
  wire [5:0] T_991;
  wire [7:0] T_995;
  wire [5:0] T_996;
  wire [7:0] T_1000;
  wire [5:0] T_1001;
  wire [7:0] T_1005;
  wire [5:0] T_1006;
  wire [7:0] T_1010;
  wire [5:0] T_1011;
  wire [7:0] T_1015;
  wire [5:0] T_1016;
  wire [7:0] T_1020;
  wire [5:0] T_1021;
  wire [7:0] T_1025;
  wire [5:0] T_1026;
  wire [7:0] T_1030;
  wire [5:0] T_1031;
  wire [7:0] T_1035;
  wire [5:0] T_1036;
  wire [7:0] T_1040;
  wire [5:0] T_1041;
  wire [7:0] T_1045;
  wire [5:0] T_1046;
  wire [7:0] T_1050;
  wire [5:0] T_1051;
  wire [7:0] T_1055;
  wire [5:0] T_1056;
  wire [7:0] T_1060;
  wire [5:0] T_1061;
  wire [7:0] T_1065;
  wire [5:0] T_1066;
  wire [7:0] T_1070;
  wire [5:0] T_1071;
  wire [7:0] T_1075;
  wire [5:0] T_1076;
  wire [7:0] T_1080;
  wire [5:0] T_1081;
  wire [7:0] T_1085;
  wire [5:0] T_1086;
  wire [7:0] T_1090;
  wire [5:0] T_1091;
  wire [7:0] T_1095;
  wire [5:0] T_1096;
  wire [7:0] T_1100;
  wire [5:0] T_1101;
  wire [7:0] T_1105;
  wire [5:0] T_1106;
  wire [7:0] T_1110;
  wire [5:0] T_1111;
  wire [7:0] T_1115;
  wire [5:0] T_1116;
  wire [7:0] T_1120;
  wire [5:0] T_1121;
  wire [7:0] T_1125;
  wire [5:0] T_1126;
  wire [7:0] T_1130;
  wire [5:0] T_1131;
  wire [7:0] T_1135;
  wire [5:0] T_1136;
  wire [7:0] T_1140;
  wire [5:0] T_1141;
  wire [7:0] T_1145;
  wire [5:0] T_1146;
  wire [7:0] T_1150;
  wire [5:0] T_1151;
  wire [7:0] T_1155;
  wire [5:0] T_1156;
  wire [7:0] T_1160;
  wire [5:0] T_1161;
  wire [7:0] T_1165;
  wire [5:0] T_1166;
  wire [7:0] T_1170;
  wire [5:0] T_1171;
  wire [7:0] T_1175;
  wire [5:0] T_1176;
  wire [7:0] T_1180;
  wire [5:0] T_1181;
  wire [7:0] T_1185;
  wire [5:0] T_1186;
  wire [7:0] T_1190;
  wire [5:0] T_1191;
  wire [7:0] T_1195;
  wire [5:0] T_1196;
  reg  useRAS_0;
  reg [31:0] GEN_153;
  reg  useRAS_1;
  reg [31:0] GEN_154;
  reg  useRAS_2;
  reg [31:0] GEN_155;
  reg  useRAS_3;
  reg [31:0] GEN_156;
  reg  useRAS_4;
  reg [31:0] GEN_157;
  reg  useRAS_5;
  reg [31:0] GEN_158;
  reg  useRAS_6;
  reg [31:0] GEN_159;
  reg  useRAS_7;
  reg [31:0] GEN_160;
  reg  useRAS_8;
  reg [31:0] GEN_161;
  reg  useRAS_9;
  reg [31:0] GEN_162;
  reg  useRAS_10;
  reg [31:0] GEN_163;
  reg  useRAS_11;
  reg [31:0] GEN_164;
  reg  useRAS_12;
  reg [31:0] GEN_165;
  reg  useRAS_13;
  reg [31:0] GEN_166;
  reg  useRAS_14;
  reg [31:0] GEN_167;
  reg  useRAS_15;
  reg [31:0] GEN_168;
  reg  useRAS_16;
  reg [31:0] GEN_169;
  reg  useRAS_17;
  reg [31:0] GEN_170;
  reg  useRAS_18;
  reg [31:0] GEN_171;
  reg  useRAS_19;
  reg [31:0] GEN_172;
  reg  useRAS_20;
  reg [31:0] GEN_173;
  reg  useRAS_21;
  reg [31:0] GEN_174;
  reg  useRAS_22;
  reg [31:0] GEN_175;
  reg  useRAS_23;
  reg [31:0] GEN_177;
  reg  useRAS_24;
  reg [31:0] GEN_178;
  reg  useRAS_25;
  reg [31:0] GEN_179;
  reg  useRAS_26;
  reg [31:0] GEN_180;
  reg  useRAS_27;
  reg [31:0] GEN_181;
  reg  useRAS_28;
  reg [31:0] GEN_182;
  reg  useRAS_29;
  reg [31:0] GEN_183;
  reg  useRAS_30;
  reg [31:0] GEN_184;
  reg  useRAS_31;
  reg [31:0] GEN_185;
  reg  useRAS_32;
  reg [31:0] GEN_186;
  reg  useRAS_33;
  reg [31:0] GEN_187;
  reg  useRAS_34;
  reg [31:0] GEN_188;
  reg  useRAS_35;
  reg [31:0] GEN_189;
  reg  useRAS_36;
  reg [31:0] GEN_190;
  reg  useRAS_37;
  reg [31:0] GEN_191;
  reg  useRAS_38;
  reg [31:0] GEN_192;
  reg  useRAS_39;
  reg [31:0] GEN_193;
  reg  useRAS_40;
  reg [31:0] GEN_194;
  reg  useRAS_41;
  reg [31:0] GEN_195;
  reg  useRAS_42;
  reg [31:0] GEN_196;
  reg  useRAS_43;
  reg [31:0] GEN_197;
  reg  useRAS_44;
  reg [31:0] GEN_198;
  reg  useRAS_45;
  reg [31:0] GEN_199;
  reg  useRAS_46;
  reg [31:0] GEN_200;
  reg  useRAS_47;
  reg [31:0] GEN_201;
  reg  useRAS_48;
  reg [31:0] GEN_202;
  reg  useRAS_49;
  reg [31:0] GEN_203;
  reg  useRAS_50;
  reg [31:0] GEN_204;
  reg  useRAS_51;
  reg [31:0] GEN_205;
  reg  useRAS_52;
  reg [31:0] GEN_206;
  reg  useRAS_53;
  reg [31:0] GEN_207;
  reg  useRAS_54;
  reg [31:0] GEN_208;
  reg  useRAS_55;
  reg [31:0] GEN_209;
  reg  useRAS_56;
  reg [31:0] GEN_210;
  reg  useRAS_57;
  reg [31:0] GEN_211;
  reg  useRAS_58;
  reg [31:0] GEN_212;
  reg  useRAS_59;
  reg [31:0] GEN_213;
  reg  useRAS_60;
  reg [31:0] GEN_214;
  reg  useRAS_61;
  reg [31:0] GEN_215;
  reg  isJump_0;
  reg [31:0] GEN_216;
  reg  isJump_1;
  reg [31:0] GEN_217;
  reg  isJump_2;
  reg [31:0] GEN_218;
  reg  isJump_3;
  reg [31:0] GEN_219;
  reg  isJump_4;
  reg [31:0] GEN_220;
  reg  isJump_5;
  reg [31:0] GEN_221;
  reg  isJump_6;
  reg [31:0] GEN_222;
  reg  isJump_7;
  reg [31:0] GEN_223;
  reg  isJump_8;
  reg [31:0] GEN_224;
  reg  isJump_9;
  reg [31:0] GEN_225;
  reg  isJump_10;
  reg [31:0] GEN_226;
  reg  isJump_11;
  reg [31:0] GEN_227;
  reg  isJump_12;
  reg [31:0] GEN_228;
  reg  isJump_13;
  reg [31:0] GEN_229;
  reg  isJump_14;
  reg [31:0] GEN_230;
  reg  isJump_15;
  reg [31:0] GEN_231;
  reg  isJump_16;
  reg [31:0] GEN_232;
  reg  isJump_17;
  reg [31:0] GEN_233;
  reg  isJump_18;
  reg [31:0] GEN_234;
  reg  isJump_19;
  reg [31:0] GEN_235;
  reg  isJump_20;
  reg [31:0] GEN_236;
  reg  isJump_21;
  reg [31:0] GEN_237;
  reg  isJump_22;
  reg [31:0] GEN_238;
  reg  isJump_23;
  reg [31:0] GEN_240;
  reg  isJump_24;
  reg [31:0] GEN_241;
  reg  isJump_25;
  reg [31:0] GEN_242;
  reg  isJump_26;
  reg [31:0] GEN_243;
  reg  isJump_27;
  reg [31:0] GEN_244;
  reg  isJump_28;
  reg [31:0] GEN_245;
  reg  isJump_29;
  reg [31:0] GEN_246;
  reg  isJump_30;
  reg [31:0] GEN_247;
  reg  isJump_31;
  reg [31:0] GEN_248;
  reg  isJump_32;
  reg [31:0] GEN_249;
  reg  isJump_33;
  reg [31:0] GEN_250;
  reg  isJump_34;
  reg [31:0] GEN_251;
  reg  isJump_35;
  reg [31:0] GEN_252;
  reg  isJump_36;
  reg [31:0] GEN_253;
  reg  isJump_37;
  reg [31:0] GEN_254;
  reg  isJump_38;
  reg [31:0] GEN_255;
  reg  isJump_39;
  reg [31:0] GEN_256;
  reg  isJump_40;
  reg [31:0] GEN_257;
  reg  isJump_41;
  reg [31:0] GEN_258;
  reg  isJump_42;
  reg [31:0] GEN_259;
  reg  isJump_43;
  reg [31:0] GEN_260;
  reg  isJump_44;
  reg [31:0] GEN_323;
  reg  isJump_45;
  reg [31:0] GEN_386;
  reg  isJump_46;
  reg [31:0] GEN_387;
  reg  isJump_47;
  reg [31:0] GEN_388;
  reg  isJump_48;
  reg [31:0] GEN_389;
  reg  isJump_49;
  reg [31:0] GEN_390;
  reg  isJump_50;
  reg [31:0] GEN_391;
  reg  isJump_51;
  reg [31:0] GEN_392;
  reg  isJump_52;
  reg [31:0] GEN_394;
  reg  isJump_53;
  reg [31:0] GEN_395;
  reg  isJump_54;
  reg [31:0] GEN_396;
  reg  isJump_55;
  reg [31:0] GEN_397;
  reg  isJump_56;
  reg [31:0] GEN_399;
  reg  isJump_57;
  reg [31:0] GEN_400;
  reg  isJump_58;
  reg [31:0] GEN_401;
  reg  isJump_59;
  reg [31:0] GEN_402;
  reg  isJump_60;
  reg [31:0] GEN_404;
  reg  isJump_61;
  reg [31:0] GEN_405;
  reg  brIdx [0:61];
  reg [31:0] GEN_406;
  wire  brIdx_T_3612_data;
  wire [5:0] brIdx_T_3612_addr;
  wire  brIdx_T_3612_en;
  wire  brIdx_T_2876_data;
  wire [5:0] brIdx_T_2876_addr;
  wire  brIdx_T_2876_mask;
  wire  brIdx_T_2876_en;
  reg  T_1215;
  reg [31:0] GEN_407;
  reg  T_1216_prediction_valid;
  reg [31:0] GEN_409;
  reg  T_1216_prediction_bits_taken;
  reg [31:0] GEN_410;
  reg  T_1216_prediction_bits_mask;
  reg [31:0] GEN_411;
  reg  T_1216_prediction_bits_bridx;
  reg [31:0] GEN_412;
  reg [38:0] T_1216_prediction_bits_target;
  reg [63:0] GEN_414;
  reg [5:0] T_1216_prediction_bits_entry;
  reg [31:0] GEN_415;
  reg [6:0] T_1216_prediction_bits_bht_history;
  reg [31:0] GEN_416;
  reg [1:0] T_1216_prediction_bits_bht_value;
  reg [31:0] GEN_417;
  reg [38:0] T_1216_pc;
  reg [63:0] GEN_419;
  reg [38:0] T_1216_target;
  reg [63:0] GEN_420;
  reg  T_1216_taken;
  reg [31:0] GEN_426;
  reg  T_1216_isJump;
  reg [31:0] GEN_427;
  reg  T_1216_isReturn;
  reg [31:0] GEN_428;
  reg [38:0] T_1216_br_pc;
  reg [63:0] GEN_429;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [38:0] GEN_8;
  wire [5:0] GEN_9;
  wire [6:0] GEN_10;
  wire [1:0] GEN_11;
  wire [38:0] GEN_12;
  wire [38:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [38:0] GEN_17;
  wire  r_btb_update_valid;
  wire  r_btb_update_bits_prediction_valid;
  wire  r_btb_update_bits_prediction_bits_taken;
  wire  r_btb_update_bits_prediction_bits_mask;
  wire  r_btb_update_bits_prediction_bits_bridx;
  wire [38:0] r_btb_update_bits_prediction_bits_target;
  wire [5:0] r_btb_update_bits_prediction_bits_entry;
  wire [6:0] r_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] r_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] r_btb_update_bits_pc;
  wire [38:0] r_btb_update_bits_target;
  wire  r_btb_update_bits_taken;
  wire  r_btb_update_bits_isJump;
  wire  r_btb_update_bits_isReturn;
  wire [38:0] r_btb_update_bits_br_pc;
  wire [26:0] T_1398;
  wire  T_1401;
  wire  T_1404;
  wire  T_1407;
  wire  T_1410;
  wire  T_1413;
  wire  T_1416;
  wire  T_1422_0;
  wire  T_1422_1;
  wire  T_1422_2;
  wire  T_1422_3;
  wire  T_1422_4;
  wire  T_1422_5;
  wire [1:0] T_1424;
  wire [2:0] T_1425;
  wire [1:0] T_1426;
  wire [2:0] T_1427;
  wire [5:0] T_1428;
  wire [5:0] pageHit;
  wire [11:0] T_1429;
  wire  T_1432;
  wire  T_1435;
  wire  T_1438;
  wire  T_1441;
  wire  T_1444;
  wire  T_1447;
  wire  T_1450;
  wire  T_1453;
  wire  T_1456;
  wire  T_1459;
  wire  T_1462;
  wire  T_1465;
  wire  T_1468;
  wire  T_1471;
  wire  T_1474;
  wire  T_1477;
  wire  T_1480;
  wire  T_1483;
  wire  T_1486;
  wire  T_1489;
  wire  T_1492;
  wire  T_1495;
  wire  T_1498;
  wire  T_1501;
  wire  T_1504;
  wire  T_1507;
  wire  T_1510;
  wire  T_1513;
  wire  T_1516;
  wire  T_1519;
  wire  T_1522;
  wire  T_1525;
  wire  T_1528;
  wire  T_1531;
  wire  T_1534;
  wire  T_1537;
  wire  T_1540;
  wire  T_1543;
  wire  T_1546;
  wire  T_1549;
  wire  T_1552;
  wire  T_1555;
  wire  T_1558;
  wire  T_1561;
  wire  T_1564;
  wire  T_1567;
  wire  T_1570;
  wire  T_1573;
  wire  T_1576;
  wire  T_1579;
  wire  T_1582;
  wire  T_1585;
  wire  T_1588;
  wire  T_1591;
  wire  T_1594;
  wire  T_1597;
  wire  T_1600;
  wire  T_1603;
  wire  T_1606;
  wire  T_1609;
  wire  T_1612;
  wire  T_1615;
  wire  T_1621_0;
  wire  T_1621_1;
  wire  T_1621_2;
  wire  T_1621_3;
  wire  T_1621_4;
  wire  T_1621_5;
  wire  T_1621_6;
  wire  T_1621_7;
  wire  T_1621_8;
  wire  T_1621_9;
  wire  T_1621_10;
  wire  T_1621_11;
  wire  T_1621_12;
  wire  T_1621_13;
  wire  T_1621_14;
  wire  T_1621_15;
  wire  T_1621_16;
  wire  T_1621_17;
  wire  T_1621_18;
  wire  T_1621_19;
  wire  T_1621_20;
  wire  T_1621_21;
  wire  T_1621_22;
  wire  T_1621_23;
  wire  T_1621_24;
  wire  T_1621_25;
  wire  T_1621_26;
  wire  T_1621_27;
  wire  T_1621_28;
  wire  T_1621_29;
  wire  T_1621_30;
  wire  T_1621_31;
  wire  T_1621_32;
  wire  T_1621_33;
  wire  T_1621_34;
  wire  T_1621_35;
  wire  T_1621_36;
  wire  T_1621_37;
  wire  T_1621_38;
  wire  T_1621_39;
  wire  T_1621_40;
  wire  T_1621_41;
  wire  T_1621_42;
  wire  T_1621_43;
  wire  T_1621_44;
  wire  T_1621_45;
  wire  T_1621_46;
  wire  T_1621_47;
  wire  T_1621_48;
  wire  T_1621_49;
  wire  T_1621_50;
  wire  T_1621_51;
  wire  T_1621_52;
  wire  T_1621_53;
  wire  T_1621_54;
  wire  T_1621_55;
  wire  T_1621_56;
  wire  T_1621_57;
  wire  T_1621_58;
  wire  T_1621_59;
  wire  T_1621_60;
  wire  T_1621_61;
  wire [1:0] T_1623;
  wire [2:0] T_1624;
  wire [1:0] T_1625;
  wire [1:0] T_1626;
  wire [3:0] T_1627;
  wire [6:0] T_1628;
  wire [1:0] T_1629;
  wire [1:0] T_1630;
  wire [3:0] T_1631;
  wire [1:0] T_1632;
  wire [1:0] T_1633;
  wire [3:0] T_1634;
  wire [7:0] T_1635;
  wire [14:0] T_1636;
  wire [1:0] T_1637;
  wire [1:0] T_1638;
  wire [3:0] T_1639;
  wire [1:0] T_1640;
  wire [1:0] T_1641;
  wire [3:0] T_1642;
  wire [7:0] T_1643;
  wire [1:0] T_1644;
  wire [1:0] T_1645;
  wire [3:0] T_1646;
  wire [1:0] T_1647;
  wire [1:0] T_1648;
  wire [3:0] T_1649;
  wire [7:0] T_1650;
  wire [15:0] T_1651;
  wire [30:0] T_1652;
  wire [1:0] T_1653;
  wire [2:0] T_1654;
  wire [1:0] T_1655;
  wire [1:0] T_1656;
  wire [3:0] T_1657;
  wire [6:0] T_1658;
  wire [1:0] T_1659;
  wire [1:0] T_1660;
  wire [3:0] T_1661;
  wire [1:0] T_1662;
  wire [1:0] T_1663;
  wire [3:0] T_1664;
  wire [7:0] T_1665;
  wire [14:0] T_1666;
  wire [1:0] T_1667;
  wire [1:0] T_1668;
  wire [3:0] T_1669;
  wire [1:0] T_1670;
  wire [1:0] T_1671;
  wire [3:0] T_1672;
  wire [7:0] T_1673;
  wire [1:0] T_1674;
  wire [1:0] T_1675;
  wire [3:0] T_1676;
  wire [1:0] T_1677;
  wire [1:0] T_1678;
  wire [3:0] T_1679;
  wire [7:0] T_1680;
  wire [15:0] T_1681;
  wire [30:0] T_1682;
  wire [61:0] T_1683;
  wire [5:0] T_1684;
  wire [5:0] T_1685;
  wire [5:0] T_1686;
  wire [5:0] T_1687;
  wire [5:0] T_1688;
  wire [5:0] T_1689;
  wire [5:0] T_1690;
  wire [5:0] T_1691;
  wire [5:0] T_1692;
  wire [5:0] T_1693;
  wire [5:0] T_1694;
  wire [5:0] T_1695;
  wire [5:0] T_1696;
  wire [5:0] T_1697;
  wire [5:0] T_1698;
  wire [5:0] T_1699;
  wire [5:0] T_1700;
  wire [5:0] T_1701;
  wire [5:0] T_1702;
  wire [5:0] T_1703;
  wire [5:0] T_1704;
  wire [5:0] T_1705;
  wire [5:0] T_1706;
  wire [5:0] T_1707;
  wire [5:0] T_1708;
  wire [5:0] T_1709;
  wire [5:0] T_1710;
  wire [5:0] T_1711;
  wire [5:0] T_1712;
  wire [5:0] T_1713;
  wire [5:0] T_1714;
  wire [5:0] T_1715;
  wire [5:0] T_1716;
  wire [5:0] T_1717;
  wire [5:0] T_1718;
  wire [5:0] T_1719;
  wire [5:0] T_1720;
  wire [5:0] T_1721;
  wire [5:0] T_1722;
  wire [5:0] T_1723;
  wire [5:0] T_1724;
  wire [5:0] T_1725;
  wire [5:0] T_1726;
  wire [5:0] T_1727;
  wire [5:0] T_1728;
  wire [5:0] T_1729;
  wire [5:0] T_1730;
  wire [5:0] T_1731;
  wire [5:0] T_1732;
  wire [5:0] T_1733;
  wire [5:0] T_1734;
  wire [5:0] T_1735;
  wire [5:0] T_1736;
  wire [5:0] T_1737;
  wire [5:0] T_1738;
  wire [5:0] T_1739;
  wire [5:0] T_1740;
  wire [5:0] T_1741;
  wire [5:0] T_1742;
  wire [5:0] T_1743;
  wire [5:0] T_1744;
  wire [5:0] T_1745;
  wire [5:0] GEN_581;
  wire  T_1747;
  wire  T_1749;
  wire  T_1751;
  wire  T_1753;
  wire  T_1755;
  wire  T_1757;
  wire  T_1759;
  wire  T_1761;
  wire  T_1763;
  wire  T_1765;
  wire  T_1767;
  wire  T_1769;
  wire  T_1771;
  wire  T_1773;
  wire  T_1775;
  wire  T_1777;
  wire  T_1779;
  wire  T_1781;
  wire  T_1783;
  wire  T_1785;
  wire  T_1787;
  wire  T_1789;
  wire  T_1791;
  wire  T_1793;
  wire  T_1795;
  wire  T_1797;
  wire  T_1799;
  wire  T_1801;
  wire  T_1803;
  wire  T_1805;
  wire  T_1807;
  wire  T_1809;
  wire  T_1811;
  wire  T_1813;
  wire  T_1815;
  wire  T_1817;
  wire  T_1819;
  wire  T_1821;
  wire  T_1823;
  wire  T_1825;
  wire  T_1827;
  wire  T_1829;
  wire  T_1831;
  wire  T_1833;
  wire  T_1835;
  wire  T_1837;
  wire  T_1839;
  wire  T_1841;
  wire  T_1843;
  wire  T_1845;
  wire  T_1847;
  wire  T_1849;
  wire  T_1851;
  wire  T_1853;
  wire  T_1855;
  wire  T_1857;
  wire  T_1859;
  wire  T_1861;
  wire  T_1863;
  wire  T_1865;
  wire  T_1867;
  wire  T_1869;
  wire  T_1875_0;
  wire  T_1875_1;
  wire  T_1875_2;
  wire  T_1875_3;
  wire  T_1875_4;
  wire  T_1875_5;
  wire  T_1875_6;
  wire  T_1875_7;
  wire  T_1875_8;
  wire  T_1875_9;
  wire  T_1875_10;
  wire  T_1875_11;
  wire  T_1875_12;
  wire  T_1875_13;
  wire  T_1875_14;
  wire  T_1875_15;
  wire  T_1875_16;
  wire  T_1875_17;
  wire  T_1875_18;
  wire  T_1875_19;
  wire  T_1875_20;
  wire  T_1875_21;
  wire  T_1875_22;
  wire  T_1875_23;
  wire  T_1875_24;
  wire  T_1875_25;
  wire  T_1875_26;
  wire  T_1875_27;
  wire  T_1875_28;
  wire  T_1875_29;
  wire  T_1875_30;
  wire  T_1875_31;
  wire  T_1875_32;
  wire  T_1875_33;
  wire  T_1875_34;
  wire  T_1875_35;
  wire  T_1875_36;
  wire  T_1875_37;
  wire  T_1875_38;
  wire  T_1875_39;
  wire  T_1875_40;
  wire  T_1875_41;
  wire  T_1875_42;
  wire  T_1875_43;
  wire  T_1875_44;
  wire  T_1875_45;
  wire  T_1875_46;
  wire  T_1875_47;
  wire  T_1875_48;
  wire  T_1875_49;
  wire  T_1875_50;
  wire  T_1875_51;
  wire  T_1875_52;
  wire  T_1875_53;
  wire  T_1875_54;
  wire  T_1875_55;
  wire  T_1875_56;
  wire  T_1875_57;
  wire  T_1875_58;
  wire  T_1875_59;
  wire  T_1875_60;
  wire  T_1875_61;
  wire [1:0] T_1877;
  wire [2:0] T_1878;
  wire [1:0] T_1879;
  wire [1:0] T_1880;
  wire [3:0] T_1881;
  wire [6:0] T_1882;
  wire [1:0] T_1883;
  wire [1:0] T_1884;
  wire [3:0] T_1885;
  wire [1:0] T_1886;
  wire [1:0] T_1887;
  wire [3:0] T_1888;
  wire [7:0] T_1889;
  wire [14:0] T_1890;
  wire [1:0] T_1891;
  wire [1:0] T_1892;
  wire [3:0] T_1893;
  wire [1:0] T_1894;
  wire [1:0] T_1895;
  wire [3:0] T_1896;
  wire [7:0] T_1897;
  wire [1:0] T_1898;
  wire [1:0] T_1899;
  wire [3:0] T_1900;
  wire [1:0] T_1901;
  wire [1:0] T_1902;
  wire [3:0] T_1903;
  wire [7:0] T_1904;
  wire [15:0] T_1905;
  wire [30:0] T_1906;
  wire [1:0] T_1907;
  wire [2:0] T_1908;
  wire [1:0] T_1909;
  wire [1:0] T_1910;
  wire [3:0] T_1911;
  wire [6:0] T_1912;
  wire [1:0] T_1913;
  wire [1:0] T_1914;
  wire [3:0] T_1915;
  wire [1:0] T_1916;
  wire [1:0] T_1917;
  wire [3:0] T_1918;
  wire [7:0] T_1919;
  wire [14:0] T_1920;
  wire [1:0] T_1921;
  wire [1:0] T_1922;
  wire [3:0] T_1923;
  wire [1:0] T_1924;
  wire [1:0] T_1925;
  wire [3:0] T_1926;
  wire [7:0] T_1927;
  wire [1:0] T_1928;
  wire [1:0] T_1929;
  wire [3:0] T_1930;
  wire [1:0] T_1931;
  wire [1:0] T_1932;
  wire [3:0] T_1933;
  wire [7:0] T_1934;
  wire [15:0] T_1935;
  wire [30:0] T_1936;
  wire [61:0] T_1937;
  wire [61:0] T_1938;
  wire [61:0] hits;
  wire [26:0] T_1939;
  wire  T_1942;
  wire  T_1945;
  wire  T_1948;
  wire  T_1951;
  wire  T_1954;
  wire  T_1957;
  wire  T_1963_0;
  wire  T_1963_1;
  wire  T_1963_2;
  wire  T_1963_3;
  wire  T_1963_4;
  wire  T_1963_5;
  wire [1:0] T_1965;
  wire [2:0] T_1966;
  wire [1:0] T_1967;
  wire [2:0] T_1968;
  wire [5:0] T_1969;
  wire [5:0] updatePageHit;
  wire [11:0] T_1970;
  wire  T_1973;
  wire  T_1976;
  wire  T_1979;
  wire  T_1982;
  wire  T_1985;
  wire  T_1988;
  wire  T_1991;
  wire  T_1994;
  wire  T_1997;
  wire  T_2000;
  wire  T_2003;
  wire  T_2006;
  wire  T_2009;
  wire  T_2012;
  wire  T_2015;
  wire  T_2018;
  wire  T_2021;
  wire  T_2024;
  wire  T_2027;
  wire  T_2030;
  wire  T_2033;
  wire  T_2036;
  wire  T_2039;
  wire  T_2042;
  wire  T_2045;
  wire  T_2048;
  wire  T_2051;
  wire  T_2054;
  wire  T_2057;
  wire  T_2060;
  wire  T_2063;
  wire  T_2066;
  wire  T_2069;
  wire  T_2072;
  wire  T_2075;
  wire  T_2078;
  wire  T_2081;
  wire  T_2084;
  wire  T_2087;
  wire  T_2090;
  wire  T_2093;
  wire  T_2096;
  wire  T_2099;
  wire  T_2102;
  wire  T_2105;
  wire  T_2108;
  wire  T_2111;
  wire  T_2114;
  wire  T_2117;
  wire  T_2120;
  wire  T_2123;
  wire  T_2126;
  wire  T_2129;
  wire  T_2132;
  wire  T_2135;
  wire  T_2138;
  wire  T_2141;
  wire  T_2144;
  wire  T_2147;
  wire  T_2150;
  wire  T_2153;
  wire  T_2156;
  wire  T_2162_0;
  wire  T_2162_1;
  wire  T_2162_2;
  wire  T_2162_3;
  wire  T_2162_4;
  wire  T_2162_5;
  wire  T_2162_6;
  wire  T_2162_7;
  wire  T_2162_8;
  wire  T_2162_9;
  wire  T_2162_10;
  wire  T_2162_11;
  wire  T_2162_12;
  wire  T_2162_13;
  wire  T_2162_14;
  wire  T_2162_15;
  wire  T_2162_16;
  wire  T_2162_17;
  wire  T_2162_18;
  wire  T_2162_19;
  wire  T_2162_20;
  wire  T_2162_21;
  wire  T_2162_22;
  wire  T_2162_23;
  wire  T_2162_24;
  wire  T_2162_25;
  wire  T_2162_26;
  wire  T_2162_27;
  wire  T_2162_28;
  wire  T_2162_29;
  wire  T_2162_30;
  wire  T_2162_31;
  wire  T_2162_32;
  wire  T_2162_33;
  wire  T_2162_34;
  wire  T_2162_35;
  wire  T_2162_36;
  wire  T_2162_37;
  wire  T_2162_38;
  wire  T_2162_39;
  wire  T_2162_40;
  wire  T_2162_41;
  wire  T_2162_42;
  wire  T_2162_43;
  wire  T_2162_44;
  wire  T_2162_45;
  wire  T_2162_46;
  wire  T_2162_47;
  wire  T_2162_48;
  wire  T_2162_49;
  wire  T_2162_50;
  wire  T_2162_51;
  wire  T_2162_52;
  wire  T_2162_53;
  wire  T_2162_54;
  wire  T_2162_55;
  wire  T_2162_56;
  wire  T_2162_57;
  wire  T_2162_58;
  wire  T_2162_59;
  wire  T_2162_60;
  wire  T_2162_61;
  wire [5:0] T_2225;
  wire [5:0] T_2226;
  wire [5:0] T_2227;
  wire [5:0] T_2228;
  wire [5:0] T_2229;
  wire [5:0] T_2230;
  wire [5:0] T_2231;
  wire [5:0] T_2232;
  wire [5:0] T_2233;
  wire [5:0] T_2234;
  wire [5:0] T_2235;
  wire [5:0] T_2236;
  wire [5:0] T_2237;
  wire [5:0] T_2238;
  wire [5:0] T_2239;
  wire [5:0] T_2240;
  wire [5:0] T_2241;
  wire [5:0] T_2242;
  wire [5:0] T_2243;
  wire [5:0] T_2244;
  wire [5:0] T_2245;
  wire [5:0] T_2246;
  wire [5:0] T_2247;
  wire [5:0] T_2248;
  wire [5:0] T_2249;
  wire [5:0] T_2250;
  wire [5:0] T_2251;
  wire [5:0] T_2252;
  wire [5:0] T_2253;
  wire [5:0] T_2254;
  wire [5:0] T_2255;
  wire [5:0] T_2256;
  wire [5:0] T_2257;
  wire [5:0] T_2258;
  wire [5:0] T_2259;
  wire [5:0] T_2260;
  wire [5:0] T_2261;
  wire [5:0] T_2262;
  wire [5:0] T_2263;
  wire [5:0] T_2264;
  wire [5:0] T_2265;
  wire [5:0] T_2266;
  wire [5:0] T_2267;
  wire [5:0] T_2268;
  wire [5:0] T_2269;
  wire [5:0] T_2270;
  wire [5:0] T_2271;
  wire [5:0] T_2272;
  wire [5:0] T_2273;
  wire [5:0] T_2274;
  wire [5:0] T_2275;
  wire [5:0] T_2276;
  wire [5:0] T_2277;
  wire [5:0] T_2278;
  wire [5:0] T_2279;
  wire [5:0] T_2280;
  wire [5:0] T_2281;
  wire [5:0] T_2282;
  wire [5:0] T_2283;
  wire [5:0] T_2284;
  wire [5:0] T_2285;
  wire [5:0] T_2286;
  wire  T_2288;
  wire  T_2290;
  wire  T_2292;
  wire  T_2294;
  wire  T_2296;
  wire  T_2298;
  wire  T_2300;
  wire  T_2302;
  wire  T_2304;
  wire  T_2306;
  wire  T_2308;
  wire  T_2310;
  wire  T_2312;
  wire  T_2314;
  wire  T_2316;
  wire  T_2318;
  wire  T_2320;
  wire  T_2322;
  wire  T_2324;
  wire  T_2326;
  wire  T_2328;
  wire  T_2330;
  wire  T_2332;
  wire  T_2334;
  wire  T_2336;
  wire  T_2338;
  wire  T_2340;
  wire  T_2342;
  wire  T_2344;
  wire  T_2346;
  wire  T_2348;
  wire  T_2350;
  wire  T_2352;
  wire  T_2354;
  wire  T_2356;
  wire  T_2358;
  wire  T_2360;
  wire  T_2362;
  wire  T_2364;
  wire  T_2366;
  wire  T_2368;
  wire  T_2370;
  wire  T_2372;
  wire  T_2374;
  wire  T_2376;
  wire  T_2378;
  wire  T_2380;
  wire  T_2382;
  wire  T_2384;
  wire  T_2386;
  wire  T_2388;
  wire  T_2390;
  wire  T_2392;
  wire  T_2394;
  wire  T_2396;
  wire  T_2398;
  wire  T_2400;
  wire  T_2402;
  wire  T_2404;
  wire  T_2406;
  wire  T_2408;
  wire  T_2410;
  wire  T_2416_0;
  wire  T_2416_1;
  wire  T_2416_2;
  wire  T_2416_3;
  wire  T_2416_4;
  wire  T_2416_5;
  wire  T_2416_6;
  wire  T_2416_7;
  wire  T_2416_8;
  wire  T_2416_9;
  wire  T_2416_10;
  wire  T_2416_11;
  wire  T_2416_12;
  wire  T_2416_13;
  wire  T_2416_14;
  wire  T_2416_15;
  wire  T_2416_16;
  wire  T_2416_17;
  wire  T_2416_18;
  wire  T_2416_19;
  wire  T_2416_20;
  wire  T_2416_21;
  wire  T_2416_22;
  wire  T_2416_23;
  wire  T_2416_24;
  wire  T_2416_25;
  wire  T_2416_26;
  wire  T_2416_27;
  wire  T_2416_28;
  wire  T_2416_29;
  wire  T_2416_30;
  wire  T_2416_31;
  wire  T_2416_32;
  wire  T_2416_33;
  wire  T_2416_34;
  wire  T_2416_35;
  wire  T_2416_36;
  wire  T_2416_37;
  wire  T_2416_38;
  wire  T_2416_39;
  wire  T_2416_40;
  wire  T_2416_41;
  wire  T_2416_42;
  wire  T_2416_43;
  wire  T_2416_44;
  wire  T_2416_45;
  wire  T_2416_46;
  wire  T_2416_47;
  wire  T_2416_48;
  wire  T_2416_49;
  wire  T_2416_50;
  wire  T_2416_51;
  wire  T_2416_52;
  wire  T_2416_53;
  wire  T_2416_54;
  wire  T_2416_55;
  wire  T_2416_56;
  wire  T_2416_57;
  wire  T_2416_58;
  wire  T_2416_59;
  wire  T_2416_60;
  wire  T_2416_61;
  wire  T_2481;
  wire  T_2482;
  reg [5:0] nextRepl;
  reg [31:0] GEN_430;
  wire  T_2485;
  wire [5:0] GEN_705;
  wire [6:0] T_2487;
  wire [5:0] T_2488;
  wire [5:0] GEN_18;
  wire [5:0] GEN_19;
  wire  useUpdatePageHit;
  wire  doIdxPageRepl;
  wire [5:0] idxPageRepl;
  wire [5:0] idxPageUpdateOH;
  wire [1:0] T_2494;
  wire [3:0] T_2495;
  wire [1:0] GEN_707;
  wire  T_2497;
  wire [3:0] GEN_708;
  wire [3:0] T_2498;
  wire [1:0] T_2499;
  wire [1:0] T_2500;
  wire  T_2502;
  wire [1:0] T_2503;
  wire  T_2504;
  wire [1:0] T_2505;
  wire [2:0] idxPageUpdate;
  wire [5:0] idxPageReplEn;
  wire  samePage;
  wire [5:0] T_2509;
  wire [5:0] T_2510;
  wire  usePageHit;
  wire  T_2513;
  wire  T_2515;
  wire  doTgtPageRepl;
  wire [4:0] T_2516;
  wire [5:0] GEN_711;
  wire [5:0] T_2517;
  wire  T_2518;
  wire [5:0] GEN_712;
  wire [5:0] T_2519;
  wire [5:0] tgtPageRepl;
  wire [5:0] T_2520;
  wire [1:0] T_2521;
  wire [3:0] T_2522;
  wire  T_2524;
  wire [3:0] GEN_714;
  wire [3:0] T_2525;
  wire [1:0] T_2526;
  wire [1:0] T_2527;
  wire  T_2529;
  wire [1:0] T_2530;
  wire  T_2531;
  wire [1:0] T_2532;
  wire [2:0] tgtPageUpdate;
  wire [5:0] tgtPageReplEn;
  wire  doPageRepl;
  wire [5:0] pageReplEn;
  wire  T_2534;
  reg [2:0] T_2536;
  reg [31:0] GEN_434;
  wire  T_2538;
  wire [2:0] GEN_716;
  wire [3:0] T_2540;
  wire [2:0] T_2541;
  wire [2:0] GEN_20;
  wire [2:0] GEN_21;
  wire [7:0] T_2545;
  wire  T_2546;
  wire  T_2547;
  wire  T_2549;
  wire [5:0] T_2550;
  wire [5:0] T_2551;
  wire [5:0] T_2552;
  wire  T_2554;
  wire [5:0] T_2555;
  wire [5:0] T_2556;
  wire  T_2558;
  wire [5:0] T_2559;
  wire [5:0] T_2560;
  wire  T_2562;
  wire [5:0] T_2563;
  wire [5:0] T_2564;
  wire  T_2566;
  wire [5:0] T_2567;
  wire [5:0] T_2568;
  wire  T_2570;
  wire [5:0] T_2571;
  wire [5:0] T_2572;
  wire  T_2574;
  wire [5:0] T_2575;
  wire [5:0] T_2576;
  wire  T_2578;
  wire [5:0] T_2579;
  wire [5:0] T_2580;
  wire  T_2582;
  wire [5:0] T_2583;
  wire [5:0] T_2584;
  wire  T_2586;
  wire [5:0] T_2587;
  wire [5:0] T_2588;
  wire  T_2590;
  wire [5:0] T_2591;
  wire [5:0] T_2592;
  wire  T_2594;
  wire [5:0] T_2595;
  wire [5:0] T_2596;
  wire  T_2598;
  wire [5:0] T_2599;
  wire [5:0] T_2600;
  wire  T_2602;
  wire [5:0] T_2603;
  wire [5:0] T_2604;
  wire  T_2606;
  wire [5:0] T_2607;
  wire [5:0] T_2608;
  wire  T_2610;
  wire [5:0] T_2611;
  wire [5:0] T_2612;
  wire  T_2614;
  wire [5:0] T_2615;
  wire [5:0] T_2616;
  wire  T_2618;
  wire [5:0] T_2619;
  wire [5:0] T_2620;
  wire  T_2622;
  wire [5:0] T_2623;
  wire [5:0] T_2624;
  wire  T_2626;
  wire [5:0] T_2627;
  wire [5:0] T_2628;
  wire  T_2630;
  wire [5:0] T_2631;
  wire [5:0] T_2632;
  wire  T_2634;
  wire [5:0] T_2635;
  wire [5:0] T_2636;
  wire  T_2638;
  wire [5:0] T_2639;
  wire [5:0] T_2640;
  wire  T_2642;
  wire [5:0] T_2643;
  wire [5:0] T_2644;
  wire  T_2646;
  wire [5:0] T_2647;
  wire [5:0] T_2648;
  wire  T_2650;
  wire [5:0] T_2651;
  wire [5:0] T_2652;
  wire  T_2654;
  wire [5:0] T_2655;
  wire [5:0] T_2656;
  wire  T_2658;
  wire [5:0] T_2659;
  wire [5:0] T_2660;
  wire  T_2662;
  wire [5:0] T_2663;
  wire [5:0] T_2664;
  wire  T_2666;
  wire [5:0] T_2667;
  wire [5:0] T_2668;
  wire  T_2670;
  wire [5:0] T_2671;
  wire [5:0] T_2672;
  wire  T_2674;
  wire [5:0] T_2675;
  wire [5:0] T_2676;
  wire  T_2678;
  wire [5:0] T_2679;
  wire [5:0] T_2680;
  wire  T_2682;
  wire [5:0] T_2683;
  wire [5:0] T_2684;
  wire  T_2686;
  wire [5:0] T_2687;
  wire [5:0] T_2688;
  wire  T_2690;
  wire [5:0] T_2691;
  wire [5:0] T_2692;
  wire  T_2694;
  wire [5:0] T_2695;
  wire [5:0] T_2696;
  wire  T_2698;
  wire [5:0] T_2699;
  wire [5:0] T_2700;
  wire  T_2702;
  wire [5:0] T_2703;
  wire [5:0] T_2704;
  wire  T_2706;
  wire [5:0] T_2707;
  wire [5:0] T_2708;
  wire  T_2710;
  wire [5:0] T_2711;
  wire [5:0] T_2712;
  wire  T_2714;
  wire [5:0] T_2715;
  wire [5:0] T_2716;
  wire  T_2718;
  wire [5:0] T_2719;
  wire [5:0] T_2720;
  wire  T_2722;
  wire [5:0] T_2723;
  wire [5:0] T_2724;
  wire  T_2726;
  wire [5:0] T_2727;
  wire [5:0] T_2728;
  wire  T_2730;
  wire [5:0] T_2731;
  wire [5:0] T_2732;
  wire  T_2734;
  wire [5:0] T_2735;
  wire [5:0] T_2736;
  wire  T_2738;
  wire [5:0] T_2739;
  wire [5:0] T_2740;
  wire  T_2742;
  wire [5:0] T_2743;
  wire [5:0] T_2744;
  wire  T_2746;
  wire [5:0] T_2747;
  wire [5:0] T_2748;
  wire  T_2750;
  wire [5:0] T_2751;
  wire [5:0] T_2752;
  wire  T_2754;
  wire [5:0] T_2755;
  wire [5:0] T_2756;
  wire  T_2758;
  wire [5:0] T_2759;
  wire [5:0] T_2760;
  wire  T_2762;
  wire [5:0] T_2763;
  wire [5:0] T_2764;
  wire  T_2766;
  wire [5:0] T_2767;
  wire [5:0] T_2768;
  wire  T_2770;
  wire [5:0] T_2771;
  wire [5:0] T_2772;
  wire  T_2774;
  wire [5:0] T_2775;
  wire [5:0] T_2776;
  wire  T_2778;
  wire [5:0] T_2779;
  wire [5:0] T_2780;
  wire  T_2782;
  wire [5:0] T_2783;
  wire [5:0] T_2784;
  wire  T_2786;
  wire [5:0] T_2787;
  wire [5:0] T_2788;
  wire  T_2790;
  wire [5:0] T_2791;
  wire [5:0] T_2792;
  wire  T_2794;
  wire [5:0] T_2795;
  wire [5:0] T_2796;
  wire  T_2798;
  wire  T_2804_0;
  wire  T_2804_1;
  wire  T_2804_2;
  wire  T_2804_3;
  wire  T_2804_4;
  wire  T_2804_5;
  wire  T_2804_6;
  wire  T_2804_7;
  wire  T_2804_8;
  wire  T_2804_9;
  wire  T_2804_10;
  wire  T_2804_11;
  wire  T_2804_12;
  wire  T_2804_13;
  wire  T_2804_14;
  wire  T_2804_15;
  wire  T_2804_16;
  wire  T_2804_17;
  wire  T_2804_18;
  wire  T_2804_19;
  wire  T_2804_20;
  wire  T_2804_21;
  wire  T_2804_22;
  wire  T_2804_23;
  wire  T_2804_24;
  wire  T_2804_25;
  wire  T_2804_26;
  wire  T_2804_27;
  wire  T_2804_28;
  wire  T_2804_29;
  wire  T_2804_30;
  wire  T_2804_31;
  wire  T_2804_32;
  wire  T_2804_33;
  wire  T_2804_34;
  wire  T_2804_35;
  wire  T_2804_36;
  wire  T_2804_37;
  wire  T_2804_38;
  wire  T_2804_39;
  wire  T_2804_40;
  wire  T_2804_41;
  wire  T_2804_42;
  wire  T_2804_43;
  wire  T_2804_44;
  wire  T_2804_45;
  wire  T_2804_46;
  wire  T_2804_47;
  wire  T_2804_48;
  wire  T_2804_49;
  wire  T_2804_50;
  wire  T_2804_51;
  wire  T_2804_52;
  wire  T_2804_53;
  wire  T_2804_54;
  wire  T_2804_55;
  wire  T_2804_56;
  wire  T_2804_57;
  wire  T_2804_58;
  wire  T_2804_59;
  wire  T_2804_60;
  wire  T_2804_61;
  wire [1:0] T_2806;
  wire [2:0] T_2807;
  wire [1:0] T_2808;
  wire [1:0] T_2809;
  wire [3:0] T_2810;
  wire [6:0] T_2811;
  wire [1:0] T_2812;
  wire [1:0] T_2813;
  wire [3:0] T_2814;
  wire [1:0] T_2815;
  wire [1:0] T_2816;
  wire [3:0] T_2817;
  wire [7:0] T_2818;
  wire [14:0] T_2819;
  wire [1:0] T_2820;
  wire [1:0] T_2821;
  wire [3:0] T_2822;
  wire [1:0] T_2823;
  wire [1:0] T_2824;
  wire [3:0] T_2825;
  wire [7:0] T_2826;
  wire [1:0] T_2827;
  wire [1:0] T_2828;
  wire [3:0] T_2829;
  wire [1:0] T_2830;
  wire [1:0] T_2831;
  wire [3:0] T_2832;
  wire [7:0] T_2833;
  wire [15:0] T_2834;
  wire [30:0] T_2835;
  wire [1:0] T_2836;
  wire [2:0] T_2837;
  wire [1:0] T_2838;
  wire [1:0] T_2839;
  wire [3:0] T_2840;
  wire [6:0] T_2841;
  wire [1:0] T_2842;
  wire [1:0] T_2843;
  wire [3:0] T_2844;
  wire [1:0] T_2845;
  wire [1:0] T_2846;
  wire [3:0] T_2847;
  wire [7:0] T_2848;
  wire [14:0] T_2849;
  wire [1:0] T_2850;
  wire [1:0] T_2851;
  wire [3:0] T_2852;
  wire [1:0] T_2853;
  wire [1:0] T_2854;
  wire [3:0] T_2855;
  wire [7:0] T_2856;
  wire [1:0] T_2857;
  wire [1:0] T_2858;
  wire [3:0] T_2859;
  wire [1:0] T_2860;
  wire [1:0] T_2861;
  wire [3:0] T_2862;
  wire [7:0] T_2863;
  wire [15:0] T_2864;
  wire [30:0] T_2865;
  wire [61:0] T_2866;
  wire [63:0] GEN_780;
  wire [63:0] T_2868;
  wire [61:0] T_2869;
  wire [61:0] T_2870;
  wire [63:0] GEN_781;
  wire [63:0] T_2871;
  wire  GEN_0;
  wire  GEN_22;
  wire  GEN_23;
  wire [5:0] GEN_784;
  wire  GEN_24;
  wire [5:0] GEN_785;
  wire  GEN_25;
  wire [5:0] GEN_786;
  wire  GEN_26;
  wire [5:0] GEN_787;
  wire  GEN_27;
  wire [5:0] GEN_788;
  wire  GEN_28;
  wire [5:0] GEN_789;
  wire  GEN_29;
  wire [5:0] GEN_790;
  wire  GEN_30;
  wire [5:0] GEN_791;
  wire  GEN_31;
  wire [5:0] GEN_792;
  wire  GEN_32;
  wire [5:0] GEN_793;
  wire  GEN_33;
  wire [5:0] GEN_794;
  wire  GEN_34;
  wire [5:0] GEN_795;
  wire  GEN_35;
  wire [5:0] GEN_796;
  wire  GEN_36;
  wire [5:0] GEN_797;
  wire  GEN_37;
  wire [5:0] GEN_798;
  wire  GEN_38;
  wire [5:0] GEN_799;
  wire  GEN_39;
  wire [5:0] GEN_800;
  wire  GEN_40;
  wire [5:0] GEN_801;
  wire  GEN_41;
  wire [5:0] GEN_802;
  wire  GEN_42;
  wire [5:0] GEN_803;
  wire  GEN_43;
  wire [5:0] GEN_804;
  wire  GEN_44;
  wire [5:0] GEN_805;
  wire  GEN_45;
  wire [5:0] GEN_806;
  wire  GEN_46;
  wire [5:0] GEN_807;
  wire  GEN_47;
  wire [5:0] GEN_808;
  wire  GEN_48;
  wire [5:0] GEN_809;
  wire  GEN_49;
  wire [5:0] GEN_810;
  wire  GEN_50;
  wire [5:0] GEN_811;
  wire  GEN_51;
  wire [5:0] GEN_812;
  wire  GEN_52;
  wire [5:0] GEN_813;
  wire  GEN_53;
  wire  GEN_54;
  wire  GEN_55;
  wire  GEN_56;
  wire  GEN_57;
  wire  GEN_58;
  wire  GEN_59;
  wire  GEN_60;
  wire  GEN_61;
  wire  GEN_62;
  wire  GEN_63;
  wire  GEN_64;
  wire  GEN_65;
  wire  GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  GEN_75;
  wire  GEN_76;
  wire  GEN_77;
  wire  GEN_78;
  wire  GEN_79;
  wire  GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_1;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire  GEN_89;
  wire  GEN_90;
  wire  GEN_91;
  wire  GEN_92;
  wire  GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_132;
  wire  GEN_133;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire [5:0] T_2881;
  wire  T_2883;
  wire  T_2884;
  wire [26:0] T_2887;
  wire  T_2888;
  wire  T_2889;
  wire  T_2892;
  wire  T_2893;
  wire  T_2896;
  wire  T_2897;
  wire  T_2900;
  wire [26:0] T_2903;
  wire  T_2904;
  wire  T_2905;
  wire  T_2908;
  wire  T_2909;
  wire  T_2912;
  wire  T_2913;
  wire [5:0] T_2916;
  wire [5:0] GEN_176;
  wire [63:0] GEN_239;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_292;
  wire  GEN_293;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_324;
  wire  GEN_325;
  wire  GEN_326;
  wire  GEN_327;
  wire  GEN_328;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_360;
  wire  GEN_361;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_393;
  wire  GEN_398;
  wire  GEN_403;
  wire  GEN_408;
  wire  GEN_413;
  wire  GEN_418;
  wire [5:0] GEN_421;
  wire [63:0] GEN_422;
  wire [5:0] GEN_423;
  wire [61:0] GEN_847;
  wire  T_2920;
  wire  T_2921;
  wire  T_2922;
  wire  T_2923;
  wire  T_2924;
  wire  T_2925;
  wire  T_2926;
  wire  T_2927;
  wire  T_2928;
  wire  T_2929;
  wire  T_2930;
  wire  T_2931;
  wire  T_2932;
  wire  T_2933;
  wire  T_2934;
  wire  T_2935;
  wire  T_2936;
  wire  T_2937;
  wire  T_2938;
  wire  T_2939;
  wire  T_2940;
  wire  T_2941;
  wire  T_2942;
  wire  T_2943;
  wire  T_2944;
  wire  T_2945;
  wire  T_2946;
  wire  T_2947;
  wire  T_2948;
  wire  T_2949;
  wire  T_2950;
  wire  T_2951;
  wire  T_2952;
  wire  T_2953;
  wire  T_2954;
  wire  T_2955;
  wire  T_2956;
  wire  T_2957;
  wire  T_2958;
  wire  T_2959;
  wire  T_2960;
  wire  T_2961;
  wire  T_2962;
  wire  T_2963;
  wire  T_2964;
  wire  T_2965;
  wire  T_2966;
  wire  T_2967;
  wire  T_2968;
  wire  T_2969;
  wire  T_2970;
  wire  T_2971;
  wire  T_2972;
  wire  T_2973;
  wire  T_2974;
  wire  T_2975;
  wire  T_2976;
  wire  T_2977;
  wire  T_2978;
  wire  T_2979;
  wire  T_2980;
  wire  T_2981;
  wire  T_2982;
  wire [5:0] T_2984;
  wire [5:0] T_2986;
  wire [5:0] T_2988;
  wire [5:0] T_2990;
  wire [5:0] T_2992;
  wire [5:0] T_2994;
  wire [5:0] T_2996;
  wire [5:0] T_2998;
  wire [5:0] T_3000;
  wire [5:0] T_3002;
  wire [5:0] T_3004;
  wire [5:0] T_3006;
  wire [5:0] T_3008;
  wire [5:0] T_3010;
  wire [5:0] T_3012;
  wire [5:0] T_3014;
  wire [5:0] T_3016;
  wire [5:0] T_3018;
  wire [5:0] T_3020;
  wire [5:0] T_3022;
  wire [5:0] T_3024;
  wire [5:0] T_3026;
  wire [5:0] T_3028;
  wire [5:0] T_3030;
  wire [5:0] T_3032;
  wire [5:0] T_3034;
  wire [5:0] T_3036;
  wire [5:0] T_3038;
  wire [5:0] T_3040;
  wire [5:0] T_3042;
  wire [5:0] T_3044;
  wire [5:0] T_3046;
  wire [5:0] T_3048;
  wire [5:0] T_3050;
  wire [5:0] T_3052;
  wire [5:0] T_3054;
  wire [5:0] T_3056;
  wire [5:0] T_3058;
  wire [5:0] T_3060;
  wire [5:0] T_3062;
  wire [5:0] T_3064;
  wire [5:0] T_3066;
  wire [5:0] T_3068;
  wire [5:0] T_3070;
  wire [5:0] T_3072;
  wire [5:0] T_3074;
  wire [5:0] T_3076;
  wire [5:0] T_3078;
  wire [5:0] T_3080;
  wire [5:0] T_3082;
  wire [5:0] T_3084;
  wire [5:0] T_3086;
  wire [5:0] T_3088;
  wire [5:0] T_3090;
  wire [5:0] T_3092;
  wire [5:0] T_3094;
  wire [5:0] T_3096;
  wire [5:0] T_3098;
  wire [5:0] T_3100;
  wire [5:0] T_3102;
  wire [5:0] T_3104;
  wire [5:0] T_3106;
  wire [5:0] T_3108;
  wire [5:0] T_3109;
  wire [5:0] T_3110;
  wire [5:0] T_3111;
  wire [5:0] T_3112;
  wire [5:0] T_3113;
  wire [5:0] T_3114;
  wire [5:0] T_3115;
  wire [5:0] T_3116;
  wire [5:0] T_3117;
  wire [5:0] T_3118;
  wire [5:0] T_3119;
  wire [5:0] T_3120;
  wire [5:0] T_3121;
  wire [5:0] T_3122;
  wire [5:0] T_3123;
  wire [5:0] T_3124;
  wire [5:0] T_3125;
  wire [5:0] T_3126;
  wire [5:0] T_3127;
  wire [5:0] T_3128;
  wire [5:0] T_3129;
  wire [5:0] T_3130;
  wire [5:0] T_3131;
  wire [5:0] T_3132;
  wire [5:0] T_3133;
  wire [5:0] T_3134;
  wire [5:0] T_3135;
  wire [5:0] T_3136;
  wire [5:0] T_3137;
  wire [5:0] T_3138;
  wire [5:0] T_3139;
  wire [5:0] T_3140;
  wire [5:0] T_3141;
  wire [5:0] T_3142;
  wire [5:0] T_3143;
  wire [5:0] T_3144;
  wire [5:0] T_3145;
  wire [5:0] T_3146;
  wire [5:0] T_3147;
  wire [5:0] T_3148;
  wire [5:0] T_3149;
  wire [5:0] T_3150;
  wire [5:0] T_3151;
  wire [5:0] T_3152;
  wire [5:0] T_3153;
  wire [5:0] T_3154;
  wire [5:0] T_3155;
  wire [5:0] T_3156;
  wire [5:0] T_3157;
  wire [5:0] T_3158;
  wire [5:0] T_3159;
  wire [5:0] T_3160;
  wire [5:0] T_3161;
  wire [5:0] T_3162;
  wire [5:0] T_3163;
  wire [5:0] T_3164;
  wire [5:0] T_3165;
  wire [5:0] T_3166;
  wire [5:0] T_3167;
  wire [5:0] T_3168;
  wire [5:0] T_3169;
  wire  T_3170;
  wire  T_3171;
  wire  T_3172;
  wire  T_3173;
  wire  T_3174;
  wire  T_3175;
  wire [26:0] T_3189;
  wire [26:0] T_3191;
  wire [26:0] T_3193;
  wire [26:0] T_3195;
  wire [26:0] T_3197;
  wire [26:0] T_3199;
  wire [26:0] T_3201;
  wire [26:0] T_3202;
  wire [26:0] T_3203;
  wire [26:0] T_3204;
  wire [26:0] T_3205;
  wire [26:0] T_3206;
  wire [11:0] T_3394;
  wire [11:0] T_3396;
  wire [11:0] T_3398;
  wire [11:0] T_3400;
  wire [11:0] T_3402;
  wire [11:0] T_3404;
  wire [11:0] T_3406;
  wire [11:0] T_3408;
  wire [11:0] T_3410;
  wire [11:0] T_3412;
  wire [11:0] T_3414;
  wire [11:0] T_3416;
  wire [11:0] T_3418;
  wire [11:0] T_3420;
  wire [11:0] T_3422;
  wire [11:0] T_3424;
  wire [11:0] T_3426;
  wire [11:0] T_3428;
  wire [11:0] T_3430;
  wire [11:0] T_3432;
  wire [11:0] T_3434;
  wire [11:0] T_3436;
  wire [11:0] T_3438;
  wire [11:0] T_3440;
  wire [11:0] T_3442;
  wire [11:0] T_3444;
  wire [11:0] T_3446;
  wire [11:0] T_3448;
  wire [11:0] T_3450;
  wire [11:0] T_3452;
  wire [11:0] T_3454;
  wire [11:0] T_3456;
  wire [11:0] T_3458;
  wire [11:0] T_3460;
  wire [11:0] T_3462;
  wire [11:0] T_3464;
  wire [11:0] T_3466;
  wire [11:0] T_3468;
  wire [11:0] T_3470;
  wire [11:0] T_3472;
  wire [11:0] T_3474;
  wire [11:0] T_3476;
  wire [11:0] T_3478;
  wire [11:0] T_3480;
  wire [11:0] T_3482;
  wire [11:0] T_3484;
  wire [11:0] T_3486;
  wire [11:0] T_3488;
  wire [11:0] T_3490;
  wire [11:0] T_3492;
  wire [11:0] T_3494;
  wire [11:0] T_3496;
  wire [11:0] T_3498;
  wire [11:0] T_3500;
  wire [11:0] T_3502;
  wire [11:0] T_3504;
  wire [11:0] T_3506;
  wire [11:0] T_3508;
  wire [11:0] T_3510;
  wire [11:0] T_3512;
  wire [11:0] T_3514;
  wire [11:0] T_3516;
  wire [11:0] T_3518;
  wire [11:0] T_3519;
  wire [11:0] T_3520;
  wire [11:0] T_3521;
  wire [11:0] T_3522;
  wire [11:0] T_3523;
  wire [11:0] T_3524;
  wire [11:0] T_3525;
  wire [11:0] T_3526;
  wire [11:0] T_3527;
  wire [11:0] T_3528;
  wire [11:0] T_3529;
  wire [11:0] T_3530;
  wire [11:0] T_3531;
  wire [11:0] T_3532;
  wire [11:0] T_3533;
  wire [11:0] T_3534;
  wire [11:0] T_3535;
  wire [11:0] T_3536;
  wire [11:0] T_3537;
  wire [11:0] T_3538;
  wire [11:0] T_3539;
  wire [11:0] T_3540;
  wire [11:0] T_3541;
  wire [11:0] T_3542;
  wire [11:0] T_3543;
  wire [11:0] T_3544;
  wire [11:0] T_3545;
  wire [11:0] T_3546;
  wire [11:0] T_3547;
  wire [11:0] T_3548;
  wire [11:0] T_3549;
  wire [11:0] T_3550;
  wire [11:0] T_3551;
  wire [11:0] T_3552;
  wire [11:0] T_3553;
  wire [11:0] T_3554;
  wire [11:0] T_3555;
  wire [11:0] T_3556;
  wire [11:0] T_3557;
  wire [11:0] T_3558;
  wire [11:0] T_3559;
  wire [11:0] T_3560;
  wire [11:0] T_3561;
  wire [11:0] T_3562;
  wire [11:0] T_3563;
  wire [11:0] T_3564;
  wire [11:0] T_3565;
  wire [11:0] T_3566;
  wire [11:0] T_3567;
  wire [11:0] T_3568;
  wire [11:0] T_3569;
  wire [11:0] T_3570;
  wire [11:0] T_3571;
  wire [11:0] T_3572;
  wire [11:0] T_3573;
  wire [11:0] T_3574;
  wire [11:0] T_3575;
  wire [11:0] T_3576;
  wire [11:0] T_3577;
  wire [11:0] T_3578;
  wire [11:0] T_3579;
  wire [38:0] T_3580;
  wire [29:0] T_3581;
  wire [31:0] T_3582;
  wire [29:0] GEN_848;
  wire  T_3584;
  wire [31:0] GEN_849;
  wire [31:0] T_3585;
  wire [15:0] T_3586;
  wire [15:0] T_3587;
  wire [15:0] GEN_850;
  wire  T_3589;
  wire [15:0] T_3590;
  wire [7:0] T_3591;
  wire [7:0] T_3592;
  wire [7:0] GEN_851;
  wire  T_3594;
  wire [7:0] T_3595;
  wire [3:0] T_3596;
  wire [3:0] T_3597;
  wire [3:0] GEN_852;
  wire  T_3599;
  wire [3:0] T_3600;
  wire [1:0] T_3601;
  wire [1:0] T_3602;
  wire  T_3604;
  wire [1:0] T_3605;
  wire  T_3606;
  wire [1:0] T_3607;
  wire [2:0] T_3608;
  wire [3:0] T_3609;
  wire [4:0] T_3610;
  wire [5:0] T_3611;
  reg [1:0] T_3616 [0:127];
  reg [31:0] GEN_441;
  wire [1:0] T_3616_T_3942_data;
  wire [6:0] T_3616_T_3942_addr;
  wire  T_3616_T_3942_en;
  wire [1:0] T_3616_T_3949_data;
  wire [6:0] T_3616_T_3949_addr;
  wire  T_3616_T_3949_mask;
  wire  T_3616_T_3949_en;
  reg [6:0] T_3618;
  reg [31:0] GEN_451;
  wire  T_3683;
  wire  T_3686;
  wire  T_3689;
  wire  T_3692;
  wire  T_3695;
  wire  T_3698;
  wire  T_3701;
  wire  T_3704;
  wire  T_3707;
  wire  T_3710;
  wire  T_3713;
  wire  T_3716;
  wire  T_3719;
  wire  T_3722;
  wire  T_3725;
  wire  T_3728;
  wire  T_3731;
  wire  T_3734;
  wire  T_3737;
  wire  T_3740;
  wire  T_3743;
  wire  T_3746;
  wire  T_3749;
  wire  T_3752;
  wire  T_3755;
  wire  T_3758;
  wire  T_3761;
  wire  T_3764;
  wire  T_3767;
  wire  T_3770;
  wire  T_3773;
  wire  T_3776;
  wire  T_3779;
  wire  T_3782;
  wire  T_3785;
  wire  T_3788;
  wire  T_3791;
  wire  T_3794;
  wire  T_3797;
  wire  T_3800;
  wire  T_3803;
  wire  T_3806;
  wire  T_3809;
  wire  T_3812;
  wire  T_3815;
  wire  T_3818;
  wire  T_3821;
  wire  T_3824;
  wire  T_3827;
  wire  T_3830;
  wire  T_3833;
  wire  T_3836;
  wire  T_3839;
  wire  T_3842;
  wire  T_3845;
  wire  T_3848;
  wire  T_3851;
  wire  T_3854;
  wire  T_3857;
  wire  T_3860;
  wire  T_3863;
  wire  T_3866;
  wire  T_3868;
  wire  T_3869;
  wire  T_3870;
  wire  T_3871;
  wire  T_3872;
  wire  T_3873;
  wire  T_3874;
  wire  T_3875;
  wire  T_3876;
  wire  T_3877;
  wire  T_3878;
  wire  T_3879;
  wire  T_3880;
  wire  T_3881;
  wire  T_3882;
  wire  T_3883;
  wire  T_3884;
  wire  T_3885;
  wire  T_3886;
  wire  T_3887;
  wire  T_3888;
  wire  T_3889;
  wire  T_3890;
  wire  T_3891;
  wire  T_3892;
  wire  T_3893;
  wire  T_3894;
  wire  T_3895;
  wire  T_3896;
  wire  T_3897;
  wire  T_3898;
  wire  T_3899;
  wire  T_3900;
  wire  T_3901;
  wire  T_3902;
  wire  T_3903;
  wire  T_3904;
  wire  T_3905;
  wire  T_3906;
  wire  T_3907;
  wire  T_3908;
  wire  T_3909;
  wire  T_3910;
  wire  T_3911;
  wire  T_3912;
  wire  T_3913;
  wire  T_3914;
  wire  T_3915;
  wire  T_3916;
  wire  T_3917;
  wire  T_3918;
  wire  T_3919;
  wire  T_3920;
  wire  T_3921;
  wire  T_3922;
  wire  T_3923;
  wire  T_3924;
  wire  T_3925;
  wire  T_3926;
  wire  T_3927;
  wire  T_3928;
  wire  T_3929;
  wire  T_3931;
  wire  T_3932;
  wire  T_3933;
  wire [6:0] T_3937_history;
  wire [1:0] T_3937_value;
  wire [6:0] T_3940;
  wire [6:0] T_3941;
  wire  T_3943;
  wire [5:0] T_3944;
  wire [6:0] T_3945;
  wire [6:0] GEN_424;
  wire  T_3946;
  wire [6:0] T_3947;
  wire [6:0] T_3948;
  wire  T_3950;
  wire  T_3951;
  wire  T_3952;
  wire  T_3955;
  wire  T_3956;
  wire  T_3957;
  wire [1:0] T_3958;
  wire [5:0] T_3959;
  wire [6:0] T_3960;
  wire [6:0] GEN_425;
  wire [6:0] GEN_431;
  wire  T_3963;
  wire  T_3964;
  wire  GEN_432;
  reg [1:0] T_3967;
  reg [31:0] GEN_458;
  reg  T_3969;
  reg [31:0] GEN_459;
  reg [38:0] T_3976_0;
  reg [63:0] GEN_460;
  reg [38:0] T_3976_1;
  reg [63:0] GEN_461;
  wire  T_4042;
  wire  T_4045;
  wire  T_4048;
  wire  T_4051;
  wire  T_4054;
  wire  T_4057;
  wire  T_4060;
  wire  T_4063;
  wire  T_4066;
  wire  T_4069;
  wire  T_4072;
  wire  T_4075;
  wire  T_4078;
  wire  T_4081;
  wire  T_4084;
  wire  T_4087;
  wire  T_4090;
  wire  T_4093;
  wire  T_4096;
  wire  T_4099;
  wire  T_4102;
  wire  T_4105;
  wire  T_4108;
  wire  T_4111;
  wire  T_4114;
  wire  T_4117;
  wire  T_4120;
  wire  T_4123;
  wire  T_4126;
  wire  T_4129;
  wire  T_4132;
  wire  T_4135;
  wire  T_4138;
  wire  T_4141;
  wire  T_4144;
  wire  T_4147;
  wire  T_4150;
  wire  T_4153;
  wire  T_4156;
  wire  T_4159;
  wire  T_4162;
  wire  T_4165;
  wire  T_4168;
  wire  T_4171;
  wire  T_4174;
  wire  T_4177;
  wire  T_4180;
  wire  T_4183;
  wire  T_4186;
  wire  T_4189;
  wire  T_4192;
  wire  T_4195;
  wire  T_4198;
  wire  T_4201;
  wire  T_4204;
  wire  T_4207;
  wire  T_4210;
  wire  T_4213;
  wire  T_4216;
  wire  T_4219;
  wire  T_4222;
  wire  T_4225;
  wire  T_4227;
  wire  T_4228;
  wire  T_4229;
  wire  T_4230;
  wire  T_4231;
  wire  T_4232;
  wire  T_4233;
  wire  T_4234;
  wire  T_4235;
  wire  T_4236;
  wire  T_4237;
  wire  T_4238;
  wire  T_4239;
  wire  T_4240;
  wire  T_4241;
  wire  T_4242;
  wire  T_4243;
  wire  T_4244;
  wire  T_4245;
  wire  T_4246;
  wire  T_4247;
  wire  T_4248;
  wire  T_4249;
  wire  T_4250;
  wire  T_4251;
  wire  T_4252;
  wire  T_4253;
  wire  T_4254;
  wire  T_4255;
  wire  T_4256;
  wire  T_4257;
  wire  T_4258;
  wire  T_4259;
  wire  T_4260;
  wire  T_4261;
  wire  T_4262;
  wire  T_4263;
  wire  T_4264;
  wire  T_4265;
  wire  T_4266;
  wire  T_4267;
  wire  T_4268;
  wire  T_4269;
  wire  T_4270;
  wire  T_4271;
  wire  T_4272;
  wire  T_4273;
  wire  T_4274;
  wire  T_4275;
  wire  T_4276;
  wire  T_4277;
  wire  T_4278;
  wire  T_4279;
  wire  T_4280;
  wire  T_4281;
  wire  T_4282;
  wire  T_4283;
  wire  T_4284;
  wire  T_4285;
  wire  T_4286;
  wire  T_4287;
  wire  T_4288;
  wire  T_4290;
  wire  T_4292;
  wire  T_4293;
  wire [38:0] GEN_2;
  wire [38:0] GEN_433;
  wire [38:0] GEN_435;
  wire  T_4295;
  wire [1:0] GEN_855;
  wire [2:0] T_4297;
  wire [1:0] T_4298;
  wire [1:0] GEN_436;
  wire [1:0] T_4304;
  wire  T_4305;
  wire [38:0] GEN_3;
  wire [38:0] GEN_437;
  wire [38:0] GEN_438;
  wire [38:0] GEN_439;
  wire [1:0] GEN_440;
  wire [38:0] GEN_442;
  wire [38:0] GEN_443;
  wire  GEN_444;
  wire [38:0] GEN_445;
  wire  T_4308;
  wire  T_4310;
  wire  T_4311;
  wire [2:0] T_4317;
  wire [1:0] T_4318;
  wire [1:0] T_4324;
  wire  T_4325;
  wire [1:0] GEN_446;
  wire  GEN_447;
  wire [1:0] GEN_448;
  wire  GEN_449;
  wire [1:0] GEN_450;
  wire [38:0] GEN_452;
  wire [38:0] GEN_453;
  wire  GEN_454;
  wire [38:0] GEN_455;
  wire [1:0] GEN_456;
  assign io_resp_valid = T_2920;
  assign io_resp_bits_taken = GEN_432;
  assign io_resp_bits_mask = 1'h1;
  assign io_resp_bits_bridx = brIdx_T_3612_data;
  assign io_resp_bits_target = GEN_455;
  assign io_resp_bits_entry = T_3611;
  assign io_resp_bits_bht_history = T_3937_history;
  assign io_resp_bits_bht_value = T_3937_value;
  assign idxs_T_1431_addr = {{5'd0}, 1'h0};
  assign idxs_T_1431_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1431_data = idxs[idxs_T_1431_addr];
  `else
  assign idxs_T_1431_data = idxs_T_1431_addr >= 6'h3e ? $random : idxs[idxs_T_1431_addr];
  `endif
  assign idxs_T_1434_addr = {{5'd0}, 1'h1};
  assign idxs_T_1434_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1434_data = idxs[idxs_T_1434_addr];
  `else
  assign idxs_T_1434_data = idxs_T_1434_addr >= 6'h3e ? $random : idxs[idxs_T_1434_addr];
  `endif
  assign idxs_T_1437_addr = {{4'd0}, 2'h2};
  assign idxs_T_1437_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1437_data = idxs[idxs_T_1437_addr];
  `else
  assign idxs_T_1437_data = idxs_T_1437_addr >= 6'h3e ? $random : idxs[idxs_T_1437_addr];
  `endif
  assign idxs_T_1440_addr = {{4'd0}, 2'h3};
  assign idxs_T_1440_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1440_data = idxs[idxs_T_1440_addr];
  `else
  assign idxs_T_1440_data = idxs_T_1440_addr >= 6'h3e ? $random : idxs[idxs_T_1440_addr];
  `endif
  assign idxs_T_1443_addr = {{3'd0}, 3'h4};
  assign idxs_T_1443_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1443_data = idxs[idxs_T_1443_addr];
  `else
  assign idxs_T_1443_data = idxs_T_1443_addr >= 6'h3e ? $random : idxs[idxs_T_1443_addr];
  `endif
  assign idxs_T_1446_addr = {{3'd0}, 3'h5};
  assign idxs_T_1446_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1446_data = idxs[idxs_T_1446_addr];
  `else
  assign idxs_T_1446_data = idxs_T_1446_addr >= 6'h3e ? $random : idxs[idxs_T_1446_addr];
  `endif
  assign idxs_T_1449_addr = {{3'd0}, 3'h6};
  assign idxs_T_1449_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1449_data = idxs[idxs_T_1449_addr];
  `else
  assign idxs_T_1449_data = idxs_T_1449_addr >= 6'h3e ? $random : idxs[idxs_T_1449_addr];
  `endif
  assign idxs_T_1452_addr = {{3'd0}, 3'h7};
  assign idxs_T_1452_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1452_data = idxs[idxs_T_1452_addr];
  `else
  assign idxs_T_1452_data = idxs_T_1452_addr >= 6'h3e ? $random : idxs[idxs_T_1452_addr];
  `endif
  assign idxs_T_1455_addr = {{2'd0}, 4'h8};
  assign idxs_T_1455_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1455_data = idxs[idxs_T_1455_addr];
  `else
  assign idxs_T_1455_data = idxs_T_1455_addr >= 6'h3e ? $random : idxs[idxs_T_1455_addr];
  `endif
  assign idxs_T_1458_addr = {{2'd0}, 4'h9};
  assign idxs_T_1458_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1458_data = idxs[idxs_T_1458_addr];
  `else
  assign idxs_T_1458_data = idxs_T_1458_addr >= 6'h3e ? $random : idxs[idxs_T_1458_addr];
  `endif
  assign idxs_T_1461_addr = {{2'd0}, 4'ha};
  assign idxs_T_1461_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1461_data = idxs[idxs_T_1461_addr];
  `else
  assign idxs_T_1461_data = idxs_T_1461_addr >= 6'h3e ? $random : idxs[idxs_T_1461_addr];
  `endif
  assign idxs_T_1464_addr = {{2'd0}, 4'hb};
  assign idxs_T_1464_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1464_data = idxs[idxs_T_1464_addr];
  `else
  assign idxs_T_1464_data = idxs_T_1464_addr >= 6'h3e ? $random : idxs[idxs_T_1464_addr];
  `endif
  assign idxs_T_1467_addr = {{2'd0}, 4'hc};
  assign idxs_T_1467_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1467_data = idxs[idxs_T_1467_addr];
  `else
  assign idxs_T_1467_data = idxs_T_1467_addr >= 6'h3e ? $random : idxs[idxs_T_1467_addr];
  `endif
  assign idxs_T_1470_addr = {{2'd0}, 4'hd};
  assign idxs_T_1470_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1470_data = idxs[idxs_T_1470_addr];
  `else
  assign idxs_T_1470_data = idxs_T_1470_addr >= 6'h3e ? $random : idxs[idxs_T_1470_addr];
  `endif
  assign idxs_T_1473_addr = {{2'd0}, 4'he};
  assign idxs_T_1473_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1473_data = idxs[idxs_T_1473_addr];
  `else
  assign idxs_T_1473_data = idxs_T_1473_addr >= 6'h3e ? $random : idxs[idxs_T_1473_addr];
  `endif
  assign idxs_T_1476_addr = {{2'd0}, 4'hf};
  assign idxs_T_1476_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1476_data = idxs[idxs_T_1476_addr];
  `else
  assign idxs_T_1476_data = idxs_T_1476_addr >= 6'h3e ? $random : idxs[idxs_T_1476_addr];
  `endif
  assign idxs_T_1479_addr = {{1'd0}, 5'h10};
  assign idxs_T_1479_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1479_data = idxs[idxs_T_1479_addr];
  `else
  assign idxs_T_1479_data = idxs_T_1479_addr >= 6'h3e ? $random : idxs[idxs_T_1479_addr];
  `endif
  assign idxs_T_1482_addr = {{1'd0}, 5'h11};
  assign idxs_T_1482_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1482_data = idxs[idxs_T_1482_addr];
  `else
  assign idxs_T_1482_data = idxs_T_1482_addr >= 6'h3e ? $random : idxs[idxs_T_1482_addr];
  `endif
  assign idxs_T_1485_addr = {{1'd0}, 5'h12};
  assign idxs_T_1485_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1485_data = idxs[idxs_T_1485_addr];
  `else
  assign idxs_T_1485_data = idxs_T_1485_addr >= 6'h3e ? $random : idxs[idxs_T_1485_addr];
  `endif
  assign idxs_T_1488_addr = {{1'd0}, 5'h13};
  assign idxs_T_1488_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1488_data = idxs[idxs_T_1488_addr];
  `else
  assign idxs_T_1488_data = idxs_T_1488_addr >= 6'h3e ? $random : idxs[idxs_T_1488_addr];
  `endif
  assign idxs_T_1491_addr = {{1'd0}, 5'h14};
  assign idxs_T_1491_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1491_data = idxs[idxs_T_1491_addr];
  `else
  assign idxs_T_1491_data = idxs_T_1491_addr >= 6'h3e ? $random : idxs[idxs_T_1491_addr];
  `endif
  assign idxs_T_1494_addr = {{1'd0}, 5'h15};
  assign idxs_T_1494_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1494_data = idxs[idxs_T_1494_addr];
  `else
  assign idxs_T_1494_data = idxs_T_1494_addr >= 6'h3e ? $random : idxs[idxs_T_1494_addr];
  `endif
  assign idxs_T_1497_addr = {{1'd0}, 5'h16};
  assign idxs_T_1497_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1497_data = idxs[idxs_T_1497_addr];
  `else
  assign idxs_T_1497_data = idxs_T_1497_addr >= 6'h3e ? $random : idxs[idxs_T_1497_addr];
  `endif
  assign idxs_T_1500_addr = {{1'd0}, 5'h17};
  assign idxs_T_1500_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1500_data = idxs[idxs_T_1500_addr];
  `else
  assign idxs_T_1500_data = idxs_T_1500_addr >= 6'h3e ? $random : idxs[idxs_T_1500_addr];
  `endif
  assign idxs_T_1503_addr = {{1'd0}, 5'h18};
  assign idxs_T_1503_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1503_data = idxs[idxs_T_1503_addr];
  `else
  assign idxs_T_1503_data = idxs_T_1503_addr >= 6'h3e ? $random : idxs[idxs_T_1503_addr];
  `endif
  assign idxs_T_1506_addr = {{1'd0}, 5'h19};
  assign idxs_T_1506_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1506_data = idxs[idxs_T_1506_addr];
  `else
  assign idxs_T_1506_data = idxs_T_1506_addr >= 6'h3e ? $random : idxs[idxs_T_1506_addr];
  `endif
  assign idxs_T_1509_addr = {{1'd0}, 5'h1a};
  assign idxs_T_1509_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1509_data = idxs[idxs_T_1509_addr];
  `else
  assign idxs_T_1509_data = idxs_T_1509_addr >= 6'h3e ? $random : idxs[idxs_T_1509_addr];
  `endif
  assign idxs_T_1512_addr = {{1'd0}, 5'h1b};
  assign idxs_T_1512_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1512_data = idxs[idxs_T_1512_addr];
  `else
  assign idxs_T_1512_data = idxs_T_1512_addr >= 6'h3e ? $random : idxs[idxs_T_1512_addr];
  `endif
  assign idxs_T_1515_addr = {{1'd0}, 5'h1c};
  assign idxs_T_1515_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1515_data = idxs[idxs_T_1515_addr];
  `else
  assign idxs_T_1515_data = idxs_T_1515_addr >= 6'h3e ? $random : idxs[idxs_T_1515_addr];
  `endif
  assign idxs_T_1518_addr = {{1'd0}, 5'h1d};
  assign idxs_T_1518_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1518_data = idxs[idxs_T_1518_addr];
  `else
  assign idxs_T_1518_data = idxs_T_1518_addr >= 6'h3e ? $random : idxs[idxs_T_1518_addr];
  `endif
  assign idxs_T_1521_addr = {{1'd0}, 5'h1e};
  assign idxs_T_1521_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1521_data = idxs[idxs_T_1521_addr];
  `else
  assign idxs_T_1521_data = idxs_T_1521_addr >= 6'h3e ? $random : idxs[idxs_T_1521_addr];
  `endif
  assign idxs_T_1524_addr = {{1'd0}, 5'h1f};
  assign idxs_T_1524_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1524_data = idxs[idxs_T_1524_addr];
  `else
  assign idxs_T_1524_data = idxs_T_1524_addr >= 6'h3e ? $random : idxs[idxs_T_1524_addr];
  `endif
  assign idxs_T_1527_addr = 6'h20;
  assign idxs_T_1527_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1527_data = idxs[idxs_T_1527_addr];
  `else
  assign idxs_T_1527_data = idxs_T_1527_addr >= 6'h3e ? $random : idxs[idxs_T_1527_addr];
  `endif
  assign idxs_T_1530_addr = 6'h21;
  assign idxs_T_1530_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1530_data = idxs[idxs_T_1530_addr];
  `else
  assign idxs_T_1530_data = idxs_T_1530_addr >= 6'h3e ? $random : idxs[idxs_T_1530_addr];
  `endif
  assign idxs_T_1533_addr = 6'h22;
  assign idxs_T_1533_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1533_data = idxs[idxs_T_1533_addr];
  `else
  assign idxs_T_1533_data = idxs_T_1533_addr >= 6'h3e ? $random : idxs[idxs_T_1533_addr];
  `endif
  assign idxs_T_1536_addr = 6'h23;
  assign idxs_T_1536_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1536_data = idxs[idxs_T_1536_addr];
  `else
  assign idxs_T_1536_data = idxs_T_1536_addr >= 6'h3e ? $random : idxs[idxs_T_1536_addr];
  `endif
  assign idxs_T_1539_addr = 6'h24;
  assign idxs_T_1539_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1539_data = idxs[idxs_T_1539_addr];
  `else
  assign idxs_T_1539_data = idxs_T_1539_addr >= 6'h3e ? $random : idxs[idxs_T_1539_addr];
  `endif
  assign idxs_T_1542_addr = 6'h25;
  assign idxs_T_1542_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1542_data = idxs[idxs_T_1542_addr];
  `else
  assign idxs_T_1542_data = idxs_T_1542_addr >= 6'h3e ? $random : idxs[idxs_T_1542_addr];
  `endif
  assign idxs_T_1545_addr = 6'h26;
  assign idxs_T_1545_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1545_data = idxs[idxs_T_1545_addr];
  `else
  assign idxs_T_1545_data = idxs_T_1545_addr >= 6'h3e ? $random : idxs[idxs_T_1545_addr];
  `endif
  assign idxs_T_1548_addr = 6'h27;
  assign idxs_T_1548_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1548_data = idxs[idxs_T_1548_addr];
  `else
  assign idxs_T_1548_data = idxs_T_1548_addr >= 6'h3e ? $random : idxs[idxs_T_1548_addr];
  `endif
  assign idxs_T_1551_addr = 6'h28;
  assign idxs_T_1551_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1551_data = idxs[idxs_T_1551_addr];
  `else
  assign idxs_T_1551_data = idxs_T_1551_addr >= 6'h3e ? $random : idxs[idxs_T_1551_addr];
  `endif
  assign idxs_T_1554_addr = 6'h29;
  assign idxs_T_1554_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1554_data = idxs[idxs_T_1554_addr];
  `else
  assign idxs_T_1554_data = idxs_T_1554_addr >= 6'h3e ? $random : idxs[idxs_T_1554_addr];
  `endif
  assign idxs_T_1557_addr = 6'h2a;
  assign idxs_T_1557_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1557_data = idxs[idxs_T_1557_addr];
  `else
  assign idxs_T_1557_data = idxs_T_1557_addr >= 6'h3e ? $random : idxs[idxs_T_1557_addr];
  `endif
  assign idxs_T_1560_addr = 6'h2b;
  assign idxs_T_1560_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1560_data = idxs[idxs_T_1560_addr];
  `else
  assign idxs_T_1560_data = idxs_T_1560_addr >= 6'h3e ? $random : idxs[idxs_T_1560_addr];
  `endif
  assign idxs_T_1563_addr = 6'h2c;
  assign idxs_T_1563_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1563_data = idxs[idxs_T_1563_addr];
  `else
  assign idxs_T_1563_data = idxs_T_1563_addr >= 6'h3e ? $random : idxs[idxs_T_1563_addr];
  `endif
  assign idxs_T_1566_addr = 6'h2d;
  assign idxs_T_1566_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1566_data = idxs[idxs_T_1566_addr];
  `else
  assign idxs_T_1566_data = idxs_T_1566_addr >= 6'h3e ? $random : idxs[idxs_T_1566_addr];
  `endif
  assign idxs_T_1569_addr = 6'h2e;
  assign idxs_T_1569_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1569_data = idxs[idxs_T_1569_addr];
  `else
  assign idxs_T_1569_data = idxs_T_1569_addr >= 6'h3e ? $random : idxs[idxs_T_1569_addr];
  `endif
  assign idxs_T_1572_addr = 6'h2f;
  assign idxs_T_1572_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1572_data = idxs[idxs_T_1572_addr];
  `else
  assign idxs_T_1572_data = idxs_T_1572_addr >= 6'h3e ? $random : idxs[idxs_T_1572_addr];
  `endif
  assign idxs_T_1575_addr = 6'h30;
  assign idxs_T_1575_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1575_data = idxs[idxs_T_1575_addr];
  `else
  assign idxs_T_1575_data = idxs_T_1575_addr >= 6'h3e ? $random : idxs[idxs_T_1575_addr];
  `endif
  assign idxs_T_1578_addr = 6'h31;
  assign idxs_T_1578_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1578_data = idxs[idxs_T_1578_addr];
  `else
  assign idxs_T_1578_data = idxs_T_1578_addr >= 6'h3e ? $random : idxs[idxs_T_1578_addr];
  `endif
  assign idxs_T_1581_addr = 6'h32;
  assign idxs_T_1581_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1581_data = idxs[idxs_T_1581_addr];
  `else
  assign idxs_T_1581_data = idxs_T_1581_addr >= 6'h3e ? $random : idxs[idxs_T_1581_addr];
  `endif
  assign idxs_T_1584_addr = 6'h33;
  assign idxs_T_1584_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1584_data = idxs[idxs_T_1584_addr];
  `else
  assign idxs_T_1584_data = idxs_T_1584_addr >= 6'h3e ? $random : idxs[idxs_T_1584_addr];
  `endif
  assign idxs_T_1587_addr = 6'h34;
  assign idxs_T_1587_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1587_data = idxs[idxs_T_1587_addr];
  `else
  assign idxs_T_1587_data = idxs_T_1587_addr >= 6'h3e ? $random : idxs[idxs_T_1587_addr];
  `endif
  assign idxs_T_1590_addr = 6'h35;
  assign idxs_T_1590_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1590_data = idxs[idxs_T_1590_addr];
  `else
  assign idxs_T_1590_data = idxs_T_1590_addr >= 6'h3e ? $random : idxs[idxs_T_1590_addr];
  `endif
  assign idxs_T_1593_addr = 6'h36;
  assign idxs_T_1593_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1593_data = idxs[idxs_T_1593_addr];
  `else
  assign idxs_T_1593_data = idxs_T_1593_addr >= 6'h3e ? $random : idxs[idxs_T_1593_addr];
  `endif
  assign idxs_T_1596_addr = 6'h37;
  assign idxs_T_1596_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1596_data = idxs[idxs_T_1596_addr];
  `else
  assign idxs_T_1596_data = idxs_T_1596_addr >= 6'h3e ? $random : idxs[idxs_T_1596_addr];
  `endif
  assign idxs_T_1599_addr = 6'h38;
  assign idxs_T_1599_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1599_data = idxs[idxs_T_1599_addr];
  `else
  assign idxs_T_1599_data = idxs_T_1599_addr >= 6'h3e ? $random : idxs[idxs_T_1599_addr];
  `endif
  assign idxs_T_1602_addr = 6'h39;
  assign idxs_T_1602_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1602_data = idxs[idxs_T_1602_addr];
  `else
  assign idxs_T_1602_data = idxs_T_1602_addr >= 6'h3e ? $random : idxs[idxs_T_1602_addr];
  `endif
  assign idxs_T_1605_addr = 6'h3a;
  assign idxs_T_1605_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1605_data = idxs[idxs_T_1605_addr];
  `else
  assign idxs_T_1605_data = idxs_T_1605_addr >= 6'h3e ? $random : idxs[idxs_T_1605_addr];
  `endif
  assign idxs_T_1608_addr = 6'h3b;
  assign idxs_T_1608_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1608_data = idxs[idxs_T_1608_addr];
  `else
  assign idxs_T_1608_data = idxs_T_1608_addr >= 6'h3e ? $random : idxs[idxs_T_1608_addr];
  `endif
  assign idxs_T_1611_addr = 6'h3c;
  assign idxs_T_1611_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1611_data = idxs[idxs_T_1611_addr];
  `else
  assign idxs_T_1611_data = idxs_T_1611_addr >= 6'h3e ? $random : idxs[idxs_T_1611_addr];
  `endif
  assign idxs_T_1614_addr = 6'h3d;
  assign idxs_T_1614_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1614_data = idxs[idxs_T_1614_addr];
  `else
  assign idxs_T_1614_data = idxs_T_1614_addr >= 6'h3e ? $random : idxs[idxs_T_1614_addr];
  `endif
  assign idxs_T_1972_addr = {{5'd0}, 1'h0};
  assign idxs_T_1972_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1972_data = idxs[idxs_T_1972_addr];
  `else
  assign idxs_T_1972_data = idxs_T_1972_addr >= 6'h3e ? $random : idxs[idxs_T_1972_addr];
  `endif
  assign idxs_T_1975_addr = {{5'd0}, 1'h1};
  assign idxs_T_1975_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1975_data = idxs[idxs_T_1975_addr];
  `else
  assign idxs_T_1975_data = idxs_T_1975_addr >= 6'h3e ? $random : idxs[idxs_T_1975_addr];
  `endif
  assign idxs_T_1978_addr = {{4'd0}, 2'h2};
  assign idxs_T_1978_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1978_data = idxs[idxs_T_1978_addr];
  `else
  assign idxs_T_1978_data = idxs_T_1978_addr >= 6'h3e ? $random : idxs[idxs_T_1978_addr];
  `endif
  assign idxs_T_1981_addr = {{4'd0}, 2'h3};
  assign idxs_T_1981_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1981_data = idxs[idxs_T_1981_addr];
  `else
  assign idxs_T_1981_data = idxs_T_1981_addr >= 6'h3e ? $random : idxs[idxs_T_1981_addr];
  `endif
  assign idxs_T_1984_addr = {{3'd0}, 3'h4};
  assign idxs_T_1984_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1984_data = idxs[idxs_T_1984_addr];
  `else
  assign idxs_T_1984_data = idxs_T_1984_addr >= 6'h3e ? $random : idxs[idxs_T_1984_addr];
  `endif
  assign idxs_T_1987_addr = {{3'd0}, 3'h5};
  assign idxs_T_1987_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1987_data = idxs[idxs_T_1987_addr];
  `else
  assign idxs_T_1987_data = idxs_T_1987_addr >= 6'h3e ? $random : idxs[idxs_T_1987_addr];
  `endif
  assign idxs_T_1990_addr = {{3'd0}, 3'h6};
  assign idxs_T_1990_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1990_data = idxs[idxs_T_1990_addr];
  `else
  assign idxs_T_1990_data = idxs_T_1990_addr >= 6'h3e ? $random : idxs[idxs_T_1990_addr];
  `endif
  assign idxs_T_1993_addr = {{3'd0}, 3'h7};
  assign idxs_T_1993_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1993_data = idxs[idxs_T_1993_addr];
  `else
  assign idxs_T_1993_data = idxs_T_1993_addr >= 6'h3e ? $random : idxs[idxs_T_1993_addr];
  `endif
  assign idxs_T_1996_addr = {{2'd0}, 4'h8};
  assign idxs_T_1996_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1996_data = idxs[idxs_T_1996_addr];
  `else
  assign idxs_T_1996_data = idxs_T_1996_addr >= 6'h3e ? $random : idxs[idxs_T_1996_addr];
  `endif
  assign idxs_T_1999_addr = {{2'd0}, 4'h9};
  assign idxs_T_1999_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_1999_data = idxs[idxs_T_1999_addr];
  `else
  assign idxs_T_1999_data = idxs_T_1999_addr >= 6'h3e ? $random : idxs[idxs_T_1999_addr];
  `endif
  assign idxs_T_2002_addr = {{2'd0}, 4'ha};
  assign idxs_T_2002_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2002_data = idxs[idxs_T_2002_addr];
  `else
  assign idxs_T_2002_data = idxs_T_2002_addr >= 6'h3e ? $random : idxs[idxs_T_2002_addr];
  `endif
  assign idxs_T_2005_addr = {{2'd0}, 4'hb};
  assign idxs_T_2005_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2005_data = idxs[idxs_T_2005_addr];
  `else
  assign idxs_T_2005_data = idxs_T_2005_addr >= 6'h3e ? $random : idxs[idxs_T_2005_addr];
  `endif
  assign idxs_T_2008_addr = {{2'd0}, 4'hc};
  assign idxs_T_2008_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2008_data = idxs[idxs_T_2008_addr];
  `else
  assign idxs_T_2008_data = idxs_T_2008_addr >= 6'h3e ? $random : idxs[idxs_T_2008_addr];
  `endif
  assign idxs_T_2011_addr = {{2'd0}, 4'hd};
  assign idxs_T_2011_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2011_data = idxs[idxs_T_2011_addr];
  `else
  assign idxs_T_2011_data = idxs_T_2011_addr >= 6'h3e ? $random : idxs[idxs_T_2011_addr];
  `endif
  assign idxs_T_2014_addr = {{2'd0}, 4'he};
  assign idxs_T_2014_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2014_data = idxs[idxs_T_2014_addr];
  `else
  assign idxs_T_2014_data = idxs_T_2014_addr >= 6'h3e ? $random : idxs[idxs_T_2014_addr];
  `endif
  assign idxs_T_2017_addr = {{2'd0}, 4'hf};
  assign idxs_T_2017_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2017_data = idxs[idxs_T_2017_addr];
  `else
  assign idxs_T_2017_data = idxs_T_2017_addr >= 6'h3e ? $random : idxs[idxs_T_2017_addr];
  `endif
  assign idxs_T_2020_addr = {{1'd0}, 5'h10};
  assign idxs_T_2020_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2020_data = idxs[idxs_T_2020_addr];
  `else
  assign idxs_T_2020_data = idxs_T_2020_addr >= 6'h3e ? $random : idxs[idxs_T_2020_addr];
  `endif
  assign idxs_T_2023_addr = {{1'd0}, 5'h11};
  assign idxs_T_2023_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2023_data = idxs[idxs_T_2023_addr];
  `else
  assign idxs_T_2023_data = idxs_T_2023_addr >= 6'h3e ? $random : idxs[idxs_T_2023_addr];
  `endif
  assign idxs_T_2026_addr = {{1'd0}, 5'h12};
  assign idxs_T_2026_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2026_data = idxs[idxs_T_2026_addr];
  `else
  assign idxs_T_2026_data = idxs_T_2026_addr >= 6'h3e ? $random : idxs[idxs_T_2026_addr];
  `endif
  assign idxs_T_2029_addr = {{1'd0}, 5'h13};
  assign idxs_T_2029_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2029_data = idxs[idxs_T_2029_addr];
  `else
  assign idxs_T_2029_data = idxs_T_2029_addr >= 6'h3e ? $random : idxs[idxs_T_2029_addr];
  `endif
  assign idxs_T_2032_addr = {{1'd0}, 5'h14};
  assign idxs_T_2032_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2032_data = idxs[idxs_T_2032_addr];
  `else
  assign idxs_T_2032_data = idxs_T_2032_addr >= 6'h3e ? $random : idxs[idxs_T_2032_addr];
  `endif
  assign idxs_T_2035_addr = {{1'd0}, 5'h15};
  assign idxs_T_2035_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2035_data = idxs[idxs_T_2035_addr];
  `else
  assign idxs_T_2035_data = idxs_T_2035_addr >= 6'h3e ? $random : idxs[idxs_T_2035_addr];
  `endif
  assign idxs_T_2038_addr = {{1'd0}, 5'h16};
  assign idxs_T_2038_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2038_data = idxs[idxs_T_2038_addr];
  `else
  assign idxs_T_2038_data = idxs_T_2038_addr >= 6'h3e ? $random : idxs[idxs_T_2038_addr];
  `endif
  assign idxs_T_2041_addr = {{1'd0}, 5'h17};
  assign idxs_T_2041_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2041_data = idxs[idxs_T_2041_addr];
  `else
  assign idxs_T_2041_data = idxs_T_2041_addr >= 6'h3e ? $random : idxs[idxs_T_2041_addr];
  `endif
  assign idxs_T_2044_addr = {{1'd0}, 5'h18};
  assign idxs_T_2044_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2044_data = idxs[idxs_T_2044_addr];
  `else
  assign idxs_T_2044_data = idxs_T_2044_addr >= 6'h3e ? $random : idxs[idxs_T_2044_addr];
  `endif
  assign idxs_T_2047_addr = {{1'd0}, 5'h19};
  assign idxs_T_2047_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2047_data = idxs[idxs_T_2047_addr];
  `else
  assign idxs_T_2047_data = idxs_T_2047_addr >= 6'h3e ? $random : idxs[idxs_T_2047_addr];
  `endif
  assign idxs_T_2050_addr = {{1'd0}, 5'h1a};
  assign idxs_T_2050_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2050_data = idxs[idxs_T_2050_addr];
  `else
  assign idxs_T_2050_data = idxs_T_2050_addr >= 6'h3e ? $random : idxs[idxs_T_2050_addr];
  `endif
  assign idxs_T_2053_addr = {{1'd0}, 5'h1b};
  assign idxs_T_2053_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2053_data = idxs[idxs_T_2053_addr];
  `else
  assign idxs_T_2053_data = idxs_T_2053_addr >= 6'h3e ? $random : idxs[idxs_T_2053_addr];
  `endif
  assign idxs_T_2056_addr = {{1'd0}, 5'h1c};
  assign idxs_T_2056_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2056_data = idxs[idxs_T_2056_addr];
  `else
  assign idxs_T_2056_data = idxs_T_2056_addr >= 6'h3e ? $random : idxs[idxs_T_2056_addr];
  `endif
  assign idxs_T_2059_addr = {{1'd0}, 5'h1d};
  assign idxs_T_2059_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2059_data = idxs[idxs_T_2059_addr];
  `else
  assign idxs_T_2059_data = idxs_T_2059_addr >= 6'h3e ? $random : idxs[idxs_T_2059_addr];
  `endif
  assign idxs_T_2062_addr = {{1'd0}, 5'h1e};
  assign idxs_T_2062_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2062_data = idxs[idxs_T_2062_addr];
  `else
  assign idxs_T_2062_data = idxs_T_2062_addr >= 6'h3e ? $random : idxs[idxs_T_2062_addr];
  `endif
  assign idxs_T_2065_addr = {{1'd0}, 5'h1f};
  assign idxs_T_2065_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2065_data = idxs[idxs_T_2065_addr];
  `else
  assign idxs_T_2065_data = idxs_T_2065_addr >= 6'h3e ? $random : idxs[idxs_T_2065_addr];
  `endif
  assign idxs_T_2068_addr = 6'h20;
  assign idxs_T_2068_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2068_data = idxs[idxs_T_2068_addr];
  `else
  assign idxs_T_2068_data = idxs_T_2068_addr >= 6'h3e ? $random : idxs[idxs_T_2068_addr];
  `endif
  assign idxs_T_2071_addr = 6'h21;
  assign idxs_T_2071_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2071_data = idxs[idxs_T_2071_addr];
  `else
  assign idxs_T_2071_data = idxs_T_2071_addr >= 6'h3e ? $random : idxs[idxs_T_2071_addr];
  `endif
  assign idxs_T_2074_addr = 6'h22;
  assign idxs_T_2074_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2074_data = idxs[idxs_T_2074_addr];
  `else
  assign idxs_T_2074_data = idxs_T_2074_addr >= 6'h3e ? $random : idxs[idxs_T_2074_addr];
  `endif
  assign idxs_T_2077_addr = 6'h23;
  assign idxs_T_2077_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2077_data = idxs[idxs_T_2077_addr];
  `else
  assign idxs_T_2077_data = idxs_T_2077_addr >= 6'h3e ? $random : idxs[idxs_T_2077_addr];
  `endif
  assign idxs_T_2080_addr = 6'h24;
  assign idxs_T_2080_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2080_data = idxs[idxs_T_2080_addr];
  `else
  assign idxs_T_2080_data = idxs_T_2080_addr >= 6'h3e ? $random : idxs[idxs_T_2080_addr];
  `endif
  assign idxs_T_2083_addr = 6'h25;
  assign idxs_T_2083_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2083_data = idxs[idxs_T_2083_addr];
  `else
  assign idxs_T_2083_data = idxs_T_2083_addr >= 6'h3e ? $random : idxs[idxs_T_2083_addr];
  `endif
  assign idxs_T_2086_addr = 6'h26;
  assign idxs_T_2086_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2086_data = idxs[idxs_T_2086_addr];
  `else
  assign idxs_T_2086_data = idxs_T_2086_addr >= 6'h3e ? $random : idxs[idxs_T_2086_addr];
  `endif
  assign idxs_T_2089_addr = 6'h27;
  assign idxs_T_2089_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2089_data = idxs[idxs_T_2089_addr];
  `else
  assign idxs_T_2089_data = idxs_T_2089_addr >= 6'h3e ? $random : idxs[idxs_T_2089_addr];
  `endif
  assign idxs_T_2092_addr = 6'h28;
  assign idxs_T_2092_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2092_data = idxs[idxs_T_2092_addr];
  `else
  assign idxs_T_2092_data = idxs_T_2092_addr >= 6'h3e ? $random : idxs[idxs_T_2092_addr];
  `endif
  assign idxs_T_2095_addr = 6'h29;
  assign idxs_T_2095_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2095_data = idxs[idxs_T_2095_addr];
  `else
  assign idxs_T_2095_data = idxs_T_2095_addr >= 6'h3e ? $random : idxs[idxs_T_2095_addr];
  `endif
  assign idxs_T_2098_addr = 6'h2a;
  assign idxs_T_2098_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2098_data = idxs[idxs_T_2098_addr];
  `else
  assign idxs_T_2098_data = idxs_T_2098_addr >= 6'h3e ? $random : idxs[idxs_T_2098_addr];
  `endif
  assign idxs_T_2101_addr = 6'h2b;
  assign idxs_T_2101_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2101_data = idxs[idxs_T_2101_addr];
  `else
  assign idxs_T_2101_data = idxs_T_2101_addr >= 6'h3e ? $random : idxs[idxs_T_2101_addr];
  `endif
  assign idxs_T_2104_addr = 6'h2c;
  assign idxs_T_2104_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2104_data = idxs[idxs_T_2104_addr];
  `else
  assign idxs_T_2104_data = idxs_T_2104_addr >= 6'h3e ? $random : idxs[idxs_T_2104_addr];
  `endif
  assign idxs_T_2107_addr = 6'h2d;
  assign idxs_T_2107_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2107_data = idxs[idxs_T_2107_addr];
  `else
  assign idxs_T_2107_data = idxs_T_2107_addr >= 6'h3e ? $random : idxs[idxs_T_2107_addr];
  `endif
  assign idxs_T_2110_addr = 6'h2e;
  assign idxs_T_2110_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2110_data = idxs[idxs_T_2110_addr];
  `else
  assign idxs_T_2110_data = idxs_T_2110_addr >= 6'h3e ? $random : idxs[idxs_T_2110_addr];
  `endif
  assign idxs_T_2113_addr = 6'h2f;
  assign idxs_T_2113_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2113_data = idxs[idxs_T_2113_addr];
  `else
  assign idxs_T_2113_data = idxs_T_2113_addr >= 6'h3e ? $random : idxs[idxs_T_2113_addr];
  `endif
  assign idxs_T_2116_addr = 6'h30;
  assign idxs_T_2116_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2116_data = idxs[idxs_T_2116_addr];
  `else
  assign idxs_T_2116_data = idxs_T_2116_addr >= 6'h3e ? $random : idxs[idxs_T_2116_addr];
  `endif
  assign idxs_T_2119_addr = 6'h31;
  assign idxs_T_2119_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2119_data = idxs[idxs_T_2119_addr];
  `else
  assign idxs_T_2119_data = idxs_T_2119_addr >= 6'h3e ? $random : idxs[idxs_T_2119_addr];
  `endif
  assign idxs_T_2122_addr = 6'h32;
  assign idxs_T_2122_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2122_data = idxs[idxs_T_2122_addr];
  `else
  assign idxs_T_2122_data = idxs_T_2122_addr >= 6'h3e ? $random : idxs[idxs_T_2122_addr];
  `endif
  assign idxs_T_2125_addr = 6'h33;
  assign idxs_T_2125_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2125_data = idxs[idxs_T_2125_addr];
  `else
  assign idxs_T_2125_data = idxs_T_2125_addr >= 6'h3e ? $random : idxs[idxs_T_2125_addr];
  `endif
  assign idxs_T_2128_addr = 6'h34;
  assign idxs_T_2128_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2128_data = idxs[idxs_T_2128_addr];
  `else
  assign idxs_T_2128_data = idxs_T_2128_addr >= 6'h3e ? $random : idxs[idxs_T_2128_addr];
  `endif
  assign idxs_T_2131_addr = 6'h35;
  assign idxs_T_2131_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2131_data = idxs[idxs_T_2131_addr];
  `else
  assign idxs_T_2131_data = idxs_T_2131_addr >= 6'h3e ? $random : idxs[idxs_T_2131_addr];
  `endif
  assign idxs_T_2134_addr = 6'h36;
  assign idxs_T_2134_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2134_data = idxs[idxs_T_2134_addr];
  `else
  assign idxs_T_2134_data = idxs_T_2134_addr >= 6'h3e ? $random : idxs[idxs_T_2134_addr];
  `endif
  assign idxs_T_2137_addr = 6'h37;
  assign idxs_T_2137_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2137_data = idxs[idxs_T_2137_addr];
  `else
  assign idxs_T_2137_data = idxs_T_2137_addr >= 6'h3e ? $random : idxs[idxs_T_2137_addr];
  `endif
  assign idxs_T_2140_addr = 6'h38;
  assign idxs_T_2140_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2140_data = idxs[idxs_T_2140_addr];
  `else
  assign idxs_T_2140_data = idxs_T_2140_addr >= 6'h3e ? $random : idxs[idxs_T_2140_addr];
  `endif
  assign idxs_T_2143_addr = 6'h39;
  assign idxs_T_2143_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2143_data = idxs[idxs_T_2143_addr];
  `else
  assign idxs_T_2143_data = idxs_T_2143_addr >= 6'h3e ? $random : idxs[idxs_T_2143_addr];
  `endif
  assign idxs_T_2146_addr = 6'h3a;
  assign idxs_T_2146_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2146_data = idxs[idxs_T_2146_addr];
  `else
  assign idxs_T_2146_data = idxs_T_2146_addr >= 6'h3e ? $random : idxs[idxs_T_2146_addr];
  `endif
  assign idxs_T_2149_addr = 6'h3b;
  assign idxs_T_2149_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2149_data = idxs[idxs_T_2149_addr];
  `else
  assign idxs_T_2149_data = idxs_T_2149_addr >= 6'h3e ? $random : idxs[idxs_T_2149_addr];
  `endif
  assign idxs_T_2152_addr = 6'h3c;
  assign idxs_T_2152_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2152_data = idxs[idxs_T_2152_addr];
  `else
  assign idxs_T_2152_data = idxs_T_2152_addr >= 6'h3e ? $random : idxs[idxs_T_2152_addr];
  `endif
  assign idxs_T_2155_addr = 6'h3d;
  assign idxs_T_2155_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxs_T_2155_data = idxs[idxs_T_2155_addr];
  `else
  assign idxs_T_2155_data = idxs_T_2155_addr >= 6'h3e ? $random : idxs[idxs_T_2155_addr];
  `endif
  assign idxs_T_2872_data = r_btb_update_bits_pc[11:0];
  assign idxs_T_2872_addr = T_2550;
  assign idxs_T_2872_mask = r_btb_update_valid;
  assign idxs_T_2872_en = r_btb_update_valid;
  assign idxPages_T_578_addr = {{5'd0}, 1'h0};
  assign idxPages_T_578_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_578_data = idxPages[idxPages_T_578_addr];
  `else
  assign idxPages_T_578_data = idxPages_T_578_addr >= 6'h3e ? $random : idxPages[idxPages_T_578_addr];
  `endif
  assign idxPages_T_583_addr = {{5'd0}, 1'h1};
  assign idxPages_T_583_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_583_data = idxPages[idxPages_T_583_addr];
  `else
  assign idxPages_T_583_data = idxPages_T_583_addr >= 6'h3e ? $random : idxPages[idxPages_T_583_addr];
  `endif
  assign idxPages_T_588_addr = {{4'd0}, 2'h2};
  assign idxPages_T_588_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_588_data = idxPages[idxPages_T_588_addr];
  `else
  assign idxPages_T_588_data = idxPages_T_588_addr >= 6'h3e ? $random : idxPages[idxPages_T_588_addr];
  `endif
  assign idxPages_T_593_addr = {{4'd0}, 2'h3};
  assign idxPages_T_593_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_593_data = idxPages[idxPages_T_593_addr];
  `else
  assign idxPages_T_593_data = idxPages_T_593_addr >= 6'h3e ? $random : idxPages[idxPages_T_593_addr];
  `endif
  assign idxPages_T_598_addr = {{3'd0}, 3'h4};
  assign idxPages_T_598_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_598_data = idxPages[idxPages_T_598_addr];
  `else
  assign idxPages_T_598_data = idxPages_T_598_addr >= 6'h3e ? $random : idxPages[idxPages_T_598_addr];
  `endif
  assign idxPages_T_603_addr = {{3'd0}, 3'h5};
  assign idxPages_T_603_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_603_data = idxPages[idxPages_T_603_addr];
  `else
  assign idxPages_T_603_data = idxPages_T_603_addr >= 6'h3e ? $random : idxPages[idxPages_T_603_addr];
  `endif
  assign idxPages_T_608_addr = {{3'd0}, 3'h6};
  assign idxPages_T_608_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_608_data = idxPages[idxPages_T_608_addr];
  `else
  assign idxPages_T_608_data = idxPages_T_608_addr >= 6'h3e ? $random : idxPages[idxPages_T_608_addr];
  `endif
  assign idxPages_T_613_addr = {{3'd0}, 3'h7};
  assign idxPages_T_613_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_613_data = idxPages[idxPages_T_613_addr];
  `else
  assign idxPages_T_613_data = idxPages_T_613_addr >= 6'h3e ? $random : idxPages[idxPages_T_613_addr];
  `endif
  assign idxPages_T_618_addr = {{2'd0}, 4'h8};
  assign idxPages_T_618_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_618_data = idxPages[idxPages_T_618_addr];
  `else
  assign idxPages_T_618_data = idxPages_T_618_addr >= 6'h3e ? $random : idxPages[idxPages_T_618_addr];
  `endif
  assign idxPages_T_623_addr = {{2'd0}, 4'h9};
  assign idxPages_T_623_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_623_data = idxPages[idxPages_T_623_addr];
  `else
  assign idxPages_T_623_data = idxPages_T_623_addr >= 6'h3e ? $random : idxPages[idxPages_T_623_addr];
  `endif
  assign idxPages_T_628_addr = {{2'd0}, 4'ha};
  assign idxPages_T_628_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_628_data = idxPages[idxPages_T_628_addr];
  `else
  assign idxPages_T_628_data = idxPages_T_628_addr >= 6'h3e ? $random : idxPages[idxPages_T_628_addr];
  `endif
  assign idxPages_T_633_addr = {{2'd0}, 4'hb};
  assign idxPages_T_633_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_633_data = idxPages[idxPages_T_633_addr];
  `else
  assign idxPages_T_633_data = idxPages_T_633_addr >= 6'h3e ? $random : idxPages[idxPages_T_633_addr];
  `endif
  assign idxPages_T_638_addr = {{2'd0}, 4'hc};
  assign idxPages_T_638_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_638_data = idxPages[idxPages_T_638_addr];
  `else
  assign idxPages_T_638_data = idxPages_T_638_addr >= 6'h3e ? $random : idxPages[idxPages_T_638_addr];
  `endif
  assign idxPages_T_643_addr = {{2'd0}, 4'hd};
  assign idxPages_T_643_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_643_data = idxPages[idxPages_T_643_addr];
  `else
  assign idxPages_T_643_data = idxPages_T_643_addr >= 6'h3e ? $random : idxPages[idxPages_T_643_addr];
  `endif
  assign idxPages_T_648_addr = {{2'd0}, 4'he};
  assign idxPages_T_648_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_648_data = idxPages[idxPages_T_648_addr];
  `else
  assign idxPages_T_648_data = idxPages_T_648_addr >= 6'h3e ? $random : idxPages[idxPages_T_648_addr];
  `endif
  assign idxPages_T_653_addr = {{2'd0}, 4'hf};
  assign idxPages_T_653_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_653_data = idxPages[idxPages_T_653_addr];
  `else
  assign idxPages_T_653_data = idxPages_T_653_addr >= 6'h3e ? $random : idxPages[idxPages_T_653_addr];
  `endif
  assign idxPages_T_658_addr = {{1'd0}, 5'h10};
  assign idxPages_T_658_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_658_data = idxPages[idxPages_T_658_addr];
  `else
  assign idxPages_T_658_data = idxPages_T_658_addr >= 6'h3e ? $random : idxPages[idxPages_T_658_addr];
  `endif
  assign idxPages_T_663_addr = {{1'd0}, 5'h11};
  assign idxPages_T_663_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_663_data = idxPages[idxPages_T_663_addr];
  `else
  assign idxPages_T_663_data = idxPages_T_663_addr >= 6'h3e ? $random : idxPages[idxPages_T_663_addr];
  `endif
  assign idxPages_T_668_addr = {{1'd0}, 5'h12};
  assign idxPages_T_668_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_668_data = idxPages[idxPages_T_668_addr];
  `else
  assign idxPages_T_668_data = idxPages_T_668_addr >= 6'h3e ? $random : idxPages[idxPages_T_668_addr];
  `endif
  assign idxPages_T_673_addr = {{1'd0}, 5'h13};
  assign idxPages_T_673_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_673_data = idxPages[idxPages_T_673_addr];
  `else
  assign idxPages_T_673_data = idxPages_T_673_addr >= 6'h3e ? $random : idxPages[idxPages_T_673_addr];
  `endif
  assign idxPages_T_678_addr = {{1'd0}, 5'h14};
  assign idxPages_T_678_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_678_data = idxPages[idxPages_T_678_addr];
  `else
  assign idxPages_T_678_data = idxPages_T_678_addr >= 6'h3e ? $random : idxPages[idxPages_T_678_addr];
  `endif
  assign idxPages_T_683_addr = {{1'd0}, 5'h15};
  assign idxPages_T_683_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_683_data = idxPages[idxPages_T_683_addr];
  `else
  assign idxPages_T_683_data = idxPages_T_683_addr >= 6'h3e ? $random : idxPages[idxPages_T_683_addr];
  `endif
  assign idxPages_T_688_addr = {{1'd0}, 5'h16};
  assign idxPages_T_688_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_688_data = idxPages[idxPages_T_688_addr];
  `else
  assign idxPages_T_688_data = idxPages_T_688_addr >= 6'h3e ? $random : idxPages[idxPages_T_688_addr];
  `endif
  assign idxPages_T_693_addr = {{1'd0}, 5'h17};
  assign idxPages_T_693_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_693_data = idxPages[idxPages_T_693_addr];
  `else
  assign idxPages_T_693_data = idxPages_T_693_addr >= 6'h3e ? $random : idxPages[idxPages_T_693_addr];
  `endif
  assign idxPages_T_698_addr = {{1'd0}, 5'h18};
  assign idxPages_T_698_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_698_data = idxPages[idxPages_T_698_addr];
  `else
  assign idxPages_T_698_data = idxPages_T_698_addr >= 6'h3e ? $random : idxPages[idxPages_T_698_addr];
  `endif
  assign idxPages_T_703_addr = {{1'd0}, 5'h19};
  assign idxPages_T_703_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_703_data = idxPages[idxPages_T_703_addr];
  `else
  assign idxPages_T_703_data = idxPages_T_703_addr >= 6'h3e ? $random : idxPages[idxPages_T_703_addr];
  `endif
  assign idxPages_T_708_addr = {{1'd0}, 5'h1a};
  assign idxPages_T_708_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_708_data = idxPages[idxPages_T_708_addr];
  `else
  assign idxPages_T_708_data = idxPages_T_708_addr >= 6'h3e ? $random : idxPages[idxPages_T_708_addr];
  `endif
  assign idxPages_T_713_addr = {{1'd0}, 5'h1b};
  assign idxPages_T_713_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_713_data = idxPages[idxPages_T_713_addr];
  `else
  assign idxPages_T_713_data = idxPages_T_713_addr >= 6'h3e ? $random : idxPages[idxPages_T_713_addr];
  `endif
  assign idxPages_T_718_addr = {{1'd0}, 5'h1c};
  assign idxPages_T_718_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_718_data = idxPages[idxPages_T_718_addr];
  `else
  assign idxPages_T_718_data = idxPages_T_718_addr >= 6'h3e ? $random : idxPages[idxPages_T_718_addr];
  `endif
  assign idxPages_T_723_addr = {{1'd0}, 5'h1d};
  assign idxPages_T_723_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_723_data = idxPages[idxPages_T_723_addr];
  `else
  assign idxPages_T_723_data = idxPages_T_723_addr >= 6'h3e ? $random : idxPages[idxPages_T_723_addr];
  `endif
  assign idxPages_T_728_addr = {{1'd0}, 5'h1e};
  assign idxPages_T_728_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_728_data = idxPages[idxPages_T_728_addr];
  `else
  assign idxPages_T_728_data = idxPages_T_728_addr >= 6'h3e ? $random : idxPages[idxPages_T_728_addr];
  `endif
  assign idxPages_T_733_addr = {{1'd0}, 5'h1f};
  assign idxPages_T_733_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_733_data = idxPages[idxPages_T_733_addr];
  `else
  assign idxPages_T_733_data = idxPages_T_733_addr >= 6'h3e ? $random : idxPages[idxPages_T_733_addr];
  `endif
  assign idxPages_T_738_addr = 6'h20;
  assign idxPages_T_738_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_738_data = idxPages[idxPages_T_738_addr];
  `else
  assign idxPages_T_738_data = idxPages_T_738_addr >= 6'h3e ? $random : idxPages[idxPages_T_738_addr];
  `endif
  assign idxPages_T_743_addr = 6'h21;
  assign idxPages_T_743_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_743_data = idxPages[idxPages_T_743_addr];
  `else
  assign idxPages_T_743_data = idxPages_T_743_addr >= 6'h3e ? $random : idxPages[idxPages_T_743_addr];
  `endif
  assign idxPages_T_748_addr = 6'h22;
  assign idxPages_T_748_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_748_data = idxPages[idxPages_T_748_addr];
  `else
  assign idxPages_T_748_data = idxPages_T_748_addr >= 6'h3e ? $random : idxPages[idxPages_T_748_addr];
  `endif
  assign idxPages_T_753_addr = 6'h23;
  assign idxPages_T_753_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_753_data = idxPages[idxPages_T_753_addr];
  `else
  assign idxPages_T_753_data = idxPages_T_753_addr >= 6'h3e ? $random : idxPages[idxPages_T_753_addr];
  `endif
  assign idxPages_T_758_addr = 6'h24;
  assign idxPages_T_758_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_758_data = idxPages[idxPages_T_758_addr];
  `else
  assign idxPages_T_758_data = idxPages_T_758_addr >= 6'h3e ? $random : idxPages[idxPages_T_758_addr];
  `endif
  assign idxPages_T_763_addr = 6'h25;
  assign idxPages_T_763_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_763_data = idxPages[idxPages_T_763_addr];
  `else
  assign idxPages_T_763_data = idxPages_T_763_addr >= 6'h3e ? $random : idxPages[idxPages_T_763_addr];
  `endif
  assign idxPages_T_768_addr = 6'h26;
  assign idxPages_T_768_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_768_data = idxPages[idxPages_T_768_addr];
  `else
  assign idxPages_T_768_data = idxPages_T_768_addr >= 6'h3e ? $random : idxPages[idxPages_T_768_addr];
  `endif
  assign idxPages_T_773_addr = 6'h27;
  assign idxPages_T_773_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_773_data = idxPages[idxPages_T_773_addr];
  `else
  assign idxPages_T_773_data = idxPages_T_773_addr >= 6'h3e ? $random : idxPages[idxPages_T_773_addr];
  `endif
  assign idxPages_T_778_addr = 6'h28;
  assign idxPages_T_778_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_778_data = idxPages[idxPages_T_778_addr];
  `else
  assign idxPages_T_778_data = idxPages_T_778_addr >= 6'h3e ? $random : idxPages[idxPages_T_778_addr];
  `endif
  assign idxPages_T_783_addr = 6'h29;
  assign idxPages_T_783_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_783_data = idxPages[idxPages_T_783_addr];
  `else
  assign idxPages_T_783_data = idxPages_T_783_addr >= 6'h3e ? $random : idxPages[idxPages_T_783_addr];
  `endif
  assign idxPages_T_788_addr = 6'h2a;
  assign idxPages_T_788_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_788_data = idxPages[idxPages_T_788_addr];
  `else
  assign idxPages_T_788_data = idxPages_T_788_addr >= 6'h3e ? $random : idxPages[idxPages_T_788_addr];
  `endif
  assign idxPages_T_793_addr = 6'h2b;
  assign idxPages_T_793_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_793_data = idxPages[idxPages_T_793_addr];
  `else
  assign idxPages_T_793_data = idxPages_T_793_addr >= 6'h3e ? $random : idxPages[idxPages_T_793_addr];
  `endif
  assign idxPages_T_798_addr = 6'h2c;
  assign idxPages_T_798_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_798_data = idxPages[idxPages_T_798_addr];
  `else
  assign idxPages_T_798_data = idxPages_T_798_addr >= 6'h3e ? $random : idxPages[idxPages_T_798_addr];
  `endif
  assign idxPages_T_803_addr = 6'h2d;
  assign idxPages_T_803_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_803_data = idxPages[idxPages_T_803_addr];
  `else
  assign idxPages_T_803_data = idxPages_T_803_addr >= 6'h3e ? $random : idxPages[idxPages_T_803_addr];
  `endif
  assign idxPages_T_808_addr = 6'h2e;
  assign idxPages_T_808_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_808_data = idxPages[idxPages_T_808_addr];
  `else
  assign idxPages_T_808_data = idxPages_T_808_addr >= 6'h3e ? $random : idxPages[idxPages_T_808_addr];
  `endif
  assign idxPages_T_813_addr = 6'h2f;
  assign idxPages_T_813_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_813_data = idxPages[idxPages_T_813_addr];
  `else
  assign idxPages_T_813_data = idxPages_T_813_addr >= 6'h3e ? $random : idxPages[idxPages_T_813_addr];
  `endif
  assign idxPages_T_818_addr = 6'h30;
  assign idxPages_T_818_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_818_data = idxPages[idxPages_T_818_addr];
  `else
  assign idxPages_T_818_data = idxPages_T_818_addr >= 6'h3e ? $random : idxPages[idxPages_T_818_addr];
  `endif
  assign idxPages_T_823_addr = 6'h31;
  assign idxPages_T_823_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_823_data = idxPages[idxPages_T_823_addr];
  `else
  assign idxPages_T_823_data = idxPages_T_823_addr >= 6'h3e ? $random : idxPages[idxPages_T_823_addr];
  `endif
  assign idxPages_T_828_addr = 6'h32;
  assign idxPages_T_828_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_828_data = idxPages[idxPages_T_828_addr];
  `else
  assign idxPages_T_828_data = idxPages_T_828_addr >= 6'h3e ? $random : idxPages[idxPages_T_828_addr];
  `endif
  assign idxPages_T_833_addr = 6'h33;
  assign idxPages_T_833_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_833_data = idxPages[idxPages_T_833_addr];
  `else
  assign idxPages_T_833_data = idxPages_T_833_addr >= 6'h3e ? $random : idxPages[idxPages_T_833_addr];
  `endif
  assign idxPages_T_838_addr = 6'h34;
  assign idxPages_T_838_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_838_data = idxPages[idxPages_T_838_addr];
  `else
  assign idxPages_T_838_data = idxPages_T_838_addr >= 6'h3e ? $random : idxPages[idxPages_T_838_addr];
  `endif
  assign idxPages_T_843_addr = 6'h35;
  assign idxPages_T_843_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_843_data = idxPages[idxPages_T_843_addr];
  `else
  assign idxPages_T_843_data = idxPages_T_843_addr >= 6'h3e ? $random : idxPages[idxPages_T_843_addr];
  `endif
  assign idxPages_T_848_addr = 6'h36;
  assign idxPages_T_848_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_848_data = idxPages[idxPages_T_848_addr];
  `else
  assign idxPages_T_848_data = idxPages_T_848_addr >= 6'h3e ? $random : idxPages[idxPages_T_848_addr];
  `endif
  assign idxPages_T_853_addr = 6'h37;
  assign idxPages_T_853_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_853_data = idxPages[idxPages_T_853_addr];
  `else
  assign idxPages_T_853_data = idxPages_T_853_addr >= 6'h3e ? $random : idxPages[idxPages_T_853_addr];
  `endif
  assign idxPages_T_858_addr = 6'h38;
  assign idxPages_T_858_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_858_data = idxPages[idxPages_T_858_addr];
  `else
  assign idxPages_T_858_data = idxPages_T_858_addr >= 6'h3e ? $random : idxPages[idxPages_T_858_addr];
  `endif
  assign idxPages_T_863_addr = 6'h39;
  assign idxPages_T_863_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_863_data = idxPages[idxPages_T_863_addr];
  `else
  assign idxPages_T_863_data = idxPages_T_863_addr >= 6'h3e ? $random : idxPages[idxPages_T_863_addr];
  `endif
  assign idxPages_T_868_addr = 6'h3a;
  assign idxPages_T_868_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_868_data = idxPages[idxPages_T_868_addr];
  `else
  assign idxPages_T_868_data = idxPages_T_868_addr >= 6'h3e ? $random : idxPages[idxPages_T_868_addr];
  `endif
  assign idxPages_T_873_addr = 6'h3b;
  assign idxPages_T_873_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_873_data = idxPages[idxPages_T_873_addr];
  `else
  assign idxPages_T_873_data = idxPages_T_873_addr >= 6'h3e ? $random : idxPages[idxPages_T_873_addr];
  `endif
  assign idxPages_T_878_addr = 6'h3c;
  assign idxPages_T_878_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_878_data = idxPages[idxPages_T_878_addr];
  `else
  assign idxPages_T_878_data = idxPages_T_878_addr >= 6'h3e ? $random : idxPages[idxPages_T_878_addr];
  `endif
  assign idxPages_T_883_addr = 6'h3d;
  assign idxPages_T_883_en = 1'h1;
  `ifdef SYNTHESIS
  assign idxPages_T_883_data = idxPages[idxPages_T_883_addr];
  `else
  assign idxPages_T_883_data = idxPages_T_883_addr >= 6'h3e ? $random : idxPages[idxPages_T_883_addr];
  `endif
  assign idxPages_T_2874_data = idxPageUpdate;
  assign idxPages_T_2874_addr = T_2550;
  assign idxPages_T_2874_mask = r_btb_update_valid;
  assign idxPages_T_2874_en = r_btb_update_valid;
  assign tgts_T_3270_addr = {{5'd0}, 1'h0};
  assign tgts_T_3270_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3270_data = tgts[tgts_T_3270_addr];
  `else
  assign tgts_T_3270_data = tgts_T_3270_addr >= 6'h3e ? $random : tgts[tgts_T_3270_addr];
  `endif
  assign tgts_T_3272_addr = {{5'd0}, 1'h1};
  assign tgts_T_3272_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3272_data = tgts[tgts_T_3272_addr];
  `else
  assign tgts_T_3272_data = tgts_T_3272_addr >= 6'h3e ? $random : tgts[tgts_T_3272_addr];
  `endif
  assign tgts_T_3274_addr = {{4'd0}, 2'h2};
  assign tgts_T_3274_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3274_data = tgts[tgts_T_3274_addr];
  `else
  assign tgts_T_3274_data = tgts_T_3274_addr >= 6'h3e ? $random : tgts[tgts_T_3274_addr];
  `endif
  assign tgts_T_3276_addr = {{4'd0}, 2'h3};
  assign tgts_T_3276_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3276_data = tgts[tgts_T_3276_addr];
  `else
  assign tgts_T_3276_data = tgts_T_3276_addr >= 6'h3e ? $random : tgts[tgts_T_3276_addr];
  `endif
  assign tgts_T_3278_addr = {{3'd0}, 3'h4};
  assign tgts_T_3278_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3278_data = tgts[tgts_T_3278_addr];
  `else
  assign tgts_T_3278_data = tgts_T_3278_addr >= 6'h3e ? $random : tgts[tgts_T_3278_addr];
  `endif
  assign tgts_T_3280_addr = {{3'd0}, 3'h5};
  assign tgts_T_3280_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3280_data = tgts[tgts_T_3280_addr];
  `else
  assign tgts_T_3280_data = tgts_T_3280_addr >= 6'h3e ? $random : tgts[tgts_T_3280_addr];
  `endif
  assign tgts_T_3282_addr = {{3'd0}, 3'h6};
  assign tgts_T_3282_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3282_data = tgts[tgts_T_3282_addr];
  `else
  assign tgts_T_3282_data = tgts_T_3282_addr >= 6'h3e ? $random : tgts[tgts_T_3282_addr];
  `endif
  assign tgts_T_3284_addr = {{3'd0}, 3'h7};
  assign tgts_T_3284_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3284_data = tgts[tgts_T_3284_addr];
  `else
  assign tgts_T_3284_data = tgts_T_3284_addr >= 6'h3e ? $random : tgts[tgts_T_3284_addr];
  `endif
  assign tgts_T_3286_addr = {{2'd0}, 4'h8};
  assign tgts_T_3286_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3286_data = tgts[tgts_T_3286_addr];
  `else
  assign tgts_T_3286_data = tgts_T_3286_addr >= 6'h3e ? $random : tgts[tgts_T_3286_addr];
  `endif
  assign tgts_T_3288_addr = {{2'd0}, 4'h9};
  assign tgts_T_3288_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3288_data = tgts[tgts_T_3288_addr];
  `else
  assign tgts_T_3288_data = tgts_T_3288_addr >= 6'h3e ? $random : tgts[tgts_T_3288_addr];
  `endif
  assign tgts_T_3290_addr = {{2'd0}, 4'ha};
  assign tgts_T_3290_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3290_data = tgts[tgts_T_3290_addr];
  `else
  assign tgts_T_3290_data = tgts_T_3290_addr >= 6'h3e ? $random : tgts[tgts_T_3290_addr];
  `endif
  assign tgts_T_3292_addr = {{2'd0}, 4'hb};
  assign tgts_T_3292_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3292_data = tgts[tgts_T_3292_addr];
  `else
  assign tgts_T_3292_data = tgts_T_3292_addr >= 6'h3e ? $random : tgts[tgts_T_3292_addr];
  `endif
  assign tgts_T_3294_addr = {{2'd0}, 4'hc};
  assign tgts_T_3294_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3294_data = tgts[tgts_T_3294_addr];
  `else
  assign tgts_T_3294_data = tgts_T_3294_addr >= 6'h3e ? $random : tgts[tgts_T_3294_addr];
  `endif
  assign tgts_T_3296_addr = {{2'd0}, 4'hd};
  assign tgts_T_3296_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3296_data = tgts[tgts_T_3296_addr];
  `else
  assign tgts_T_3296_data = tgts_T_3296_addr >= 6'h3e ? $random : tgts[tgts_T_3296_addr];
  `endif
  assign tgts_T_3298_addr = {{2'd0}, 4'he};
  assign tgts_T_3298_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3298_data = tgts[tgts_T_3298_addr];
  `else
  assign tgts_T_3298_data = tgts_T_3298_addr >= 6'h3e ? $random : tgts[tgts_T_3298_addr];
  `endif
  assign tgts_T_3300_addr = {{2'd0}, 4'hf};
  assign tgts_T_3300_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3300_data = tgts[tgts_T_3300_addr];
  `else
  assign tgts_T_3300_data = tgts_T_3300_addr >= 6'h3e ? $random : tgts[tgts_T_3300_addr];
  `endif
  assign tgts_T_3302_addr = {{1'd0}, 5'h10};
  assign tgts_T_3302_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3302_data = tgts[tgts_T_3302_addr];
  `else
  assign tgts_T_3302_data = tgts_T_3302_addr >= 6'h3e ? $random : tgts[tgts_T_3302_addr];
  `endif
  assign tgts_T_3304_addr = {{1'd0}, 5'h11};
  assign tgts_T_3304_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3304_data = tgts[tgts_T_3304_addr];
  `else
  assign tgts_T_3304_data = tgts_T_3304_addr >= 6'h3e ? $random : tgts[tgts_T_3304_addr];
  `endif
  assign tgts_T_3306_addr = {{1'd0}, 5'h12};
  assign tgts_T_3306_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3306_data = tgts[tgts_T_3306_addr];
  `else
  assign tgts_T_3306_data = tgts_T_3306_addr >= 6'h3e ? $random : tgts[tgts_T_3306_addr];
  `endif
  assign tgts_T_3308_addr = {{1'd0}, 5'h13};
  assign tgts_T_3308_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3308_data = tgts[tgts_T_3308_addr];
  `else
  assign tgts_T_3308_data = tgts_T_3308_addr >= 6'h3e ? $random : tgts[tgts_T_3308_addr];
  `endif
  assign tgts_T_3310_addr = {{1'd0}, 5'h14};
  assign tgts_T_3310_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3310_data = tgts[tgts_T_3310_addr];
  `else
  assign tgts_T_3310_data = tgts_T_3310_addr >= 6'h3e ? $random : tgts[tgts_T_3310_addr];
  `endif
  assign tgts_T_3312_addr = {{1'd0}, 5'h15};
  assign tgts_T_3312_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3312_data = tgts[tgts_T_3312_addr];
  `else
  assign tgts_T_3312_data = tgts_T_3312_addr >= 6'h3e ? $random : tgts[tgts_T_3312_addr];
  `endif
  assign tgts_T_3314_addr = {{1'd0}, 5'h16};
  assign tgts_T_3314_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3314_data = tgts[tgts_T_3314_addr];
  `else
  assign tgts_T_3314_data = tgts_T_3314_addr >= 6'h3e ? $random : tgts[tgts_T_3314_addr];
  `endif
  assign tgts_T_3316_addr = {{1'd0}, 5'h17};
  assign tgts_T_3316_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3316_data = tgts[tgts_T_3316_addr];
  `else
  assign tgts_T_3316_data = tgts_T_3316_addr >= 6'h3e ? $random : tgts[tgts_T_3316_addr];
  `endif
  assign tgts_T_3318_addr = {{1'd0}, 5'h18};
  assign tgts_T_3318_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3318_data = tgts[tgts_T_3318_addr];
  `else
  assign tgts_T_3318_data = tgts_T_3318_addr >= 6'h3e ? $random : tgts[tgts_T_3318_addr];
  `endif
  assign tgts_T_3320_addr = {{1'd0}, 5'h19};
  assign tgts_T_3320_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3320_data = tgts[tgts_T_3320_addr];
  `else
  assign tgts_T_3320_data = tgts_T_3320_addr >= 6'h3e ? $random : tgts[tgts_T_3320_addr];
  `endif
  assign tgts_T_3322_addr = {{1'd0}, 5'h1a};
  assign tgts_T_3322_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3322_data = tgts[tgts_T_3322_addr];
  `else
  assign tgts_T_3322_data = tgts_T_3322_addr >= 6'h3e ? $random : tgts[tgts_T_3322_addr];
  `endif
  assign tgts_T_3324_addr = {{1'd0}, 5'h1b};
  assign tgts_T_3324_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3324_data = tgts[tgts_T_3324_addr];
  `else
  assign tgts_T_3324_data = tgts_T_3324_addr >= 6'h3e ? $random : tgts[tgts_T_3324_addr];
  `endif
  assign tgts_T_3326_addr = {{1'd0}, 5'h1c};
  assign tgts_T_3326_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3326_data = tgts[tgts_T_3326_addr];
  `else
  assign tgts_T_3326_data = tgts_T_3326_addr >= 6'h3e ? $random : tgts[tgts_T_3326_addr];
  `endif
  assign tgts_T_3328_addr = {{1'd0}, 5'h1d};
  assign tgts_T_3328_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3328_data = tgts[tgts_T_3328_addr];
  `else
  assign tgts_T_3328_data = tgts_T_3328_addr >= 6'h3e ? $random : tgts[tgts_T_3328_addr];
  `endif
  assign tgts_T_3330_addr = {{1'd0}, 5'h1e};
  assign tgts_T_3330_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3330_data = tgts[tgts_T_3330_addr];
  `else
  assign tgts_T_3330_data = tgts_T_3330_addr >= 6'h3e ? $random : tgts[tgts_T_3330_addr];
  `endif
  assign tgts_T_3332_addr = {{1'd0}, 5'h1f};
  assign tgts_T_3332_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3332_data = tgts[tgts_T_3332_addr];
  `else
  assign tgts_T_3332_data = tgts_T_3332_addr >= 6'h3e ? $random : tgts[tgts_T_3332_addr];
  `endif
  assign tgts_T_3334_addr = 6'h20;
  assign tgts_T_3334_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3334_data = tgts[tgts_T_3334_addr];
  `else
  assign tgts_T_3334_data = tgts_T_3334_addr >= 6'h3e ? $random : tgts[tgts_T_3334_addr];
  `endif
  assign tgts_T_3336_addr = 6'h21;
  assign tgts_T_3336_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3336_data = tgts[tgts_T_3336_addr];
  `else
  assign tgts_T_3336_data = tgts_T_3336_addr >= 6'h3e ? $random : tgts[tgts_T_3336_addr];
  `endif
  assign tgts_T_3338_addr = 6'h22;
  assign tgts_T_3338_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3338_data = tgts[tgts_T_3338_addr];
  `else
  assign tgts_T_3338_data = tgts_T_3338_addr >= 6'h3e ? $random : tgts[tgts_T_3338_addr];
  `endif
  assign tgts_T_3340_addr = 6'h23;
  assign tgts_T_3340_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3340_data = tgts[tgts_T_3340_addr];
  `else
  assign tgts_T_3340_data = tgts_T_3340_addr >= 6'h3e ? $random : tgts[tgts_T_3340_addr];
  `endif
  assign tgts_T_3342_addr = 6'h24;
  assign tgts_T_3342_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3342_data = tgts[tgts_T_3342_addr];
  `else
  assign tgts_T_3342_data = tgts_T_3342_addr >= 6'h3e ? $random : tgts[tgts_T_3342_addr];
  `endif
  assign tgts_T_3344_addr = 6'h25;
  assign tgts_T_3344_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3344_data = tgts[tgts_T_3344_addr];
  `else
  assign tgts_T_3344_data = tgts_T_3344_addr >= 6'h3e ? $random : tgts[tgts_T_3344_addr];
  `endif
  assign tgts_T_3346_addr = 6'h26;
  assign tgts_T_3346_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3346_data = tgts[tgts_T_3346_addr];
  `else
  assign tgts_T_3346_data = tgts_T_3346_addr >= 6'h3e ? $random : tgts[tgts_T_3346_addr];
  `endif
  assign tgts_T_3348_addr = 6'h27;
  assign tgts_T_3348_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3348_data = tgts[tgts_T_3348_addr];
  `else
  assign tgts_T_3348_data = tgts_T_3348_addr >= 6'h3e ? $random : tgts[tgts_T_3348_addr];
  `endif
  assign tgts_T_3350_addr = 6'h28;
  assign tgts_T_3350_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3350_data = tgts[tgts_T_3350_addr];
  `else
  assign tgts_T_3350_data = tgts_T_3350_addr >= 6'h3e ? $random : tgts[tgts_T_3350_addr];
  `endif
  assign tgts_T_3352_addr = 6'h29;
  assign tgts_T_3352_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3352_data = tgts[tgts_T_3352_addr];
  `else
  assign tgts_T_3352_data = tgts_T_3352_addr >= 6'h3e ? $random : tgts[tgts_T_3352_addr];
  `endif
  assign tgts_T_3354_addr = 6'h2a;
  assign tgts_T_3354_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3354_data = tgts[tgts_T_3354_addr];
  `else
  assign tgts_T_3354_data = tgts_T_3354_addr >= 6'h3e ? $random : tgts[tgts_T_3354_addr];
  `endif
  assign tgts_T_3356_addr = 6'h2b;
  assign tgts_T_3356_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3356_data = tgts[tgts_T_3356_addr];
  `else
  assign tgts_T_3356_data = tgts_T_3356_addr >= 6'h3e ? $random : tgts[tgts_T_3356_addr];
  `endif
  assign tgts_T_3358_addr = 6'h2c;
  assign tgts_T_3358_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3358_data = tgts[tgts_T_3358_addr];
  `else
  assign tgts_T_3358_data = tgts_T_3358_addr >= 6'h3e ? $random : tgts[tgts_T_3358_addr];
  `endif
  assign tgts_T_3360_addr = 6'h2d;
  assign tgts_T_3360_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3360_data = tgts[tgts_T_3360_addr];
  `else
  assign tgts_T_3360_data = tgts_T_3360_addr >= 6'h3e ? $random : tgts[tgts_T_3360_addr];
  `endif
  assign tgts_T_3362_addr = 6'h2e;
  assign tgts_T_3362_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3362_data = tgts[tgts_T_3362_addr];
  `else
  assign tgts_T_3362_data = tgts_T_3362_addr >= 6'h3e ? $random : tgts[tgts_T_3362_addr];
  `endif
  assign tgts_T_3364_addr = 6'h2f;
  assign tgts_T_3364_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3364_data = tgts[tgts_T_3364_addr];
  `else
  assign tgts_T_3364_data = tgts_T_3364_addr >= 6'h3e ? $random : tgts[tgts_T_3364_addr];
  `endif
  assign tgts_T_3366_addr = 6'h30;
  assign tgts_T_3366_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3366_data = tgts[tgts_T_3366_addr];
  `else
  assign tgts_T_3366_data = tgts_T_3366_addr >= 6'h3e ? $random : tgts[tgts_T_3366_addr];
  `endif
  assign tgts_T_3368_addr = 6'h31;
  assign tgts_T_3368_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3368_data = tgts[tgts_T_3368_addr];
  `else
  assign tgts_T_3368_data = tgts_T_3368_addr >= 6'h3e ? $random : tgts[tgts_T_3368_addr];
  `endif
  assign tgts_T_3370_addr = 6'h32;
  assign tgts_T_3370_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3370_data = tgts[tgts_T_3370_addr];
  `else
  assign tgts_T_3370_data = tgts_T_3370_addr >= 6'h3e ? $random : tgts[tgts_T_3370_addr];
  `endif
  assign tgts_T_3372_addr = 6'h33;
  assign tgts_T_3372_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3372_data = tgts[tgts_T_3372_addr];
  `else
  assign tgts_T_3372_data = tgts_T_3372_addr >= 6'h3e ? $random : tgts[tgts_T_3372_addr];
  `endif
  assign tgts_T_3374_addr = 6'h34;
  assign tgts_T_3374_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3374_data = tgts[tgts_T_3374_addr];
  `else
  assign tgts_T_3374_data = tgts_T_3374_addr >= 6'h3e ? $random : tgts[tgts_T_3374_addr];
  `endif
  assign tgts_T_3376_addr = 6'h35;
  assign tgts_T_3376_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3376_data = tgts[tgts_T_3376_addr];
  `else
  assign tgts_T_3376_data = tgts_T_3376_addr >= 6'h3e ? $random : tgts[tgts_T_3376_addr];
  `endif
  assign tgts_T_3378_addr = 6'h36;
  assign tgts_T_3378_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3378_data = tgts[tgts_T_3378_addr];
  `else
  assign tgts_T_3378_data = tgts_T_3378_addr >= 6'h3e ? $random : tgts[tgts_T_3378_addr];
  `endif
  assign tgts_T_3380_addr = 6'h37;
  assign tgts_T_3380_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3380_data = tgts[tgts_T_3380_addr];
  `else
  assign tgts_T_3380_data = tgts_T_3380_addr >= 6'h3e ? $random : tgts[tgts_T_3380_addr];
  `endif
  assign tgts_T_3382_addr = 6'h38;
  assign tgts_T_3382_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3382_data = tgts[tgts_T_3382_addr];
  `else
  assign tgts_T_3382_data = tgts_T_3382_addr >= 6'h3e ? $random : tgts[tgts_T_3382_addr];
  `endif
  assign tgts_T_3384_addr = 6'h39;
  assign tgts_T_3384_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3384_data = tgts[tgts_T_3384_addr];
  `else
  assign tgts_T_3384_data = tgts_T_3384_addr >= 6'h3e ? $random : tgts[tgts_T_3384_addr];
  `endif
  assign tgts_T_3386_addr = 6'h3a;
  assign tgts_T_3386_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3386_data = tgts[tgts_T_3386_addr];
  `else
  assign tgts_T_3386_data = tgts_T_3386_addr >= 6'h3e ? $random : tgts[tgts_T_3386_addr];
  `endif
  assign tgts_T_3388_addr = 6'h3b;
  assign tgts_T_3388_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3388_data = tgts[tgts_T_3388_addr];
  `else
  assign tgts_T_3388_data = tgts_T_3388_addr >= 6'h3e ? $random : tgts[tgts_T_3388_addr];
  `endif
  assign tgts_T_3390_addr = 6'h3c;
  assign tgts_T_3390_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3390_data = tgts[tgts_T_3390_addr];
  `else
  assign tgts_T_3390_data = tgts_T_3390_addr >= 6'h3e ? $random : tgts[tgts_T_3390_addr];
  `endif
  assign tgts_T_3392_addr = 6'h3d;
  assign tgts_T_3392_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgts_T_3392_data = tgts[tgts_T_3392_addr];
  `else
  assign tgts_T_3392_data = tgts_T_3392_addr >= 6'h3e ? $random : tgts[tgts_T_3392_addr];
  `endif
  assign tgts_T_2873_data = io_req_bits_addr[11:0];
  assign tgts_T_2873_addr = T_2550;
  assign tgts_T_2873_mask = r_btb_update_valid;
  assign tgts_T_2873_en = r_btb_update_valid;
  assign tgtPages_T_888_addr = {{5'd0}, 1'h0};
  assign tgtPages_T_888_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_888_data = tgtPages[tgtPages_T_888_addr];
  `else
  assign tgtPages_T_888_data = tgtPages_T_888_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_888_addr];
  `endif
  assign tgtPages_T_893_addr = {{5'd0}, 1'h1};
  assign tgtPages_T_893_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_893_data = tgtPages[tgtPages_T_893_addr];
  `else
  assign tgtPages_T_893_data = tgtPages_T_893_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_893_addr];
  `endif
  assign tgtPages_T_898_addr = {{4'd0}, 2'h2};
  assign tgtPages_T_898_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_898_data = tgtPages[tgtPages_T_898_addr];
  `else
  assign tgtPages_T_898_data = tgtPages_T_898_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_898_addr];
  `endif
  assign tgtPages_T_903_addr = {{4'd0}, 2'h3};
  assign tgtPages_T_903_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_903_data = tgtPages[tgtPages_T_903_addr];
  `else
  assign tgtPages_T_903_data = tgtPages_T_903_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_903_addr];
  `endif
  assign tgtPages_T_908_addr = {{3'd0}, 3'h4};
  assign tgtPages_T_908_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_908_data = tgtPages[tgtPages_T_908_addr];
  `else
  assign tgtPages_T_908_data = tgtPages_T_908_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_908_addr];
  `endif
  assign tgtPages_T_913_addr = {{3'd0}, 3'h5};
  assign tgtPages_T_913_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_913_data = tgtPages[tgtPages_T_913_addr];
  `else
  assign tgtPages_T_913_data = tgtPages_T_913_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_913_addr];
  `endif
  assign tgtPages_T_918_addr = {{3'd0}, 3'h6};
  assign tgtPages_T_918_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_918_data = tgtPages[tgtPages_T_918_addr];
  `else
  assign tgtPages_T_918_data = tgtPages_T_918_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_918_addr];
  `endif
  assign tgtPages_T_923_addr = {{3'd0}, 3'h7};
  assign tgtPages_T_923_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_923_data = tgtPages[tgtPages_T_923_addr];
  `else
  assign tgtPages_T_923_data = tgtPages_T_923_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_923_addr];
  `endif
  assign tgtPages_T_928_addr = {{2'd0}, 4'h8};
  assign tgtPages_T_928_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_928_data = tgtPages[tgtPages_T_928_addr];
  `else
  assign tgtPages_T_928_data = tgtPages_T_928_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_928_addr];
  `endif
  assign tgtPages_T_933_addr = {{2'd0}, 4'h9};
  assign tgtPages_T_933_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_933_data = tgtPages[tgtPages_T_933_addr];
  `else
  assign tgtPages_T_933_data = tgtPages_T_933_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_933_addr];
  `endif
  assign tgtPages_T_938_addr = {{2'd0}, 4'ha};
  assign tgtPages_T_938_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_938_data = tgtPages[tgtPages_T_938_addr];
  `else
  assign tgtPages_T_938_data = tgtPages_T_938_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_938_addr];
  `endif
  assign tgtPages_T_943_addr = {{2'd0}, 4'hb};
  assign tgtPages_T_943_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_943_data = tgtPages[tgtPages_T_943_addr];
  `else
  assign tgtPages_T_943_data = tgtPages_T_943_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_943_addr];
  `endif
  assign tgtPages_T_948_addr = {{2'd0}, 4'hc};
  assign tgtPages_T_948_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_948_data = tgtPages[tgtPages_T_948_addr];
  `else
  assign tgtPages_T_948_data = tgtPages_T_948_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_948_addr];
  `endif
  assign tgtPages_T_953_addr = {{2'd0}, 4'hd};
  assign tgtPages_T_953_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_953_data = tgtPages[tgtPages_T_953_addr];
  `else
  assign tgtPages_T_953_data = tgtPages_T_953_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_953_addr];
  `endif
  assign tgtPages_T_958_addr = {{2'd0}, 4'he};
  assign tgtPages_T_958_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_958_data = tgtPages[tgtPages_T_958_addr];
  `else
  assign tgtPages_T_958_data = tgtPages_T_958_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_958_addr];
  `endif
  assign tgtPages_T_963_addr = {{2'd0}, 4'hf};
  assign tgtPages_T_963_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_963_data = tgtPages[tgtPages_T_963_addr];
  `else
  assign tgtPages_T_963_data = tgtPages_T_963_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_963_addr];
  `endif
  assign tgtPages_T_968_addr = {{1'd0}, 5'h10};
  assign tgtPages_T_968_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_968_data = tgtPages[tgtPages_T_968_addr];
  `else
  assign tgtPages_T_968_data = tgtPages_T_968_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_968_addr];
  `endif
  assign tgtPages_T_973_addr = {{1'd0}, 5'h11};
  assign tgtPages_T_973_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_973_data = tgtPages[tgtPages_T_973_addr];
  `else
  assign tgtPages_T_973_data = tgtPages_T_973_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_973_addr];
  `endif
  assign tgtPages_T_978_addr = {{1'd0}, 5'h12};
  assign tgtPages_T_978_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_978_data = tgtPages[tgtPages_T_978_addr];
  `else
  assign tgtPages_T_978_data = tgtPages_T_978_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_978_addr];
  `endif
  assign tgtPages_T_983_addr = {{1'd0}, 5'h13};
  assign tgtPages_T_983_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_983_data = tgtPages[tgtPages_T_983_addr];
  `else
  assign tgtPages_T_983_data = tgtPages_T_983_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_983_addr];
  `endif
  assign tgtPages_T_988_addr = {{1'd0}, 5'h14};
  assign tgtPages_T_988_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_988_data = tgtPages[tgtPages_T_988_addr];
  `else
  assign tgtPages_T_988_data = tgtPages_T_988_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_988_addr];
  `endif
  assign tgtPages_T_993_addr = {{1'd0}, 5'h15};
  assign tgtPages_T_993_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_993_data = tgtPages[tgtPages_T_993_addr];
  `else
  assign tgtPages_T_993_data = tgtPages_T_993_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_993_addr];
  `endif
  assign tgtPages_T_998_addr = {{1'd0}, 5'h16};
  assign tgtPages_T_998_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_998_data = tgtPages[tgtPages_T_998_addr];
  `else
  assign tgtPages_T_998_data = tgtPages_T_998_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_998_addr];
  `endif
  assign tgtPages_T_1003_addr = {{1'd0}, 5'h17};
  assign tgtPages_T_1003_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1003_data = tgtPages[tgtPages_T_1003_addr];
  `else
  assign tgtPages_T_1003_data = tgtPages_T_1003_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1003_addr];
  `endif
  assign tgtPages_T_1008_addr = {{1'd0}, 5'h18};
  assign tgtPages_T_1008_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1008_data = tgtPages[tgtPages_T_1008_addr];
  `else
  assign tgtPages_T_1008_data = tgtPages_T_1008_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1008_addr];
  `endif
  assign tgtPages_T_1013_addr = {{1'd0}, 5'h19};
  assign tgtPages_T_1013_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1013_data = tgtPages[tgtPages_T_1013_addr];
  `else
  assign tgtPages_T_1013_data = tgtPages_T_1013_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1013_addr];
  `endif
  assign tgtPages_T_1018_addr = {{1'd0}, 5'h1a};
  assign tgtPages_T_1018_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1018_data = tgtPages[tgtPages_T_1018_addr];
  `else
  assign tgtPages_T_1018_data = tgtPages_T_1018_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1018_addr];
  `endif
  assign tgtPages_T_1023_addr = {{1'd0}, 5'h1b};
  assign tgtPages_T_1023_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1023_data = tgtPages[tgtPages_T_1023_addr];
  `else
  assign tgtPages_T_1023_data = tgtPages_T_1023_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1023_addr];
  `endif
  assign tgtPages_T_1028_addr = {{1'd0}, 5'h1c};
  assign tgtPages_T_1028_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1028_data = tgtPages[tgtPages_T_1028_addr];
  `else
  assign tgtPages_T_1028_data = tgtPages_T_1028_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1028_addr];
  `endif
  assign tgtPages_T_1033_addr = {{1'd0}, 5'h1d};
  assign tgtPages_T_1033_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1033_data = tgtPages[tgtPages_T_1033_addr];
  `else
  assign tgtPages_T_1033_data = tgtPages_T_1033_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1033_addr];
  `endif
  assign tgtPages_T_1038_addr = {{1'd0}, 5'h1e};
  assign tgtPages_T_1038_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1038_data = tgtPages[tgtPages_T_1038_addr];
  `else
  assign tgtPages_T_1038_data = tgtPages_T_1038_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1038_addr];
  `endif
  assign tgtPages_T_1043_addr = {{1'd0}, 5'h1f};
  assign tgtPages_T_1043_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1043_data = tgtPages[tgtPages_T_1043_addr];
  `else
  assign tgtPages_T_1043_data = tgtPages_T_1043_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1043_addr];
  `endif
  assign tgtPages_T_1048_addr = 6'h20;
  assign tgtPages_T_1048_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1048_data = tgtPages[tgtPages_T_1048_addr];
  `else
  assign tgtPages_T_1048_data = tgtPages_T_1048_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1048_addr];
  `endif
  assign tgtPages_T_1053_addr = 6'h21;
  assign tgtPages_T_1053_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1053_data = tgtPages[tgtPages_T_1053_addr];
  `else
  assign tgtPages_T_1053_data = tgtPages_T_1053_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1053_addr];
  `endif
  assign tgtPages_T_1058_addr = 6'h22;
  assign tgtPages_T_1058_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1058_data = tgtPages[tgtPages_T_1058_addr];
  `else
  assign tgtPages_T_1058_data = tgtPages_T_1058_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1058_addr];
  `endif
  assign tgtPages_T_1063_addr = 6'h23;
  assign tgtPages_T_1063_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1063_data = tgtPages[tgtPages_T_1063_addr];
  `else
  assign tgtPages_T_1063_data = tgtPages_T_1063_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1063_addr];
  `endif
  assign tgtPages_T_1068_addr = 6'h24;
  assign tgtPages_T_1068_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1068_data = tgtPages[tgtPages_T_1068_addr];
  `else
  assign tgtPages_T_1068_data = tgtPages_T_1068_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1068_addr];
  `endif
  assign tgtPages_T_1073_addr = 6'h25;
  assign tgtPages_T_1073_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1073_data = tgtPages[tgtPages_T_1073_addr];
  `else
  assign tgtPages_T_1073_data = tgtPages_T_1073_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1073_addr];
  `endif
  assign tgtPages_T_1078_addr = 6'h26;
  assign tgtPages_T_1078_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1078_data = tgtPages[tgtPages_T_1078_addr];
  `else
  assign tgtPages_T_1078_data = tgtPages_T_1078_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1078_addr];
  `endif
  assign tgtPages_T_1083_addr = 6'h27;
  assign tgtPages_T_1083_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1083_data = tgtPages[tgtPages_T_1083_addr];
  `else
  assign tgtPages_T_1083_data = tgtPages_T_1083_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1083_addr];
  `endif
  assign tgtPages_T_1088_addr = 6'h28;
  assign tgtPages_T_1088_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1088_data = tgtPages[tgtPages_T_1088_addr];
  `else
  assign tgtPages_T_1088_data = tgtPages_T_1088_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1088_addr];
  `endif
  assign tgtPages_T_1093_addr = 6'h29;
  assign tgtPages_T_1093_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1093_data = tgtPages[tgtPages_T_1093_addr];
  `else
  assign tgtPages_T_1093_data = tgtPages_T_1093_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1093_addr];
  `endif
  assign tgtPages_T_1098_addr = 6'h2a;
  assign tgtPages_T_1098_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1098_data = tgtPages[tgtPages_T_1098_addr];
  `else
  assign tgtPages_T_1098_data = tgtPages_T_1098_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1098_addr];
  `endif
  assign tgtPages_T_1103_addr = 6'h2b;
  assign tgtPages_T_1103_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1103_data = tgtPages[tgtPages_T_1103_addr];
  `else
  assign tgtPages_T_1103_data = tgtPages_T_1103_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1103_addr];
  `endif
  assign tgtPages_T_1108_addr = 6'h2c;
  assign tgtPages_T_1108_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1108_data = tgtPages[tgtPages_T_1108_addr];
  `else
  assign tgtPages_T_1108_data = tgtPages_T_1108_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1108_addr];
  `endif
  assign tgtPages_T_1113_addr = 6'h2d;
  assign tgtPages_T_1113_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1113_data = tgtPages[tgtPages_T_1113_addr];
  `else
  assign tgtPages_T_1113_data = tgtPages_T_1113_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1113_addr];
  `endif
  assign tgtPages_T_1118_addr = 6'h2e;
  assign tgtPages_T_1118_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1118_data = tgtPages[tgtPages_T_1118_addr];
  `else
  assign tgtPages_T_1118_data = tgtPages_T_1118_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1118_addr];
  `endif
  assign tgtPages_T_1123_addr = 6'h2f;
  assign tgtPages_T_1123_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1123_data = tgtPages[tgtPages_T_1123_addr];
  `else
  assign tgtPages_T_1123_data = tgtPages_T_1123_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1123_addr];
  `endif
  assign tgtPages_T_1128_addr = 6'h30;
  assign tgtPages_T_1128_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1128_data = tgtPages[tgtPages_T_1128_addr];
  `else
  assign tgtPages_T_1128_data = tgtPages_T_1128_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1128_addr];
  `endif
  assign tgtPages_T_1133_addr = 6'h31;
  assign tgtPages_T_1133_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1133_data = tgtPages[tgtPages_T_1133_addr];
  `else
  assign tgtPages_T_1133_data = tgtPages_T_1133_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1133_addr];
  `endif
  assign tgtPages_T_1138_addr = 6'h32;
  assign tgtPages_T_1138_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1138_data = tgtPages[tgtPages_T_1138_addr];
  `else
  assign tgtPages_T_1138_data = tgtPages_T_1138_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1138_addr];
  `endif
  assign tgtPages_T_1143_addr = 6'h33;
  assign tgtPages_T_1143_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1143_data = tgtPages[tgtPages_T_1143_addr];
  `else
  assign tgtPages_T_1143_data = tgtPages_T_1143_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1143_addr];
  `endif
  assign tgtPages_T_1148_addr = 6'h34;
  assign tgtPages_T_1148_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1148_data = tgtPages[tgtPages_T_1148_addr];
  `else
  assign tgtPages_T_1148_data = tgtPages_T_1148_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1148_addr];
  `endif
  assign tgtPages_T_1153_addr = 6'h35;
  assign tgtPages_T_1153_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1153_data = tgtPages[tgtPages_T_1153_addr];
  `else
  assign tgtPages_T_1153_data = tgtPages_T_1153_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1153_addr];
  `endif
  assign tgtPages_T_1158_addr = 6'h36;
  assign tgtPages_T_1158_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1158_data = tgtPages[tgtPages_T_1158_addr];
  `else
  assign tgtPages_T_1158_data = tgtPages_T_1158_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1158_addr];
  `endif
  assign tgtPages_T_1163_addr = 6'h37;
  assign tgtPages_T_1163_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1163_data = tgtPages[tgtPages_T_1163_addr];
  `else
  assign tgtPages_T_1163_data = tgtPages_T_1163_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1163_addr];
  `endif
  assign tgtPages_T_1168_addr = 6'h38;
  assign tgtPages_T_1168_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1168_data = tgtPages[tgtPages_T_1168_addr];
  `else
  assign tgtPages_T_1168_data = tgtPages_T_1168_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1168_addr];
  `endif
  assign tgtPages_T_1173_addr = 6'h39;
  assign tgtPages_T_1173_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1173_data = tgtPages[tgtPages_T_1173_addr];
  `else
  assign tgtPages_T_1173_data = tgtPages_T_1173_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1173_addr];
  `endif
  assign tgtPages_T_1178_addr = 6'h3a;
  assign tgtPages_T_1178_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1178_data = tgtPages[tgtPages_T_1178_addr];
  `else
  assign tgtPages_T_1178_data = tgtPages_T_1178_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1178_addr];
  `endif
  assign tgtPages_T_1183_addr = 6'h3b;
  assign tgtPages_T_1183_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1183_data = tgtPages[tgtPages_T_1183_addr];
  `else
  assign tgtPages_T_1183_data = tgtPages_T_1183_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1183_addr];
  `endif
  assign tgtPages_T_1188_addr = 6'h3c;
  assign tgtPages_T_1188_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1188_data = tgtPages[tgtPages_T_1188_addr];
  `else
  assign tgtPages_T_1188_data = tgtPages_T_1188_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1188_addr];
  `endif
  assign tgtPages_T_1193_addr = 6'h3d;
  assign tgtPages_T_1193_en = 1'h1;
  `ifdef SYNTHESIS
  assign tgtPages_T_1193_data = tgtPages[tgtPages_T_1193_addr];
  `else
  assign tgtPages_T_1193_data = tgtPages_T_1193_addr >= 6'h3e ? $random : tgtPages[tgtPages_T_1193_addr];
  `endif
  assign tgtPages_T_2875_data = tgtPageUpdate;
  assign tgtPages_T_2875_addr = T_2550;
  assign tgtPages_T_2875_mask = r_btb_update_valid;
  assign tgtPages_T_2875_en = r_btb_update_valid;
  assign pages_T_1400_addr = {{2'd0}, 1'h0};
  assign pages_T_1400_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1400_data = pages[pages_T_1400_addr];
  `else
  assign pages_T_1400_data = pages_T_1400_addr >= 3'h6 ? $random : pages[pages_T_1400_addr];
  `endif
  assign pages_T_1403_addr = {{2'd0}, 1'h1};
  assign pages_T_1403_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1403_data = pages[pages_T_1403_addr];
  `else
  assign pages_T_1403_data = pages_T_1403_addr >= 3'h6 ? $random : pages[pages_T_1403_addr];
  `endif
  assign pages_T_1406_addr = {{1'd0}, 2'h2};
  assign pages_T_1406_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1406_data = pages[pages_T_1406_addr];
  `else
  assign pages_T_1406_data = pages_T_1406_addr >= 3'h6 ? $random : pages[pages_T_1406_addr];
  `endif
  assign pages_T_1409_addr = {{1'd0}, 2'h3};
  assign pages_T_1409_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1409_data = pages[pages_T_1409_addr];
  `else
  assign pages_T_1409_data = pages_T_1409_addr >= 3'h6 ? $random : pages[pages_T_1409_addr];
  `endif
  assign pages_T_1412_addr = 3'h4;
  assign pages_T_1412_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1412_data = pages[pages_T_1412_addr];
  `else
  assign pages_T_1412_data = pages_T_1412_addr >= 3'h6 ? $random : pages[pages_T_1412_addr];
  `endif
  assign pages_T_1415_addr = 3'h5;
  assign pages_T_1415_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1415_data = pages[pages_T_1415_addr];
  `else
  assign pages_T_1415_data = pages_T_1415_addr >= 3'h6 ? $random : pages[pages_T_1415_addr];
  `endif
  assign pages_T_1941_addr = {{2'd0}, 1'h0};
  assign pages_T_1941_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1941_data = pages[pages_T_1941_addr];
  `else
  assign pages_T_1941_data = pages_T_1941_addr >= 3'h6 ? $random : pages[pages_T_1941_addr];
  `endif
  assign pages_T_1944_addr = {{2'd0}, 1'h1};
  assign pages_T_1944_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1944_data = pages[pages_T_1944_addr];
  `else
  assign pages_T_1944_data = pages_T_1944_addr >= 3'h6 ? $random : pages[pages_T_1944_addr];
  `endif
  assign pages_T_1947_addr = {{1'd0}, 2'h2};
  assign pages_T_1947_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1947_data = pages[pages_T_1947_addr];
  `else
  assign pages_T_1947_data = pages_T_1947_addr >= 3'h6 ? $random : pages[pages_T_1947_addr];
  `endif
  assign pages_T_1950_addr = {{1'd0}, 2'h3};
  assign pages_T_1950_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1950_data = pages[pages_T_1950_addr];
  `else
  assign pages_T_1950_data = pages_T_1950_addr >= 3'h6 ? $random : pages[pages_T_1950_addr];
  `endif
  assign pages_T_1953_addr = 3'h4;
  assign pages_T_1953_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1953_data = pages[pages_T_1953_addr];
  `else
  assign pages_T_1953_data = pages_T_1953_addr >= 3'h6 ? $random : pages[pages_T_1953_addr];
  `endif
  assign pages_T_1956_addr = 3'h5;
  assign pages_T_1956_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_1956_data = pages[pages_T_1956_addr];
  `else
  assign pages_T_1956_data = pages_T_1956_addr >= 3'h6 ? $random : pages[pages_T_1956_addr];
  `endif
  assign pages_T_3177_addr = {{2'd0}, 1'h0};
  assign pages_T_3177_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3177_data = pages[pages_T_3177_addr];
  `else
  assign pages_T_3177_data = pages_T_3177_addr >= 3'h6 ? $random : pages[pages_T_3177_addr];
  `endif
  assign pages_T_3179_addr = {{2'd0}, 1'h1};
  assign pages_T_3179_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3179_data = pages[pages_T_3179_addr];
  `else
  assign pages_T_3179_data = pages_T_3179_addr >= 3'h6 ? $random : pages[pages_T_3179_addr];
  `endif
  assign pages_T_3181_addr = {{1'd0}, 2'h2};
  assign pages_T_3181_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3181_data = pages[pages_T_3181_addr];
  `else
  assign pages_T_3181_data = pages_T_3181_addr >= 3'h6 ? $random : pages[pages_T_3181_addr];
  `endif
  assign pages_T_3183_addr = {{1'd0}, 2'h3};
  assign pages_T_3183_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3183_data = pages[pages_T_3183_addr];
  `else
  assign pages_T_3183_data = pages_T_3183_addr >= 3'h6 ? $random : pages[pages_T_3183_addr];
  `endif
  assign pages_T_3185_addr = 3'h4;
  assign pages_T_3185_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3185_data = pages[pages_T_3185_addr];
  `else
  assign pages_T_3185_data = pages_T_3185_addr >= 3'h6 ? $random : pages[pages_T_3185_addr];
  `endif
  assign pages_T_3187_addr = 3'h5;
  assign pages_T_3187_en = 1'h1;
  `ifdef SYNTHESIS
  assign pages_T_3187_data = pages[pages_T_3187_addr];
  `else
  assign pages_T_3187_data = pages_T_3187_addr >= 3'h6 ? $random : pages[pages_T_3187_addr];
  `endif
  assign pages_T_2891_data = T_2887;
  assign pages_T_2891_addr = {{2'd0}, 1'h0};
  assign pages_T_2891_mask = GEN_393;
  assign pages_T_2891_en = GEN_393;
  assign pages_T_2895_data = T_2887;
  assign pages_T_2895_addr = {{1'd0}, 2'h2};
  assign pages_T_2895_mask = GEN_398;
  assign pages_T_2895_en = GEN_398;
  assign pages_T_2899_data = T_2887;
  assign pages_T_2899_addr = 3'h4;
  assign pages_T_2899_mask = GEN_403;
  assign pages_T_2899_en = GEN_403;
  assign pages_T_2907_data = T_2903;
  assign pages_T_2907_addr = {{2'd0}, 1'h1};
  assign pages_T_2907_mask = GEN_408;
  assign pages_T_2907_en = GEN_408;
  assign pages_T_2911_data = T_2903;
  assign pages_T_2911_addr = {{1'd0}, 2'h3};
  assign pages_T_2911_mask = GEN_413;
  assign pages_T_2911_en = GEN_413;
  assign pages_T_2915_data = T_2903;
  assign pages_T_2915_addr = 3'h5;
  assign pages_T_2915_mask = GEN_418;
  assign pages_T_2915_en = GEN_418;
  assign GEN_457 = {{7'd0}, 1'h1};
  assign T_580 = GEN_457 << idxPages_T_578_data;
  assign T_581 = T_580[5:0];
  assign T_585 = GEN_457 << idxPages_T_583_data;
  assign T_586 = T_585[5:0];
  assign T_590 = GEN_457 << idxPages_T_588_data;
  assign T_591 = T_590[5:0];
  assign T_595 = GEN_457 << idxPages_T_593_data;
  assign T_596 = T_595[5:0];
  assign T_600 = GEN_457 << idxPages_T_598_data;
  assign T_601 = T_600[5:0];
  assign T_605 = GEN_457 << idxPages_T_603_data;
  assign T_606 = T_605[5:0];
  assign T_610 = GEN_457 << idxPages_T_608_data;
  assign T_611 = T_610[5:0];
  assign T_615 = GEN_457 << idxPages_T_613_data;
  assign T_616 = T_615[5:0];
  assign T_620 = GEN_457 << idxPages_T_618_data;
  assign T_621 = T_620[5:0];
  assign T_625 = GEN_457 << idxPages_T_623_data;
  assign T_626 = T_625[5:0];
  assign T_630 = GEN_457 << idxPages_T_628_data;
  assign T_631 = T_630[5:0];
  assign T_635 = GEN_457 << idxPages_T_633_data;
  assign T_636 = T_635[5:0];
  assign T_640 = GEN_457 << idxPages_T_638_data;
  assign T_641 = T_640[5:0];
  assign T_645 = GEN_457 << idxPages_T_643_data;
  assign T_646 = T_645[5:0];
  assign T_650 = GEN_457 << idxPages_T_648_data;
  assign T_651 = T_650[5:0];
  assign T_655 = GEN_457 << idxPages_T_653_data;
  assign T_656 = T_655[5:0];
  assign T_660 = GEN_457 << idxPages_T_658_data;
  assign T_661 = T_660[5:0];
  assign T_665 = GEN_457 << idxPages_T_663_data;
  assign T_666 = T_665[5:0];
  assign T_670 = GEN_457 << idxPages_T_668_data;
  assign T_671 = T_670[5:0];
  assign T_675 = GEN_457 << idxPages_T_673_data;
  assign T_676 = T_675[5:0];
  assign T_680 = GEN_457 << idxPages_T_678_data;
  assign T_681 = T_680[5:0];
  assign T_685 = GEN_457 << idxPages_T_683_data;
  assign T_686 = T_685[5:0];
  assign T_690 = GEN_457 << idxPages_T_688_data;
  assign T_691 = T_690[5:0];
  assign T_695 = GEN_457 << idxPages_T_693_data;
  assign T_696 = T_695[5:0];
  assign T_700 = GEN_457 << idxPages_T_698_data;
  assign T_701 = T_700[5:0];
  assign T_705 = GEN_457 << idxPages_T_703_data;
  assign T_706 = T_705[5:0];
  assign T_710 = GEN_457 << idxPages_T_708_data;
  assign T_711 = T_710[5:0];
  assign T_715 = GEN_457 << idxPages_T_713_data;
  assign T_716 = T_715[5:0];
  assign T_720 = GEN_457 << idxPages_T_718_data;
  assign T_721 = T_720[5:0];
  assign T_725 = GEN_457 << idxPages_T_723_data;
  assign T_726 = T_725[5:0];
  assign T_730 = GEN_457 << idxPages_T_728_data;
  assign T_731 = T_730[5:0];
  assign T_735 = GEN_457 << idxPages_T_733_data;
  assign T_736 = T_735[5:0];
  assign T_740 = GEN_457 << idxPages_T_738_data;
  assign T_741 = T_740[5:0];
  assign T_745 = GEN_457 << idxPages_T_743_data;
  assign T_746 = T_745[5:0];
  assign T_750 = GEN_457 << idxPages_T_748_data;
  assign T_751 = T_750[5:0];
  assign T_755 = GEN_457 << idxPages_T_753_data;
  assign T_756 = T_755[5:0];
  assign T_760 = GEN_457 << idxPages_T_758_data;
  assign T_761 = T_760[5:0];
  assign T_765 = GEN_457 << idxPages_T_763_data;
  assign T_766 = T_765[5:0];
  assign T_770 = GEN_457 << idxPages_T_768_data;
  assign T_771 = T_770[5:0];
  assign T_775 = GEN_457 << idxPages_T_773_data;
  assign T_776 = T_775[5:0];
  assign T_780 = GEN_457 << idxPages_T_778_data;
  assign T_781 = T_780[5:0];
  assign T_785 = GEN_457 << idxPages_T_783_data;
  assign T_786 = T_785[5:0];
  assign T_790 = GEN_457 << idxPages_T_788_data;
  assign T_791 = T_790[5:0];
  assign T_795 = GEN_457 << idxPages_T_793_data;
  assign T_796 = T_795[5:0];
  assign T_800 = GEN_457 << idxPages_T_798_data;
  assign T_801 = T_800[5:0];
  assign T_805 = GEN_457 << idxPages_T_803_data;
  assign T_806 = T_805[5:0];
  assign T_810 = GEN_457 << idxPages_T_808_data;
  assign T_811 = T_810[5:0];
  assign T_815 = GEN_457 << idxPages_T_813_data;
  assign T_816 = T_815[5:0];
  assign T_820 = GEN_457 << idxPages_T_818_data;
  assign T_821 = T_820[5:0];
  assign T_825 = GEN_457 << idxPages_T_823_data;
  assign T_826 = T_825[5:0];
  assign T_830 = GEN_457 << idxPages_T_828_data;
  assign T_831 = T_830[5:0];
  assign T_835 = GEN_457 << idxPages_T_833_data;
  assign T_836 = T_835[5:0];
  assign T_840 = GEN_457 << idxPages_T_838_data;
  assign T_841 = T_840[5:0];
  assign T_845 = GEN_457 << idxPages_T_843_data;
  assign T_846 = T_845[5:0];
  assign T_850 = GEN_457 << idxPages_T_848_data;
  assign T_851 = T_850[5:0];
  assign T_855 = GEN_457 << idxPages_T_853_data;
  assign T_856 = T_855[5:0];
  assign T_860 = GEN_457 << idxPages_T_858_data;
  assign T_861 = T_860[5:0];
  assign T_865 = GEN_457 << idxPages_T_863_data;
  assign T_866 = T_865[5:0];
  assign T_870 = GEN_457 << idxPages_T_868_data;
  assign T_871 = T_870[5:0];
  assign T_875 = GEN_457 << idxPages_T_873_data;
  assign T_876 = T_875[5:0];
  assign T_880 = GEN_457 << idxPages_T_878_data;
  assign T_881 = T_880[5:0];
  assign T_885 = GEN_457 << idxPages_T_883_data;
  assign T_886 = T_885[5:0];
  assign T_890 = GEN_457 << tgtPages_T_888_data;
  assign T_891 = T_890[5:0];
  assign T_895 = GEN_457 << tgtPages_T_893_data;
  assign T_896 = T_895[5:0];
  assign T_900 = GEN_457 << tgtPages_T_898_data;
  assign T_901 = T_900[5:0];
  assign T_905 = GEN_457 << tgtPages_T_903_data;
  assign T_906 = T_905[5:0];
  assign T_910 = GEN_457 << tgtPages_T_908_data;
  assign T_911 = T_910[5:0];
  assign T_915 = GEN_457 << tgtPages_T_913_data;
  assign T_916 = T_915[5:0];
  assign T_920 = GEN_457 << tgtPages_T_918_data;
  assign T_921 = T_920[5:0];
  assign T_925 = GEN_457 << tgtPages_T_923_data;
  assign T_926 = T_925[5:0];
  assign T_930 = GEN_457 << tgtPages_T_928_data;
  assign T_931 = T_930[5:0];
  assign T_935 = GEN_457 << tgtPages_T_933_data;
  assign T_936 = T_935[5:0];
  assign T_940 = GEN_457 << tgtPages_T_938_data;
  assign T_941 = T_940[5:0];
  assign T_945 = GEN_457 << tgtPages_T_943_data;
  assign T_946 = T_945[5:0];
  assign T_950 = GEN_457 << tgtPages_T_948_data;
  assign T_951 = T_950[5:0];
  assign T_955 = GEN_457 << tgtPages_T_953_data;
  assign T_956 = T_955[5:0];
  assign T_960 = GEN_457 << tgtPages_T_958_data;
  assign T_961 = T_960[5:0];
  assign T_965 = GEN_457 << tgtPages_T_963_data;
  assign T_966 = T_965[5:0];
  assign T_970 = GEN_457 << tgtPages_T_968_data;
  assign T_971 = T_970[5:0];
  assign T_975 = GEN_457 << tgtPages_T_973_data;
  assign T_976 = T_975[5:0];
  assign T_980 = GEN_457 << tgtPages_T_978_data;
  assign T_981 = T_980[5:0];
  assign T_985 = GEN_457 << tgtPages_T_983_data;
  assign T_986 = T_985[5:0];
  assign T_990 = GEN_457 << tgtPages_T_988_data;
  assign T_991 = T_990[5:0];
  assign T_995 = GEN_457 << tgtPages_T_993_data;
  assign T_996 = T_995[5:0];
  assign T_1000 = GEN_457 << tgtPages_T_998_data;
  assign T_1001 = T_1000[5:0];
  assign T_1005 = GEN_457 << tgtPages_T_1003_data;
  assign T_1006 = T_1005[5:0];
  assign T_1010 = GEN_457 << tgtPages_T_1008_data;
  assign T_1011 = T_1010[5:0];
  assign T_1015 = GEN_457 << tgtPages_T_1013_data;
  assign T_1016 = T_1015[5:0];
  assign T_1020 = GEN_457 << tgtPages_T_1018_data;
  assign T_1021 = T_1020[5:0];
  assign T_1025 = GEN_457 << tgtPages_T_1023_data;
  assign T_1026 = T_1025[5:0];
  assign T_1030 = GEN_457 << tgtPages_T_1028_data;
  assign T_1031 = T_1030[5:0];
  assign T_1035 = GEN_457 << tgtPages_T_1033_data;
  assign T_1036 = T_1035[5:0];
  assign T_1040 = GEN_457 << tgtPages_T_1038_data;
  assign T_1041 = T_1040[5:0];
  assign T_1045 = GEN_457 << tgtPages_T_1043_data;
  assign T_1046 = T_1045[5:0];
  assign T_1050 = GEN_457 << tgtPages_T_1048_data;
  assign T_1051 = T_1050[5:0];
  assign T_1055 = GEN_457 << tgtPages_T_1053_data;
  assign T_1056 = T_1055[5:0];
  assign T_1060 = GEN_457 << tgtPages_T_1058_data;
  assign T_1061 = T_1060[5:0];
  assign T_1065 = GEN_457 << tgtPages_T_1063_data;
  assign T_1066 = T_1065[5:0];
  assign T_1070 = GEN_457 << tgtPages_T_1068_data;
  assign T_1071 = T_1070[5:0];
  assign T_1075 = GEN_457 << tgtPages_T_1073_data;
  assign T_1076 = T_1075[5:0];
  assign T_1080 = GEN_457 << tgtPages_T_1078_data;
  assign T_1081 = T_1080[5:0];
  assign T_1085 = GEN_457 << tgtPages_T_1083_data;
  assign T_1086 = T_1085[5:0];
  assign T_1090 = GEN_457 << tgtPages_T_1088_data;
  assign T_1091 = T_1090[5:0];
  assign T_1095 = GEN_457 << tgtPages_T_1093_data;
  assign T_1096 = T_1095[5:0];
  assign T_1100 = GEN_457 << tgtPages_T_1098_data;
  assign T_1101 = T_1100[5:0];
  assign T_1105 = GEN_457 << tgtPages_T_1103_data;
  assign T_1106 = T_1105[5:0];
  assign T_1110 = GEN_457 << tgtPages_T_1108_data;
  assign T_1111 = T_1110[5:0];
  assign T_1115 = GEN_457 << tgtPages_T_1113_data;
  assign T_1116 = T_1115[5:0];
  assign T_1120 = GEN_457 << tgtPages_T_1118_data;
  assign T_1121 = T_1120[5:0];
  assign T_1125 = GEN_457 << tgtPages_T_1123_data;
  assign T_1126 = T_1125[5:0];
  assign T_1130 = GEN_457 << tgtPages_T_1128_data;
  assign T_1131 = T_1130[5:0];
  assign T_1135 = GEN_457 << tgtPages_T_1133_data;
  assign T_1136 = T_1135[5:0];
  assign T_1140 = GEN_457 << tgtPages_T_1138_data;
  assign T_1141 = T_1140[5:0];
  assign T_1145 = GEN_457 << tgtPages_T_1143_data;
  assign T_1146 = T_1145[5:0];
  assign T_1150 = GEN_457 << tgtPages_T_1148_data;
  assign T_1151 = T_1150[5:0];
  assign T_1155 = GEN_457 << tgtPages_T_1153_data;
  assign T_1156 = T_1155[5:0];
  assign T_1160 = GEN_457 << tgtPages_T_1158_data;
  assign T_1161 = T_1160[5:0];
  assign T_1165 = GEN_457 << tgtPages_T_1163_data;
  assign T_1166 = T_1165[5:0];
  assign T_1170 = GEN_457 << tgtPages_T_1168_data;
  assign T_1171 = T_1170[5:0];
  assign T_1175 = GEN_457 << tgtPages_T_1173_data;
  assign T_1176 = T_1175[5:0];
  assign T_1180 = GEN_457 << tgtPages_T_1178_data;
  assign T_1181 = T_1180[5:0];
  assign T_1185 = GEN_457 << tgtPages_T_1183_data;
  assign T_1186 = T_1185[5:0];
  assign T_1190 = GEN_457 << tgtPages_T_1188_data;
  assign T_1191 = T_1190[5:0];
  assign T_1195 = GEN_457 << tgtPages_T_1193_data;
  assign T_1196 = T_1195[5:0];
  assign brIdx_T_3612_addr = io_resp_bits_entry;
  assign brIdx_T_3612_en = 1'h1;
  `ifdef SYNTHESIS
  assign brIdx_T_3612_data = brIdx[brIdx_T_3612_addr];
  `else
  assign brIdx_T_3612_data = brIdx_T_3612_addr >= 6'h3e ? $random : brIdx[brIdx_T_3612_addr];
  `endif
  assign brIdx_T_2876_data = 1'h0;
  assign brIdx_T_2876_addr = T_2550;
  assign brIdx_T_2876_mask = r_btb_update_valid;
  assign brIdx_T_2876_en = r_btb_update_valid;
  assign GEN_4 = io_btb_update_valid ? io_btb_update_bits_prediction_valid : T_1216_prediction_valid;
  assign GEN_5 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_taken : T_1216_prediction_bits_taken;
  assign GEN_6 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_mask : T_1216_prediction_bits_mask;
  assign GEN_7 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bridx : T_1216_prediction_bits_bridx;
  assign GEN_8 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_target : T_1216_prediction_bits_target;
  assign GEN_9 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_entry : T_1216_prediction_bits_entry;
  assign GEN_10 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_history : T_1216_prediction_bits_bht_history;
  assign GEN_11 = io_btb_update_valid ? io_btb_update_bits_prediction_bits_bht_value : T_1216_prediction_bits_bht_value;
  assign GEN_12 = io_btb_update_valid ? io_btb_update_bits_pc : T_1216_pc;
  assign GEN_13 = io_btb_update_valid ? io_btb_update_bits_target : T_1216_target;
  assign GEN_14 = io_btb_update_valid ? io_btb_update_bits_taken : T_1216_taken;
  assign GEN_15 = io_btb_update_valid ? io_btb_update_bits_isJump : T_1216_isJump;
  assign GEN_16 = io_btb_update_valid ? io_btb_update_bits_isReturn : T_1216_isReturn;
  assign GEN_17 = io_btb_update_valid ? io_btb_update_bits_br_pc : T_1216_br_pc;
  assign r_btb_update_valid = T_1215;
  assign r_btb_update_bits_prediction_valid = T_1216_prediction_valid;
  assign r_btb_update_bits_prediction_bits_taken = T_1216_prediction_bits_taken;
  assign r_btb_update_bits_prediction_bits_mask = T_1216_prediction_bits_mask;
  assign r_btb_update_bits_prediction_bits_bridx = T_1216_prediction_bits_bridx;
  assign r_btb_update_bits_prediction_bits_target = T_1216_prediction_bits_target;
  assign r_btb_update_bits_prediction_bits_entry = T_1216_prediction_bits_entry;
  assign r_btb_update_bits_prediction_bits_bht_history = T_1216_prediction_bits_bht_history;
  assign r_btb_update_bits_prediction_bits_bht_value = T_1216_prediction_bits_bht_value;
  assign r_btb_update_bits_pc = T_1216_pc;
  assign r_btb_update_bits_target = T_1216_target;
  assign r_btb_update_bits_taken = T_1216_taken;
  assign r_btb_update_bits_isJump = T_1216_isJump;
  assign r_btb_update_bits_isReturn = T_1216_isReturn;
  assign r_btb_update_bits_br_pc = T_1216_br_pc;
  assign T_1398 = io_req_bits_addr[38:12];
  assign T_1401 = pages_T_1400_data == T_1398;
  assign T_1404 = pages_T_1403_data == T_1398;
  assign T_1407 = pages_T_1406_data == T_1398;
  assign T_1410 = pages_T_1409_data == T_1398;
  assign T_1413 = pages_T_1412_data == T_1398;
  assign T_1416 = pages_T_1415_data == T_1398;
  assign T_1422_0 = T_1401;
  assign T_1422_1 = T_1404;
  assign T_1422_2 = T_1407;
  assign T_1422_3 = T_1410;
  assign T_1422_4 = T_1413;
  assign T_1422_5 = T_1416;
  assign T_1424 = {T_1422_2,T_1422_1};
  assign T_1425 = {T_1424,T_1422_0};
  assign T_1426 = {T_1422_5,T_1422_4};
  assign T_1427 = {T_1426,T_1422_3};
  assign T_1428 = {T_1427,T_1425};
  assign pageHit = T_1428 & pageValid;
  assign T_1429 = io_req_bits_addr[11:0];
  assign T_1432 = idxs_T_1431_data == T_1429;
  assign T_1435 = idxs_T_1434_data == T_1429;
  assign T_1438 = idxs_T_1437_data == T_1429;
  assign T_1441 = idxs_T_1440_data == T_1429;
  assign T_1444 = idxs_T_1443_data == T_1429;
  assign T_1447 = idxs_T_1446_data == T_1429;
  assign T_1450 = idxs_T_1449_data == T_1429;
  assign T_1453 = idxs_T_1452_data == T_1429;
  assign T_1456 = idxs_T_1455_data == T_1429;
  assign T_1459 = idxs_T_1458_data == T_1429;
  assign T_1462 = idxs_T_1461_data == T_1429;
  assign T_1465 = idxs_T_1464_data == T_1429;
  assign T_1468 = idxs_T_1467_data == T_1429;
  assign T_1471 = idxs_T_1470_data == T_1429;
  assign T_1474 = idxs_T_1473_data == T_1429;
  assign T_1477 = idxs_T_1476_data == T_1429;
  assign T_1480 = idxs_T_1479_data == T_1429;
  assign T_1483 = idxs_T_1482_data == T_1429;
  assign T_1486 = idxs_T_1485_data == T_1429;
  assign T_1489 = idxs_T_1488_data == T_1429;
  assign T_1492 = idxs_T_1491_data == T_1429;
  assign T_1495 = idxs_T_1494_data == T_1429;
  assign T_1498 = idxs_T_1497_data == T_1429;
  assign T_1501 = idxs_T_1500_data == T_1429;
  assign T_1504 = idxs_T_1503_data == T_1429;
  assign T_1507 = idxs_T_1506_data == T_1429;
  assign T_1510 = idxs_T_1509_data == T_1429;
  assign T_1513 = idxs_T_1512_data == T_1429;
  assign T_1516 = idxs_T_1515_data == T_1429;
  assign T_1519 = idxs_T_1518_data == T_1429;
  assign T_1522 = idxs_T_1521_data == T_1429;
  assign T_1525 = idxs_T_1524_data == T_1429;
  assign T_1528 = idxs_T_1527_data == T_1429;
  assign T_1531 = idxs_T_1530_data == T_1429;
  assign T_1534 = idxs_T_1533_data == T_1429;
  assign T_1537 = idxs_T_1536_data == T_1429;
  assign T_1540 = idxs_T_1539_data == T_1429;
  assign T_1543 = idxs_T_1542_data == T_1429;
  assign T_1546 = idxs_T_1545_data == T_1429;
  assign T_1549 = idxs_T_1548_data == T_1429;
  assign T_1552 = idxs_T_1551_data == T_1429;
  assign T_1555 = idxs_T_1554_data == T_1429;
  assign T_1558 = idxs_T_1557_data == T_1429;
  assign T_1561 = idxs_T_1560_data == T_1429;
  assign T_1564 = idxs_T_1563_data == T_1429;
  assign T_1567 = idxs_T_1566_data == T_1429;
  assign T_1570 = idxs_T_1569_data == T_1429;
  assign T_1573 = idxs_T_1572_data == T_1429;
  assign T_1576 = idxs_T_1575_data == T_1429;
  assign T_1579 = idxs_T_1578_data == T_1429;
  assign T_1582 = idxs_T_1581_data == T_1429;
  assign T_1585 = idxs_T_1584_data == T_1429;
  assign T_1588 = idxs_T_1587_data == T_1429;
  assign T_1591 = idxs_T_1590_data == T_1429;
  assign T_1594 = idxs_T_1593_data == T_1429;
  assign T_1597 = idxs_T_1596_data == T_1429;
  assign T_1600 = idxs_T_1599_data == T_1429;
  assign T_1603 = idxs_T_1602_data == T_1429;
  assign T_1606 = idxs_T_1605_data == T_1429;
  assign T_1609 = idxs_T_1608_data == T_1429;
  assign T_1612 = idxs_T_1611_data == T_1429;
  assign T_1615 = idxs_T_1614_data == T_1429;
  assign T_1621_0 = T_1432;
  assign T_1621_1 = T_1435;
  assign T_1621_2 = T_1438;
  assign T_1621_3 = T_1441;
  assign T_1621_4 = T_1444;
  assign T_1621_5 = T_1447;
  assign T_1621_6 = T_1450;
  assign T_1621_7 = T_1453;
  assign T_1621_8 = T_1456;
  assign T_1621_9 = T_1459;
  assign T_1621_10 = T_1462;
  assign T_1621_11 = T_1465;
  assign T_1621_12 = T_1468;
  assign T_1621_13 = T_1471;
  assign T_1621_14 = T_1474;
  assign T_1621_15 = T_1477;
  assign T_1621_16 = T_1480;
  assign T_1621_17 = T_1483;
  assign T_1621_18 = T_1486;
  assign T_1621_19 = T_1489;
  assign T_1621_20 = T_1492;
  assign T_1621_21 = T_1495;
  assign T_1621_22 = T_1498;
  assign T_1621_23 = T_1501;
  assign T_1621_24 = T_1504;
  assign T_1621_25 = T_1507;
  assign T_1621_26 = T_1510;
  assign T_1621_27 = T_1513;
  assign T_1621_28 = T_1516;
  assign T_1621_29 = T_1519;
  assign T_1621_30 = T_1522;
  assign T_1621_31 = T_1525;
  assign T_1621_32 = T_1528;
  assign T_1621_33 = T_1531;
  assign T_1621_34 = T_1534;
  assign T_1621_35 = T_1537;
  assign T_1621_36 = T_1540;
  assign T_1621_37 = T_1543;
  assign T_1621_38 = T_1546;
  assign T_1621_39 = T_1549;
  assign T_1621_40 = T_1552;
  assign T_1621_41 = T_1555;
  assign T_1621_42 = T_1558;
  assign T_1621_43 = T_1561;
  assign T_1621_44 = T_1564;
  assign T_1621_45 = T_1567;
  assign T_1621_46 = T_1570;
  assign T_1621_47 = T_1573;
  assign T_1621_48 = T_1576;
  assign T_1621_49 = T_1579;
  assign T_1621_50 = T_1582;
  assign T_1621_51 = T_1585;
  assign T_1621_52 = T_1588;
  assign T_1621_53 = T_1591;
  assign T_1621_54 = T_1594;
  assign T_1621_55 = T_1597;
  assign T_1621_56 = T_1600;
  assign T_1621_57 = T_1603;
  assign T_1621_58 = T_1606;
  assign T_1621_59 = T_1609;
  assign T_1621_60 = T_1612;
  assign T_1621_61 = T_1615;
  assign T_1623 = {T_1621_2,T_1621_1};
  assign T_1624 = {T_1623,T_1621_0};
  assign T_1625 = {T_1621_4,T_1621_3};
  assign T_1626 = {T_1621_6,T_1621_5};
  assign T_1627 = {T_1626,T_1625};
  assign T_1628 = {T_1627,T_1624};
  assign T_1629 = {T_1621_8,T_1621_7};
  assign T_1630 = {T_1621_10,T_1621_9};
  assign T_1631 = {T_1630,T_1629};
  assign T_1632 = {T_1621_12,T_1621_11};
  assign T_1633 = {T_1621_14,T_1621_13};
  assign T_1634 = {T_1633,T_1632};
  assign T_1635 = {T_1634,T_1631};
  assign T_1636 = {T_1635,T_1628};
  assign T_1637 = {T_1621_16,T_1621_15};
  assign T_1638 = {T_1621_18,T_1621_17};
  assign T_1639 = {T_1638,T_1637};
  assign T_1640 = {T_1621_20,T_1621_19};
  assign T_1641 = {T_1621_22,T_1621_21};
  assign T_1642 = {T_1641,T_1640};
  assign T_1643 = {T_1642,T_1639};
  assign T_1644 = {T_1621_24,T_1621_23};
  assign T_1645 = {T_1621_26,T_1621_25};
  assign T_1646 = {T_1645,T_1644};
  assign T_1647 = {T_1621_28,T_1621_27};
  assign T_1648 = {T_1621_30,T_1621_29};
  assign T_1649 = {T_1648,T_1647};
  assign T_1650 = {T_1649,T_1646};
  assign T_1651 = {T_1650,T_1643};
  assign T_1652 = {T_1651,T_1636};
  assign T_1653 = {T_1621_33,T_1621_32};
  assign T_1654 = {T_1653,T_1621_31};
  assign T_1655 = {T_1621_35,T_1621_34};
  assign T_1656 = {T_1621_37,T_1621_36};
  assign T_1657 = {T_1656,T_1655};
  assign T_1658 = {T_1657,T_1654};
  assign T_1659 = {T_1621_39,T_1621_38};
  assign T_1660 = {T_1621_41,T_1621_40};
  assign T_1661 = {T_1660,T_1659};
  assign T_1662 = {T_1621_43,T_1621_42};
  assign T_1663 = {T_1621_45,T_1621_44};
  assign T_1664 = {T_1663,T_1662};
  assign T_1665 = {T_1664,T_1661};
  assign T_1666 = {T_1665,T_1658};
  assign T_1667 = {T_1621_47,T_1621_46};
  assign T_1668 = {T_1621_49,T_1621_48};
  assign T_1669 = {T_1668,T_1667};
  assign T_1670 = {T_1621_51,T_1621_50};
  assign T_1671 = {T_1621_53,T_1621_52};
  assign T_1672 = {T_1671,T_1670};
  assign T_1673 = {T_1672,T_1669};
  assign T_1674 = {T_1621_55,T_1621_54};
  assign T_1675 = {T_1621_57,T_1621_56};
  assign T_1676 = {T_1675,T_1674};
  assign T_1677 = {T_1621_59,T_1621_58};
  assign T_1678 = {T_1621_61,T_1621_60};
  assign T_1679 = {T_1678,T_1677};
  assign T_1680 = {T_1679,T_1676};
  assign T_1681 = {T_1680,T_1673};
  assign T_1682 = {T_1681,T_1666};
  assign T_1683 = {T_1682,T_1652};
  assign T_1684 = T_581 & pageHit;
  assign T_1685 = T_586 & pageHit;
  assign T_1686 = T_591 & pageHit;
  assign T_1687 = T_596 & pageHit;
  assign T_1688 = T_601 & pageHit;
  assign T_1689 = T_606 & pageHit;
  assign T_1690 = T_611 & pageHit;
  assign T_1691 = T_616 & pageHit;
  assign T_1692 = T_621 & pageHit;
  assign T_1693 = T_626 & pageHit;
  assign T_1694 = T_631 & pageHit;
  assign T_1695 = T_636 & pageHit;
  assign T_1696 = T_641 & pageHit;
  assign T_1697 = T_646 & pageHit;
  assign T_1698 = T_651 & pageHit;
  assign T_1699 = T_656 & pageHit;
  assign T_1700 = T_661 & pageHit;
  assign T_1701 = T_666 & pageHit;
  assign T_1702 = T_671 & pageHit;
  assign T_1703 = T_676 & pageHit;
  assign T_1704 = T_681 & pageHit;
  assign T_1705 = T_686 & pageHit;
  assign T_1706 = T_691 & pageHit;
  assign T_1707 = T_696 & pageHit;
  assign T_1708 = T_701 & pageHit;
  assign T_1709 = T_706 & pageHit;
  assign T_1710 = T_711 & pageHit;
  assign T_1711 = T_716 & pageHit;
  assign T_1712 = T_721 & pageHit;
  assign T_1713 = T_726 & pageHit;
  assign T_1714 = T_731 & pageHit;
  assign T_1715 = T_736 & pageHit;
  assign T_1716 = T_741 & pageHit;
  assign T_1717 = T_746 & pageHit;
  assign T_1718 = T_751 & pageHit;
  assign T_1719 = T_756 & pageHit;
  assign T_1720 = T_761 & pageHit;
  assign T_1721 = T_766 & pageHit;
  assign T_1722 = T_771 & pageHit;
  assign T_1723 = T_776 & pageHit;
  assign T_1724 = T_781 & pageHit;
  assign T_1725 = T_786 & pageHit;
  assign T_1726 = T_791 & pageHit;
  assign T_1727 = T_796 & pageHit;
  assign T_1728 = T_801 & pageHit;
  assign T_1729 = T_806 & pageHit;
  assign T_1730 = T_811 & pageHit;
  assign T_1731 = T_816 & pageHit;
  assign T_1732 = T_821 & pageHit;
  assign T_1733 = T_826 & pageHit;
  assign T_1734 = T_831 & pageHit;
  assign T_1735 = T_836 & pageHit;
  assign T_1736 = T_841 & pageHit;
  assign T_1737 = T_846 & pageHit;
  assign T_1738 = T_851 & pageHit;
  assign T_1739 = T_856 & pageHit;
  assign T_1740 = T_861 & pageHit;
  assign T_1741 = T_866 & pageHit;
  assign T_1742 = T_871 & pageHit;
  assign T_1743 = T_876 & pageHit;
  assign T_1744 = T_881 & pageHit;
  assign T_1745 = T_886 & pageHit;
  assign GEN_581 = {{5'd0}, 1'h0};
  assign T_1747 = T_1684 != GEN_581;
  assign T_1749 = T_1685 != GEN_581;
  assign T_1751 = T_1686 != GEN_581;
  assign T_1753 = T_1687 != GEN_581;
  assign T_1755 = T_1688 != GEN_581;
  assign T_1757 = T_1689 != GEN_581;
  assign T_1759 = T_1690 != GEN_581;
  assign T_1761 = T_1691 != GEN_581;
  assign T_1763 = T_1692 != GEN_581;
  assign T_1765 = T_1693 != GEN_581;
  assign T_1767 = T_1694 != GEN_581;
  assign T_1769 = T_1695 != GEN_581;
  assign T_1771 = T_1696 != GEN_581;
  assign T_1773 = T_1697 != GEN_581;
  assign T_1775 = T_1698 != GEN_581;
  assign T_1777 = T_1699 != GEN_581;
  assign T_1779 = T_1700 != GEN_581;
  assign T_1781 = T_1701 != GEN_581;
  assign T_1783 = T_1702 != GEN_581;
  assign T_1785 = T_1703 != GEN_581;
  assign T_1787 = T_1704 != GEN_581;
  assign T_1789 = T_1705 != GEN_581;
  assign T_1791 = T_1706 != GEN_581;
  assign T_1793 = T_1707 != GEN_581;
  assign T_1795 = T_1708 != GEN_581;
  assign T_1797 = T_1709 != GEN_581;
  assign T_1799 = T_1710 != GEN_581;
  assign T_1801 = T_1711 != GEN_581;
  assign T_1803 = T_1712 != GEN_581;
  assign T_1805 = T_1713 != GEN_581;
  assign T_1807 = T_1714 != GEN_581;
  assign T_1809 = T_1715 != GEN_581;
  assign T_1811 = T_1716 != GEN_581;
  assign T_1813 = T_1717 != GEN_581;
  assign T_1815 = T_1718 != GEN_581;
  assign T_1817 = T_1719 != GEN_581;
  assign T_1819 = T_1720 != GEN_581;
  assign T_1821 = T_1721 != GEN_581;
  assign T_1823 = T_1722 != GEN_581;
  assign T_1825 = T_1723 != GEN_581;
  assign T_1827 = T_1724 != GEN_581;
  assign T_1829 = T_1725 != GEN_581;
  assign T_1831 = T_1726 != GEN_581;
  assign T_1833 = T_1727 != GEN_581;
  assign T_1835 = T_1728 != GEN_581;
  assign T_1837 = T_1729 != GEN_581;
  assign T_1839 = T_1730 != GEN_581;
  assign T_1841 = T_1731 != GEN_581;
  assign T_1843 = T_1732 != GEN_581;
  assign T_1845 = T_1733 != GEN_581;
  assign T_1847 = T_1734 != GEN_581;
  assign T_1849 = T_1735 != GEN_581;
  assign T_1851 = T_1736 != GEN_581;
  assign T_1853 = T_1737 != GEN_581;
  assign T_1855 = T_1738 != GEN_581;
  assign T_1857 = T_1739 != GEN_581;
  assign T_1859 = T_1740 != GEN_581;
  assign T_1861 = T_1741 != GEN_581;
  assign T_1863 = T_1742 != GEN_581;
  assign T_1865 = T_1743 != GEN_581;
  assign T_1867 = T_1744 != GEN_581;
  assign T_1869 = T_1745 != GEN_581;
  assign T_1875_0 = T_1747;
  assign T_1875_1 = T_1749;
  assign T_1875_2 = T_1751;
  assign T_1875_3 = T_1753;
  assign T_1875_4 = T_1755;
  assign T_1875_5 = T_1757;
  assign T_1875_6 = T_1759;
  assign T_1875_7 = T_1761;
  assign T_1875_8 = T_1763;
  assign T_1875_9 = T_1765;
  assign T_1875_10 = T_1767;
  assign T_1875_11 = T_1769;
  assign T_1875_12 = T_1771;
  assign T_1875_13 = T_1773;
  assign T_1875_14 = T_1775;
  assign T_1875_15 = T_1777;
  assign T_1875_16 = T_1779;
  assign T_1875_17 = T_1781;
  assign T_1875_18 = T_1783;
  assign T_1875_19 = T_1785;
  assign T_1875_20 = T_1787;
  assign T_1875_21 = T_1789;
  assign T_1875_22 = T_1791;
  assign T_1875_23 = T_1793;
  assign T_1875_24 = T_1795;
  assign T_1875_25 = T_1797;
  assign T_1875_26 = T_1799;
  assign T_1875_27 = T_1801;
  assign T_1875_28 = T_1803;
  assign T_1875_29 = T_1805;
  assign T_1875_30 = T_1807;
  assign T_1875_31 = T_1809;
  assign T_1875_32 = T_1811;
  assign T_1875_33 = T_1813;
  assign T_1875_34 = T_1815;
  assign T_1875_35 = T_1817;
  assign T_1875_36 = T_1819;
  assign T_1875_37 = T_1821;
  assign T_1875_38 = T_1823;
  assign T_1875_39 = T_1825;
  assign T_1875_40 = T_1827;
  assign T_1875_41 = T_1829;
  assign T_1875_42 = T_1831;
  assign T_1875_43 = T_1833;
  assign T_1875_44 = T_1835;
  assign T_1875_45 = T_1837;
  assign T_1875_46 = T_1839;
  assign T_1875_47 = T_1841;
  assign T_1875_48 = T_1843;
  assign T_1875_49 = T_1845;
  assign T_1875_50 = T_1847;
  assign T_1875_51 = T_1849;
  assign T_1875_52 = T_1851;
  assign T_1875_53 = T_1853;
  assign T_1875_54 = T_1855;
  assign T_1875_55 = T_1857;
  assign T_1875_56 = T_1859;
  assign T_1875_57 = T_1861;
  assign T_1875_58 = T_1863;
  assign T_1875_59 = T_1865;
  assign T_1875_60 = T_1867;
  assign T_1875_61 = T_1869;
  assign T_1877 = {T_1875_2,T_1875_1};
  assign T_1878 = {T_1877,T_1875_0};
  assign T_1879 = {T_1875_4,T_1875_3};
  assign T_1880 = {T_1875_6,T_1875_5};
  assign T_1881 = {T_1880,T_1879};
  assign T_1882 = {T_1881,T_1878};
  assign T_1883 = {T_1875_8,T_1875_7};
  assign T_1884 = {T_1875_10,T_1875_9};
  assign T_1885 = {T_1884,T_1883};
  assign T_1886 = {T_1875_12,T_1875_11};
  assign T_1887 = {T_1875_14,T_1875_13};
  assign T_1888 = {T_1887,T_1886};
  assign T_1889 = {T_1888,T_1885};
  assign T_1890 = {T_1889,T_1882};
  assign T_1891 = {T_1875_16,T_1875_15};
  assign T_1892 = {T_1875_18,T_1875_17};
  assign T_1893 = {T_1892,T_1891};
  assign T_1894 = {T_1875_20,T_1875_19};
  assign T_1895 = {T_1875_22,T_1875_21};
  assign T_1896 = {T_1895,T_1894};
  assign T_1897 = {T_1896,T_1893};
  assign T_1898 = {T_1875_24,T_1875_23};
  assign T_1899 = {T_1875_26,T_1875_25};
  assign T_1900 = {T_1899,T_1898};
  assign T_1901 = {T_1875_28,T_1875_27};
  assign T_1902 = {T_1875_30,T_1875_29};
  assign T_1903 = {T_1902,T_1901};
  assign T_1904 = {T_1903,T_1900};
  assign T_1905 = {T_1904,T_1897};
  assign T_1906 = {T_1905,T_1890};
  assign T_1907 = {T_1875_33,T_1875_32};
  assign T_1908 = {T_1907,T_1875_31};
  assign T_1909 = {T_1875_35,T_1875_34};
  assign T_1910 = {T_1875_37,T_1875_36};
  assign T_1911 = {T_1910,T_1909};
  assign T_1912 = {T_1911,T_1908};
  assign T_1913 = {T_1875_39,T_1875_38};
  assign T_1914 = {T_1875_41,T_1875_40};
  assign T_1915 = {T_1914,T_1913};
  assign T_1916 = {T_1875_43,T_1875_42};
  assign T_1917 = {T_1875_45,T_1875_44};
  assign T_1918 = {T_1917,T_1916};
  assign T_1919 = {T_1918,T_1915};
  assign T_1920 = {T_1919,T_1912};
  assign T_1921 = {T_1875_47,T_1875_46};
  assign T_1922 = {T_1875_49,T_1875_48};
  assign T_1923 = {T_1922,T_1921};
  assign T_1924 = {T_1875_51,T_1875_50};
  assign T_1925 = {T_1875_53,T_1875_52};
  assign T_1926 = {T_1925,T_1924};
  assign T_1927 = {T_1926,T_1923};
  assign T_1928 = {T_1875_55,T_1875_54};
  assign T_1929 = {T_1875_57,T_1875_56};
  assign T_1930 = {T_1929,T_1928};
  assign T_1931 = {T_1875_59,T_1875_58};
  assign T_1932 = {T_1875_61,T_1875_60};
  assign T_1933 = {T_1932,T_1931};
  assign T_1934 = {T_1933,T_1930};
  assign T_1935 = {T_1934,T_1927};
  assign T_1936 = {T_1935,T_1920};
  assign T_1937 = {T_1936,T_1906};
  assign T_1938 = idxValid & T_1683;
  assign hits = T_1938 & T_1937;
  assign T_1939 = r_btb_update_bits_pc[38:12];
  assign T_1942 = pages_T_1941_data == T_1939;
  assign T_1945 = pages_T_1944_data == T_1939;
  assign T_1948 = pages_T_1947_data == T_1939;
  assign T_1951 = pages_T_1950_data == T_1939;
  assign T_1954 = pages_T_1953_data == T_1939;
  assign T_1957 = pages_T_1956_data == T_1939;
  assign T_1963_0 = T_1942;
  assign T_1963_1 = T_1945;
  assign T_1963_2 = T_1948;
  assign T_1963_3 = T_1951;
  assign T_1963_4 = T_1954;
  assign T_1963_5 = T_1957;
  assign T_1965 = {T_1963_2,T_1963_1};
  assign T_1966 = {T_1965,T_1963_0};
  assign T_1967 = {T_1963_5,T_1963_4};
  assign T_1968 = {T_1967,T_1963_3};
  assign T_1969 = {T_1968,T_1966};
  assign updatePageHit = T_1969 & pageValid;
  assign T_1970 = r_btb_update_bits_pc[11:0];
  assign T_1973 = idxs_T_1972_data == T_1970;
  assign T_1976 = idxs_T_1975_data == T_1970;
  assign T_1979 = idxs_T_1978_data == T_1970;
  assign T_1982 = idxs_T_1981_data == T_1970;
  assign T_1985 = idxs_T_1984_data == T_1970;
  assign T_1988 = idxs_T_1987_data == T_1970;
  assign T_1991 = idxs_T_1990_data == T_1970;
  assign T_1994 = idxs_T_1993_data == T_1970;
  assign T_1997 = idxs_T_1996_data == T_1970;
  assign T_2000 = idxs_T_1999_data == T_1970;
  assign T_2003 = idxs_T_2002_data == T_1970;
  assign T_2006 = idxs_T_2005_data == T_1970;
  assign T_2009 = idxs_T_2008_data == T_1970;
  assign T_2012 = idxs_T_2011_data == T_1970;
  assign T_2015 = idxs_T_2014_data == T_1970;
  assign T_2018 = idxs_T_2017_data == T_1970;
  assign T_2021 = idxs_T_2020_data == T_1970;
  assign T_2024 = idxs_T_2023_data == T_1970;
  assign T_2027 = idxs_T_2026_data == T_1970;
  assign T_2030 = idxs_T_2029_data == T_1970;
  assign T_2033 = idxs_T_2032_data == T_1970;
  assign T_2036 = idxs_T_2035_data == T_1970;
  assign T_2039 = idxs_T_2038_data == T_1970;
  assign T_2042 = idxs_T_2041_data == T_1970;
  assign T_2045 = idxs_T_2044_data == T_1970;
  assign T_2048 = idxs_T_2047_data == T_1970;
  assign T_2051 = idxs_T_2050_data == T_1970;
  assign T_2054 = idxs_T_2053_data == T_1970;
  assign T_2057 = idxs_T_2056_data == T_1970;
  assign T_2060 = idxs_T_2059_data == T_1970;
  assign T_2063 = idxs_T_2062_data == T_1970;
  assign T_2066 = idxs_T_2065_data == T_1970;
  assign T_2069 = idxs_T_2068_data == T_1970;
  assign T_2072 = idxs_T_2071_data == T_1970;
  assign T_2075 = idxs_T_2074_data == T_1970;
  assign T_2078 = idxs_T_2077_data == T_1970;
  assign T_2081 = idxs_T_2080_data == T_1970;
  assign T_2084 = idxs_T_2083_data == T_1970;
  assign T_2087 = idxs_T_2086_data == T_1970;
  assign T_2090 = idxs_T_2089_data == T_1970;
  assign T_2093 = idxs_T_2092_data == T_1970;
  assign T_2096 = idxs_T_2095_data == T_1970;
  assign T_2099 = idxs_T_2098_data == T_1970;
  assign T_2102 = idxs_T_2101_data == T_1970;
  assign T_2105 = idxs_T_2104_data == T_1970;
  assign T_2108 = idxs_T_2107_data == T_1970;
  assign T_2111 = idxs_T_2110_data == T_1970;
  assign T_2114 = idxs_T_2113_data == T_1970;
  assign T_2117 = idxs_T_2116_data == T_1970;
  assign T_2120 = idxs_T_2119_data == T_1970;
  assign T_2123 = idxs_T_2122_data == T_1970;
  assign T_2126 = idxs_T_2125_data == T_1970;
  assign T_2129 = idxs_T_2128_data == T_1970;
  assign T_2132 = idxs_T_2131_data == T_1970;
  assign T_2135 = idxs_T_2134_data == T_1970;
  assign T_2138 = idxs_T_2137_data == T_1970;
  assign T_2141 = idxs_T_2140_data == T_1970;
  assign T_2144 = idxs_T_2143_data == T_1970;
  assign T_2147 = idxs_T_2146_data == T_1970;
  assign T_2150 = idxs_T_2149_data == T_1970;
  assign T_2153 = idxs_T_2152_data == T_1970;
  assign T_2156 = idxs_T_2155_data == T_1970;
  assign T_2162_0 = T_1973;
  assign T_2162_1 = T_1976;
  assign T_2162_2 = T_1979;
  assign T_2162_3 = T_1982;
  assign T_2162_4 = T_1985;
  assign T_2162_5 = T_1988;
  assign T_2162_6 = T_1991;
  assign T_2162_7 = T_1994;
  assign T_2162_8 = T_1997;
  assign T_2162_9 = T_2000;
  assign T_2162_10 = T_2003;
  assign T_2162_11 = T_2006;
  assign T_2162_12 = T_2009;
  assign T_2162_13 = T_2012;
  assign T_2162_14 = T_2015;
  assign T_2162_15 = T_2018;
  assign T_2162_16 = T_2021;
  assign T_2162_17 = T_2024;
  assign T_2162_18 = T_2027;
  assign T_2162_19 = T_2030;
  assign T_2162_20 = T_2033;
  assign T_2162_21 = T_2036;
  assign T_2162_22 = T_2039;
  assign T_2162_23 = T_2042;
  assign T_2162_24 = T_2045;
  assign T_2162_25 = T_2048;
  assign T_2162_26 = T_2051;
  assign T_2162_27 = T_2054;
  assign T_2162_28 = T_2057;
  assign T_2162_29 = T_2060;
  assign T_2162_30 = T_2063;
  assign T_2162_31 = T_2066;
  assign T_2162_32 = T_2069;
  assign T_2162_33 = T_2072;
  assign T_2162_34 = T_2075;
  assign T_2162_35 = T_2078;
  assign T_2162_36 = T_2081;
  assign T_2162_37 = T_2084;
  assign T_2162_38 = T_2087;
  assign T_2162_39 = T_2090;
  assign T_2162_40 = T_2093;
  assign T_2162_41 = T_2096;
  assign T_2162_42 = T_2099;
  assign T_2162_43 = T_2102;
  assign T_2162_44 = T_2105;
  assign T_2162_45 = T_2108;
  assign T_2162_46 = T_2111;
  assign T_2162_47 = T_2114;
  assign T_2162_48 = T_2117;
  assign T_2162_49 = T_2120;
  assign T_2162_50 = T_2123;
  assign T_2162_51 = T_2126;
  assign T_2162_52 = T_2129;
  assign T_2162_53 = T_2132;
  assign T_2162_54 = T_2135;
  assign T_2162_55 = T_2138;
  assign T_2162_56 = T_2141;
  assign T_2162_57 = T_2144;
  assign T_2162_58 = T_2147;
  assign T_2162_59 = T_2150;
  assign T_2162_60 = T_2153;
  assign T_2162_61 = T_2156;
  assign T_2225 = T_581 & updatePageHit;
  assign T_2226 = T_586 & updatePageHit;
  assign T_2227 = T_591 & updatePageHit;
  assign T_2228 = T_596 & updatePageHit;
  assign T_2229 = T_601 & updatePageHit;
  assign T_2230 = T_606 & updatePageHit;
  assign T_2231 = T_611 & updatePageHit;
  assign T_2232 = T_616 & updatePageHit;
  assign T_2233 = T_621 & updatePageHit;
  assign T_2234 = T_626 & updatePageHit;
  assign T_2235 = T_631 & updatePageHit;
  assign T_2236 = T_636 & updatePageHit;
  assign T_2237 = T_641 & updatePageHit;
  assign T_2238 = T_646 & updatePageHit;
  assign T_2239 = T_651 & updatePageHit;
  assign T_2240 = T_656 & updatePageHit;
  assign T_2241 = T_661 & updatePageHit;
  assign T_2242 = T_666 & updatePageHit;
  assign T_2243 = T_671 & updatePageHit;
  assign T_2244 = T_676 & updatePageHit;
  assign T_2245 = T_681 & updatePageHit;
  assign T_2246 = T_686 & updatePageHit;
  assign T_2247 = T_691 & updatePageHit;
  assign T_2248 = T_696 & updatePageHit;
  assign T_2249 = T_701 & updatePageHit;
  assign T_2250 = T_706 & updatePageHit;
  assign T_2251 = T_711 & updatePageHit;
  assign T_2252 = T_716 & updatePageHit;
  assign T_2253 = T_721 & updatePageHit;
  assign T_2254 = T_726 & updatePageHit;
  assign T_2255 = T_731 & updatePageHit;
  assign T_2256 = T_736 & updatePageHit;
  assign T_2257 = T_741 & updatePageHit;
  assign T_2258 = T_746 & updatePageHit;
  assign T_2259 = T_751 & updatePageHit;
  assign T_2260 = T_756 & updatePageHit;
  assign T_2261 = T_761 & updatePageHit;
  assign T_2262 = T_766 & updatePageHit;
  assign T_2263 = T_771 & updatePageHit;
  assign T_2264 = T_776 & updatePageHit;
  assign T_2265 = T_781 & updatePageHit;
  assign T_2266 = T_786 & updatePageHit;
  assign T_2267 = T_791 & updatePageHit;
  assign T_2268 = T_796 & updatePageHit;
  assign T_2269 = T_801 & updatePageHit;
  assign T_2270 = T_806 & updatePageHit;
  assign T_2271 = T_811 & updatePageHit;
  assign T_2272 = T_816 & updatePageHit;
  assign T_2273 = T_821 & updatePageHit;
  assign T_2274 = T_826 & updatePageHit;
  assign T_2275 = T_831 & updatePageHit;
  assign T_2276 = T_836 & updatePageHit;
  assign T_2277 = T_841 & updatePageHit;
  assign T_2278 = T_846 & updatePageHit;
  assign T_2279 = T_851 & updatePageHit;
  assign T_2280 = T_856 & updatePageHit;
  assign T_2281 = T_861 & updatePageHit;
  assign T_2282 = T_866 & updatePageHit;
  assign T_2283 = T_871 & updatePageHit;
  assign T_2284 = T_876 & updatePageHit;
  assign T_2285 = T_881 & updatePageHit;
  assign T_2286 = T_886 & updatePageHit;
  assign T_2288 = T_2225 != GEN_581;
  assign T_2290 = T_2226 != GEN_581;
  assign T_2292 = T_2227 != GEN_581;
  assign T_2294 = T_2228 != GEN_581;
  assign T_2296 = T_2229 != GEN_581;
  assign T_2298 = T_2230 != GEN_581;
  assign T_2300 = T_2231 != GEN_581;
  assign T_2302 = T_2232 != GEN_581;
  assign T_2304 = T_2233 != GEN_581;
  assign T_2306 = T_2234 != GEN_581;
  assign T_2308 = T_2235 != GEN_581;
  assign T_2310 = T_2236 != GEN_581;
  assign T_2312 = T_2237 != GEN_581;
  assign T_2314 = T_2238 != GEN_581;
  assign T_2316 = T_2239 != GEN_581;
  assign T_2318 = T_2240 != GEN_581;
  assign T_2320 = T_2241 != GEN_581;
  assign T_2322 = T_2242 != GEN_581;
  assign T_2324 = T_2243 != GEN_581;
  assign T_2326 = T_2244 != GEN_581;
  assign T_2328 = T_2245 != GEN_581;
  assign T_2330 = T_2246 != GEN_581;
  assign T_2332 = T_2247 != GEN_581;
  assign T_2334 = T_2248 != GEN_581;
  assign T_2336 = T_2249 != GEN_581;
  assign T_2338 = T_2250 != GEN_581;
  assign T_2340 = T_2251 != GEN_581;
  assign T_2342 = T_2252 != GEN_581;
  assign T_2344 = T_2253 != GEN_581;
  assign T_2346 = T_2254 != GEN_581;
  assign T_2348 = T_2255 != GEN_581;
  assign T_2350 = T_2256 != GEN_581;
  assign T_2352 = T_2257 != GEN_581;
  assign T_2354 = T_2258 != GEN_581;
  assign T_2356 = T_2259 != GEN_581;
  assign T_2358 = T_2260 != GEN_581;
  assign T_2360 = T_2261 != GEN_581;
  assign T_2362 = T_2262 != GEN_581;
  assign T_2364 = T_2263 != GEN_581;
  assign T_2366 = T_2264 != GEN_581;
  assign T_2368 = T_2265 != GEN_581;
  assign T_2370 = T_2266 != GEN_581;
  assign T_2372 = T_2267 != GEN_581;
  assign T_2374 = T_2268 != GEN_581;
  assign T_2376 = T_2269 != GEN_581;
  assign T_2378 = T_2270 != GEN_581;
  assign T_2380 = T_2271 != GEN_581;
  assign T_2382 = T_2272 != GEN_581;
  assign T_2384 = T_2273 != GEN_581;
  assign T_2386 = T_2274 != GEN_581;
  assign T_2388 = T_2275 != GEN_581;
  assign T_2390 = T_2276 != GEN_581;
  assign T_2392 = T_2277 != GEN_581;
  assign T_2394 = T_2278 != GEN_581;
  assign T_2396 = T_2279 != GEN_581;
  assign T_2398 = T_2280 != GEN_581;
  assign T_2400 = T_2281 != GEN_581;
  assign T_2402 = T_2282 != GEN_581;
  assign T_2404 = T_2283 != GEN_581;
  assign T_2406 = T_2284 != GEN_581;
  assign T_2408 = T_2285 != GEN_581;
  assign T_2410 = T_2286 != GEN_581;
  assign T_2416_0 = T_2288;
  assign T_2416_1 = T_2290;
  assign T_2416_2 = T_2292;
  assign T_2416_3 = T_2294;
  assign T_2416_4 = T_2296;
  assign T_2416_5 = T_2298;
  assign T_2416_6 = T_2300;
  assign T_2416_7 = T_2302;
  assign T_2416_8 = T_2304;
  assign T_2416_9 = T_2306;
  assign T_2416_10 = T_2308;
  assign T_2416_11 = T_2310;
  assign T_2416_12 = T_2312;
  assign T_2416_13 = T_2314;
  assign T_2416_14 = T_2316;
  assign T_2416_15 = T_2318;
  assign T_2416_16 = T_2320;
  assign T_2416_17 = T_2322;
  assign T_2416_18 = T_2324;
  assign T_2416_19 = T_2326;
  assign T_2416_20 = T_2328;
  assign T_2416_21 = T_2330;
  assign T_2416_22 = T_2332;
  assign T_2416_23 = T_2334;
  assign T_2416_24 = T_2336;
  assign T_2416_25 = T_2338;
  assign T_2416_26 = T_2340;
  assign T_2416_27 = T_2342;
  assign T_2416_28 = T_2344;
  assign T_2416_29 = T_2346;
  assign T_2416_30 = T_2348;
  assign T_2416_31 = T_2350;
  assign T_2416_32 = T_2352;
  assign T_2416_33 = T_2354;
  assign T_2416_34 = T_2356;
  assign T_2416_35 = T_2358;
  assign T_2416_36 = T_2360;
  assign T_2416_37 = T_2362;
  assign T_2416_38 = T_2364;
  assign T_2416_39 = T_2366;
  assign T_2416_40 = T_2368;
  assign T_2416_41 = T_2370;
  assign T_2416_42 = T_2372;
  assign T_2416_43 = T_2374;
  assign T_2416_44 = T_2376;
  assign T_2416_45 = T_2378;
  assign T_2416_46 = T_2380;
  assign T_2416_47 = T_2382;
  assign T_2416_48 = T_2384;
  assign T_2416_49 = T_2386;
  assign T_2416_50 = T_2388;
  assign T_2416_51 = T_2390;
  assign T_2416_52 = T_2392;
  assign T_2416_53 = T_2394;
  assign T_2416_54 = T_2396;
  assign T_2416_55 = T_2398;
  assign T_2416_56 = T_2400;
  assign T_2416_57 = T_2402;
  assign T_2416_58 = T_2404;
  assign T_2416_59 = T_2406;
  assign T_2416_60 = T_2408;
  assign T_2416_61 = T_2410;
  assign T_2481 = r_btb_update_bits_prediction_valid == 1'h0;
  assign T_2482 = r_btb_update_valid & T_2481;
  assign T_2485 = nextRepl == 6'h3d;
  assign GEN_705 = {{5'd0}, 1'h1};
  assign T_2487 = nextRepl + GEN_705;
  assign T_2488 = T_2487[5:0];
  assign GEN_18 = T_2485 ? {{5'd0}, 1'h0} : T_2488;
  assign GEN_19 = T_2482 ? GEN_18 : nextRepl;
  assign useUpdatePageHit = updatePageHit != GEN_581;
  assign doIdxPageRepl = useUpdatePageHit == 1'h0;
  assign idxPageRepl = T_2545[5:0];
  assign idxPageUpdateOH = useUpdatePageHit ? updatePageHit : idxPageRepl;
  assign T_2494 = idxPageUpdateOH[5:4];
  assign T_2495 = idxPageUpdateOH[3:0];
  assign GEN_707 = {{1'd0}, 1'h0};
  assign T_2497 = T_2494 != GEN_707;
  assign GEN_708 = {{2'd0}, T_2494};
  assign T_2498 = GEN_708 | T_2495;
  assign T_2499 = T_2498[3:2];
  assign T_2500 = T_2498[1:0];
  assign T_2502 = T_2499 != GEN_707;
  assign T_2503 = T_2499 | T_2500;
  assign T_2504 = T_2503[1];
  assign T_2505 = {T_2502,T_2504};
  assign idxPageUpdate = {T_2497,T_2505};
  assign idxPageReplEn = doIdxPageRepl ? idxPageRepl : {{5'd0}, 1'h0};
  assign samePage = T_1939 == T_1398;
  assign T_2509 = ~ idxPageReplEn;
  assign T_2510 = pageHit & T_2509;
  assign usePageHit = T_2510 != GEN_581;
  assign T_2513 = samePage == 1'h0;
  assign T_2515 = usePageHit == 1'h0;
  assign doTgtPageRepl = T_2513 & T_2515;
  assign T_2516 = idxPageUpdateOH[4:0];
  assign GEN_711 = {{1'd0}, T_2516};
  assign T_2517 = GEN_711 << 1;
  assign T_2518 = idxPageUpdateOH[5];
  assign GEN_712 = {{5'd0}, T_2518};
  assign T_2519 = T_2517 | GEN_712;
  assign tgtPageRepl = samePage ? idxPageUpdateOH : T_2519;
  assign T_2520 = usePageHit ? pageHit : tgtPageRepl;
  assign T_2521 = T_2520[5:4];
  assign T_2522 = T_2520[3:0];
  assign T_2524 = T_2521 != GEN_707;
  assign GEN_714 = {{2'd0}, T_2521};
  assign T_2525 = GEN_714 | T_2522;
  assign T_2526 = T_2525[3:2];
  assign T_2527 = T_2525[1:0];
  assign T_2529 = T_2526 != GEN_707;
  assign T_2530 = T_2526 | T_2527;
  assign T_2531 = T_2530[1];
  assign T_2532 = {T_2529,T_2531};
  assign tgtPageUpdate = {T_2524,T_2532};
  assign tgtPageReplEn = doTgtPageRepl ? tgtPageRepl : {{5'd0}, 1'h0};
  assign doPageRepl = doIdxPageRepl | doTgtPageRepl;
  assign pageReplEn = idxPageReplEn | tgtPageReplEn;
  assign T_2534 = r_btb_update_valid & doPageRepl;
  assign T_2538 = T_2536 == 3'h5;
  assign GEN_716 = {{2'd0}, 1'h1};
  assign T_2540 = T_2536 + GEN_716;
  assign T_2541 = T_2540[2:0];
  assign GEN_20 = T_2538 ? {{2'd0}, 1'h0} : T_2541;
  assign GEN_21 = T_2534 ? GEN_20 : T_2536;
  assign T_2545 = GEN_457 << T_2536;
  assign T_2546 = io_req_bits_addr == r_btb_update_bits_target;
  assign T_2547 = T_2546 | reset;
  assign T_2549 = T_2547 == 1'h0;
  assign T_2550 = r_btb_update_bits_prediction_valid ? r_btb_update_bits_prediction_bits_entry : nextRepl;
  assign T_2551 = T_581 | T_891;
  assign T_2552 = pageReplEn & T_2551;
  assign T_2554 = T_2552 != GEN_581;
  assign T_2555 = T_586 | T_896;
  assign T_2556 = pageReplEn & T_2555;
  assign T_2558 = T_2556 != GEN_581;
  assign T_2559 = T_591 | T_901;
  assign T_2560 = pageReplEn & T_2559;
  assign T_2562 = T_2560 != GEN_581;
  assign T_2563 = T_596 | T_906;
  assign T_2564 = pageReplEn & T_2563;
  assign T_2566 = T_2564 != GEN_581;
  assign T_2567 = T_601 | T_911;
  assign T_2568 = pageReplEn & T_2567;
  assign T_2570 = T_2568 != GEN_581;
  assign T_2571 = T_606 | T_916;
  assign T_2572 = pageReplEn & T_2571;
  assign T_2574 = T_2572 != GEN_581;
  assign T_2575 = T_611 | T_921;
  assign T_2576 = pageReplEn & T_2575;
  assign T_2578 = T_2576 != GEN_581;
  assign T_2579 = T_616 | T_926;
  assign T_2580 = pageReplEn & T_2579;
  assign T_2582 = T_2580 != GEN_581;
  assign T_2583 = T_621 | T_931;
  assign T_2584 = pageReplEn & T_2583;
  assign T_2586 = T_2584 != GEN_581;
  assign T_2587 = T_626 | T_936;
  assign T_2588 = pageReplEn & T_2587;
  assign T_2590 = T_2588 != GEN_581;
  assign T_2591 = T_631 | T_941;
  assign T_2592 = pageReplEn & T_2591;
  assign T_2594 = T_2592 != GEN_581;
  assign T_2595 = T_636 | T_946;
  assign T_2596 = pageReplEn & T_2595;
  assign T_2598 = T_2596 != GEN_581;
  assign T_2599 = T_641 | T_951;
  assign T_2600 = pageReplEn & T_2599;
  assign T_2602 = T_2600 != GEN_581;
  assign T_2603 = T_646 | T_956;
  assign T_2604 = pageReplEn & T_2603;
  assign T_2606 = T_2604 != GEN_581;
  assign T_2607 = T_651 | T_961;
  assign T_2608 = pageReplEn & T_2607;
  assign T_2610 = T_2608 != GEN_581;
  assign T_2611 = T_656 | T_966;
  assign T_2612 = pageReplEn & T_2611;
  assign T_2614 = T_2612 != GEN_581;
  assign T_2615 = T_661 | T_971;
  assign T_2616 = pageReplEn & T_2615;
  assign T_2618 = T_2616 != GEN_581;
  assign T_2619 = T_666 | T_976;
  assign T_2620 = pageReplEn & T_2619;
  assign T_2622 = T_2620 != GEN_581;
  assign T_2623 = T_671 | T_981;
  assign T_2624 = pageReplEn & T_2623;
  assign T_2626 = T_2624 != GEN_581;
  assign T_2627 = T_676 | T_986;
  assign T_2628 = pageReplEn & T_2627;
  assign T_2630 = T_2628 != GEN_581;
  assign T_2631 = T_681 | T_991;
  assign T_2632 = pageReplEn & T_2631;
  assign T_2634 = T_2632 != GEN_581;
  assign T_2635 = T_686 | T_996;
  assign T_2636 = pageReplEn & T_2635;
  assign T_2638 = T_2636 != GEN_581;
  assign T_2639 = T_691 | T_1001;
  assign T_2640 = pageReplEn & T_2639;
  assign T_2642 = T_2640 != GEN_581;
  assign T_2643 = T_696 | T_1006;
  assign T_2644 = pageReplEn & T_2643;
  assign T_2646 = T_2644 != GEN_581;
  assign T_2647 = T_701 | T_1011;
  assign T_2648 = pageReplEn & T_2647;
  assign T_2650 = T_2648 != GEN_581;
  assign T_2651 = T_706 | T_1016;
  assign T_2652 = pageReplEn & T_2651;
  assign T_2654 = T_2652 != GEN_581;
  assign T_2655 = T_711 | T_1021;
  assign T_2656 = pageReplEn & T_2655;
  assign T_2658 = T_2656 != GEN_581;
  assign T_2659 = T_716 | T_1026;
  assign T_2660 = pageReplEn & T_2659;
  assign T_2662 = T_2660 != GEN_581;
  assign T_2663 = T_721 | T_1031;
  assign T_2664 = pageReplEn & T_2663;
  assign T_2666 = T_2664 != GEN_581;
  assign T_2667 = T_726 | T_1036;
  assign T_2668 = pageReplEn & T_2667;
  assign T_2670 = T_2668 != GEN_581;
  assign T_2671 = T_731 | T_1041;
  assign T_2672 = pageReplEn & T_2671;
  assign T_2674 = T_2672 != GEN_581;
  assign T_2675 = T_736 | T_1046;
  assign T_2676 = pageReplEn & T_2675;
  assign T_2678 = T_2676 != GEN_581;
  assign T_2679 = T_741 | T_1051;
  assign T_2680 = pageReplEn & T_2679;
  assign T_2682 = T_2680 != GEN_581;
  assign T_2683 = T_746 | T_1056;
  assign T_2684 = pageReplEn & T_2683;
  assign T_2686 = T_2684 != GEN_581;
  assign T_2687 = T_751 | T_1061;
  assign T_2688 = pageReplEn & T_2687;
  assign T_2690 = T_2688 != GEN_581;
  assign T_2691 = T_756 | T_1066;
  assign T_2692 = pageReplEn & T_2691;
  assign T_2694 = T_2692 != GEN_581;
  assign T_2695 = T_761 | T_1071;
  assign T_2696 = pageReplEn & T_2695;
  assign T_2698 = T_2696 != GEN_581;
  assign T_2699 = T_766 | T_1076;
  assign T_2700 = pageReplEn & T_2699;
  assign T_2702 = T_2700 != GEN_581;
  assign T_2703 = T_771 | T_1081;
  assign T_2704 = pageReplEn & T_2703;
  assign T_2706 = T_2704 != GEN_581;
  assign T_2707 = T_776 | T_1086;
  assign T_2708 = pageReplEn & T_2707;
  assign T_2710 = T_2708 != GEN_581;
  assign T_2711 = T_781 | T_1091;
  assign T_2712 = pageReplEn & T_2711;
  assign T_2714 = T_2712 != GEN_581;
  assign T_2715 = T_786 | T_1096;
  assign T_2716 = pageReplEn & T_2715;
  assign T_2718 = T_2716 != GEN_581;
  assign T_2719 = T_791 | T_1101;
  assign T_2720 = pageReplEn & T_2719;
  assign T_2722 = T_2720 != GEN_581;
  assign T_2723 = T_796 | T_1106;
  assign T_2724 = pageReplEn & T_2723;
  assign T_2726 = T_2724 != GEN_581;
  assign T_2727 = T_801 | T_1111;
  assign T_2728 = pageReplEn & T_2727;
  assign T_2730 = T_2728 != GEN_581;
  assign T_2731 = T_806 | T_1116;
  assign T_2732 = pageReplEn & T_2731;
  assign T_2734 = T_2732 != GEN_581;
  assign T_2735 = T_811 | T_1121;
  assign T_2736 = pageReplEn & T_2735;
  assign T_2738 = T_2736 != GEN_581;
  assign T_2739 = T_816 | T_1126;
  assign T_2740 = pageReplEn & T_2739;
  assign T_2742 = T_2740 != GEN_581;
  assign T_2743 = T_821 | T_1131;
  assign T_2744 = pageReplEn & T_2743;
  assign T_2746 = T_2744 != GEN_581;
  assign T_2747 = T_826 | T_1136;
  assign T_2748 = pageReplEn & T_2747;
  assign T_2750 = T_2748 != GEN_581;
  assign T_2751 = T_831 | T_1141;
  assign T_2752 = pageReplEn & T_2751;
  assign T_2754 = T_2752 != GEN_581;
  assign T_2755 = T_836 | T_1146;
  assign T_2756 = pageReplEn & T_2755;
  assign T_2758 = T_2756 != GEN_581;
  assign T_2759 = T_841 | T_1151;
  assign T_2760 = pageReplEn & T_2759;
  assign T_2762 = T_2760 != GEN_581;
  assign T_2763 = T_846 | T_1156;
  assign T_2764 = pageReplEn & T_2763;
  assign T_2766 = T_2764 != GEN_581;
  assign T_2767 = T_851 | T_1161;
  assign T_2768 = pageReplEn & T_2767;
  assign T_2770 = T_2768 != GEN_581;
  assign T_2771 = T_856 | T_1166;
  assign T_2772 = pageReplEn & T_2771;
  assign T_2774 = T_2772 != GEN_581;
  assign T_2775 = T_861 | T_1171;
  assign T_2776 = pageReplEn & T_2775;
  assign T_2778 = T_2776 != GEN_581;
  assign T_2779 = T_866 | T_1176;
  assign T_2780 = pageReplEn & T_2779;
  assign T_2782 = T_2780 != GEN_581;
  assign T_2783 = T_871 | T_1181;
  assign T_2784 = pageReplEn & T_2783;
  assign T_2786 = T_2784 != GEN_581;
  assign T_2787 = T_876 | T_1186;
  assign T_2788 = pageReplEn & T_2787;
  assign T_2790 = T_2788 != GEN_581;
  assign T_2791 = T_881 | T_1191;
  assign T_2792 = pageReplEn & T_2791;
  assign T_2794 = T_2792 != GEN_581;
  assign T_2795 = T_886 | T_1196;
  assign T_2796 = pageReplEn & T_2795;
  assign T_2798 = T_2796 != GEN_581;
  assign T_2804_0 = T_2554;
  assign T_2804_1 = T_2558;
  assign T_2804_2 = T_2562;
  assign T_2804_3 = T_2566;
  assign T_2804_4 = T_2570;
  assign T_2804_5 = T_2574;
  assign T_2804_6 = T_2578;
  assign T_2804_7 = T_2582;
  assign T_2804_8 = T_2586;
  assign T_2804_9 = T_2590;
  assign T_2804_10 = T_2594;
  assign T_2804_11 = T_2598;
  assign T_2804_12 = T_2602;
  assign T_2804_13 = T_2606;
  assign T_2804_14 = T_2610;
  assign T_2804_15 = T_2614;
  assign T_2804_16 = T_2618;
  assign T_2804_17 = T_2622;
  assign T_2804_18 = T_2626;
  assign T_2804_19 = T_2630;
  assign T_2804_20 = T_2634;
  assign T_2804_21 = T_2638;
  assign T_2804_22 = T_2642;
  assign T_2804_23 = T_2646;
  assign T_2804_24 = T_2650;
  assign T_2804_25 = T_2654;
  assign T_2804_26 = T_2658;
  assign T_2804_27 = T_2662;
  assign T_2804_28 = T_2666;
  assign T_2804_29 = T_2670;
  assign T_2804_30 = T_2674;
  assign T_2804_31 = T_2678;
  assign T_2804_32 = T_2682;
  assign T_2804_33 = T_2686;
  assign T_2804_34 = T_2690;
  assign T_2804_35 = T_2694;
  assign T_2804_36 = T_2698;
  assign T_2804_37 = T_2702;
  assign T_2804_38 = T_2706;
  assign T_2804_39 = T_2710;
  assign T_2804_40 = T_2714;
  assign T_2804_41 = T_2718;
  assign T_2804_42 = T_2722;
  assign T_2804_43 = T_2726;
  assign T_2804_44 = T_2730;
  assign T_2804_45 = T_2734;
  assign T_2804_46 = T_2738;
  assign T_2804_47 = T_2742;
  assign T_2804_48 = T_2746;
  assign T_2804_49 = T_2750;
  assign T_2804_50 = T_2754;
  assign T_2804_51 = T_2758;
  assign T_2804_52 = T_2762;
  assign T_2804_53 = T_2766;
  assign T_2804_54 = T_2770;
  assign T_2804_55 = T_2774;
  assign T_2804_56 = T_2778;
  assign T_2804_57 = T_2782;
  assign T_2804_58 = T_2786;
  assign T_2804_59 = T_2790;
  assign T_2804_60 = T_2794;
  assign T_2804_61 = T_2798;
  assign T_2806 = {T_2804_2,T_2804_1};
  assign T_2807 = {T_2806,T_2804_0};
  assign T_2808 = {T_2804_4,T_2804_3};
  assign T_2809 = {T_2804_6,T_2804_5};
  assign T_2810 = {T_2809,T_2808};
  assign T_2811 = {T_2810,T_2807};
  assign T_2812 = {T_2804_8,T_2804_7};
  assign T_2813 = {T_2804_10,T_2804_9};
  assign T_2814 = {T_2813,T_2812};
  assign T_2815 = {T_2804_12,T_2804_11};
  assign T_2816 = {T_2804_14,T_2804_13};
  assign T_2817 = {T_2816,T_2815};
  assign T_2818 = {T_2817,T_2814};
  assign T_2819 = {T_2818,T_2811};
  assign T_2820 = {T_2804_16,T_2804_15};
  assign T_2821 = {T_2804_18,T_2804_17};
  assign T_2822 = {T_2821,T_2820};
  assign T_2823 = {T_2804_20,T_2804_19};
  assign T_2824 = {T_2804_22,T_2804_21};
  assign T_2825 = {T_2824,T_2823};
  assign T_2826 = {T_2825,T_2822};
  assign T_2827 = {T_2804_24,T_2804_23};
  assign T_2828 = {T_2804_26,T_2804_25};
  assign T_2829 = {T_2828,T_2827};
  assign T_2830 = {T_2804_28,T_2804_27};
  assign T_2831 = {T_2804_30,T_2804_29};
  assign T_2832 = {T_2831,T_2830};
  assign T_2833 = {T_2832,T_2829};
  assign T_2834 = {T_2833,T_2826};
  assign T_2835 = {T_2834,T_2819};
  assign T_2836 = {T_2804_33,T_2804_32};
  assign T_2837 = {T_2836,T_2804_31};
  assign T_2838 = {T_2804_35,T_2804_34};
  assign T_2839 = {T_2804_37,T_2804_36};
  assign T_2840 = {T_2839,T_2838};
  assign T_2841 = {T_2840,T_2837};
  assign T_2842 = {T_2804_39,T_2804_38};
  assign T_2843 = {T_2804_41,T_2804_40};
  assign T_2844 = {T_2843,T_2842};
  assign T_2845 = {T_2804_43,T_2804_42};
  assign T_2846 = {T_2804_45,T_2804_44};
  assign T_2847 = {T_2846,T_2845};
  assign T_2848 = {T_2847,T_2844};
  assign T_2849 = {T_2848,T_2841};
  assign T_2850 = {T_2804_47,T_2804_46};
  assign T_2851 = {T_2804_49,T_2804_48};
  assign T_2852 = {T_2851,T_2850};
  assign T_2853 = {T_2804_51,T_2804_50};
  assign T_2854 = {T_2804_53,T_2804_52};
  assign T_2855 = {T_2854,T_2853};
  assign T_2856 = {T_2855,T_2852};
  assign T_2857 = {T_2804_55,T_2804_54};
  assign T_2858 = {T_2804_57,T_2804_56};
  assign T_2859 = {T_2858,T_2857};
  assign T_2860 = {T_2804_59,T_2804_58};
  assign T_2861 = {T_2804_61,T_2804_60};
  assign T_2862 = {T_2861,T_2860};
  assign T_2863 = {T_2862,T_2859};
  assign T_2864 = {T_2863,T_2856};
  assign T_2865 = {T_2864,T_2849};
  assign T_2866 = {T_2865,T_2835};
  assign GEN_780 = {{63'd0}, 1'h1};
  assign T_2868 = GEN_780 << T_2550;
  assign T_2869 = ~ T_2866;
  assign T_2870 = idxValid & T_2869;
  assign GEN_781 = {{2'd0}, T_2870};
  assign T_2871 = GEN_781 | T_2868;
  assign GEN_0 = r_btb_update_bits_isReturn;
  assign GEN_22 = GEN_581 == T_2550 ? GEN_0 : useRAS_0;
  assign GEN_23 = GEN_705 == T_2550 ? GEN_0 : useRAS_1;
  assign GEN_784 = {{4'd0}, 2'h2};
  assign GEN_24 = GEN_784 == T_2550 ? GEN_0 : useRAS_2;
  assign GEN_785 = {{4'd0}, 2'h3};
  assign GEN_25 = GEN_785 == T_2550 ? GEN_0 : useRAS_3;
  assign GEN_786 = {{3'd0}, 3'h4};
  assign GEN_26 = GEN_786 == T_2550 ? GEN_0 : useRAS_4;
  assign GEN_787 = {{3'd0}, 3'h5};
  assign GEN_27 = GEN_787 == T_2550 ? GEN_0 : useRAS_5;
  assign GEN_788 = {{3'd0}, 3'h6};
  assign GEN_28 = GEN_788 == T_2550 ? GEN_0 : useRAS_6;
  assign GEN_789 = {{3'd0}, 3'h7};
  assign GEN_29 = GEN_789 == T_2550 ? GEN_0 : useRAS_7;
  assign GEN_790 = {{2'd0}, 4'h8};
  assign GEN_30 = GEN_790 == T_2550 ? GEN_0 : useRAS_8;
  assign GEN_791 = {{2'd0}, 4'h9};
  assign GEN_31 = GEN_791 == T_2550 ? GEN_0 : useRAS_9;
  assign GEN_792 = {{2'd0}, 4'ha};
  assign GEN_32 = GEN_792 == T_2550 ? GEN_0 : useRAS_10;
  assign GEN_793 = {{2'd0}, 4'hb};
  assign GEN_33 = GEN_793 == T_2550 ? GEN_0 : useRAS_11;
  assign GEN_794 = {{2'd0}, 4'hc};
  assign GEN_34 = GEN_794 == T_2550 ? GEN_0 : useRAS_12;
  assign GEN_795 = {{2'd0}, 4'hd};
  assign GEN_35 = GEN_795 == T_2550 ? GEN_0 : useRAS_13;
  assign GEN_796 = {{2'd0}, 4'he};
  assign GEN_36 = GEN_796 == T_2550 ? GEN_0 : useRAS_14;
  assign GEN_797 = {{2'd0}, 4'hf};
  assign GEN_37 = GEN_797 == T_2550 ? GEN_0 : useRAS_15;
  assign GEN_798 = {{1'd0}, 5'h10};
  assign GEN_38 = GEN_798 == T_2550 ? GEN_0 : useRAS_16;
  assign GEN_799 = {{1'd0}, 5'h11};
  assign GEN_39 = GEN_799 == T_2550 ? GEN_0 : useRAS_17;
  assign GEN_800 = {{1'd0}, 5'h12};
  assign GEN_40 = GEN_800 == T_2550 ? GEN_0 : useRAS_18;
  assign GEN_801 = {{1'd0}, 5'h13};
  assign GEN_41 = GEN_801 == T_2550 ? GEN_0 : useRAS_19;
  assign GEN_802 = {{1'd0}, 5'h14};
  assign GEN_42 = GEN_802 == T_2550 ? GEN_0 : useRAS_20;
  assign GEN_803 = {{1'd0}, 5'h15};
  assign GEN_43 = GEN_803 == T_2550 ? GEN_0 : useRAS_21;
  assign GEN_804 = {{1'd0}, 5'h16};
  assign GEN_44 = GEN_804 == T_2550 ? GEN_0 : useRAS_22;
  assign GEN_805 = {{1'd0}, 5'h17};
  assign GEN_45 = GEN_805 == T_2550 ? GEN_0 : useRAS_23;
  assign GEN_806 = {{1'd0}, 5'h18};
  assign GEN_46 = GEN_806 == T_2550 ? GEN_0 : useRAS_24;
  assign GEN_807 = {{1'd0}, 5'h19};
  assign GEN_47 = GEN_807 == T_2550 ? GEN_0 : useRAS_25;
  assign GEN_808 = {{1'd0}, 5'h1a};
  assign GEN_48 = GEN_808 == T_2550 ? GEN_0 : useRAS_26;
  assign GEN_809 = {{1'd0}, 5'h1b};
  assign GEN_49 = GEN_809 == T_2550 ? GEN_0 : useRAS_27;
  assign GEN_810 = {{1'd0}, 5'h1c};
  assign GEN_50 = GEN_810 == T_2550 ? GEN_0 : useRAS_28;
  assign GEN_811 = {{1'd0}, 5'h1d};
  assign GEN_51 = GEN_811 == T_2550 ? GEN_0 : useRAS_29;
  assign GEN_812 = {{1'd0}, 5'h1e};
  assign GEN_52 = GEN_812 == T_2550 ? GEN_0 : useRAS_30;
  assign GEN_813 = {{1'd0}, 5'h1f};
  assign GEN_53 = GEN_813 == T_2550 ? GEN_0 : useRAS_31;
  assign GEN_54 = 6'h20 == T_2550 ? GEN_0 : useRAS_32;
  assign GEN_55 = 6'h21 == T_2550 ? GEN_0 : useRAS_33;
  assign GEN_56 = 6'h22 == T_2550 ? GEN_0 : useRAS_34;
  assign GEN_57 = 6'h23 == T_2550 ? GEN_0 : useRAS_35;
  assign GEN_58 = 6'h24 == T_2550 ? GEN_0 : useRAS_36;
  assign GEN_59 = 6'h25 == T_2550 ? GEN_0 : useRAS_37;
  assign GEN_60 = 6'h26 == T_2550 ? GEN_0 : useRAS_38;
  assign GEN_61 = 6'h27 == T_2550 ? GEN_0 : useRAS_39;
  assign GEN_62 = 6'h28 == T_2550 ? GEN_0 : useRAS_40;
  assign GEN_63 = 6'h29 == T_2550 ? GEN_0 : useRAS_41;
  assign GEN_64 = 6'h2a == T_2550 ? GEN_0 : useRAS_42;
  assign GEN_65 = 6'h2b == T_2550 ? GEN_0 : useRAS_43;
  assign GEN_66 = 6'h2c == T_2550 ? GEN_0 : useRAS_44;
  assign GEN_67 = 6'h2d == T_2550 ? GEN_0 : useRAS_45;
  assign GEN_68 = 6'h2e == T_2550 ? GEN_0 : useRAS_46;
  assign GEN_69 = 6'h2f == T_2550 ? GEN_0 : useRAS_47;
  assign GEN_70 = 6'h30 == T_2550 ? GEN_0 : useRAS_48;
  assign GEN_71 = 6'h31 == T_2550 ? GEN_0 : useRAS_49;
  assign GEN_72 = 6'h32 == T_2550 ? GEN_0 : useRAS_50;
  assign GEN_73 = 6'h33 == T_2550 ? GEN_0 : useRAS_51;
  assign GEN_74 = 6'h34 == T_2550 ? GEN_0 : useRAS_52;
  assign GEN_75 = 6'h35 == T_2550 ? GEN_0 : useRAS_53;
  assign GEN_76 = 6'h36 == T_2550 ? GEN_0 : useRAS_54;
  assign GEN_77 = 6'h37 == T_2550 ? GEN_0 : useRAS_55;
  assign GEN_78 = 6'h38 == T_2550 ? GEN_0 : useRAS_56;
  assign GEN_79 = 6'h39 == T_2550 ? GEN_0 : useRAS_57;
  assign GEN_80 = 6'h3a == T_2550 ? GEN_0 : useRAS_58;
  assign GEN_81 = 6'h3b == T_2550 ? GEN_0 : useRAS_59;
  assign GEN_82 = 6'h3c == T_2550 ? GEN_0 : useRAS_60;
  assign GEN_83 = 6'h3d == T_2550 ? GEN_0 : useRAS_61;
  assign GEN_1 = r_btb_update_bits_isJump;
  assign GEN_84 = GEN_581 == T_2550 ? GEN_1 : isJump_0;
  assign GEN_85 = GEN_705 == T_2550 ? GEN_1 : isJump_1;
  assign GEN_86 = GEN_784 == T_2550 ? GEN_1 : isJump_2;
  assign GEN_87 = GEN_785 == T_2550 ? GEN_1 : isJump_3;
  assign GEN_88 = GEN_786 == T_2550 ? GEN_1 : isJump_4;
  assign GEN_89 = GEN_787 == T_2550 ? GEN_1 : isJump_5;
  assign GEN_90 = GEN_788 == T_2550 ? GEN_1 : isJump_6;
  assign GEN_91 = GEN_789 == T_2550 ? GEN_1 : isJump_7;
  assign GEN_92 = GEN_790 == T_2550 ? GEN_1 : isJump_8;
  assign GEN_93 = GEN_791 == T_2550 ? GEN_1 : isJump_9;
  assign GEN_94 = GEN_792 == T_2550 ? GEN_1 : isJump_10;
  assign GEN_95 = GEN_793 == T_2550 ? GEN_1 : isJump_11;
  assign GEN_96 = GEN_794 == T_2550 ? GEN_1 : isJump_12;
  assign GEN_97 = GEN_795 == T_2550 ? GEN_1 : isJump_13;
  assign GEN_98 = GEN_796 == T_2550 ? GEN_1 : isJump_14;
  assign GEN_99 = GEN_797 == T_2550 ? GEN_1 : isJump_15;
  assign GEN_100 = GEN_798 == T_2550 ? GEN_1 : isJump_16;
  assign GEN_101 = GEN_799 == T_2550 ? GEN_1 : isJump_17;
  assign GEN_102 = GEN_800 == T_2550 ? GEN_1 : isJump_18;
  assign GEN_103 = GEN_801 == T_2550 ? GEN_1 : isJump_19;
  assign GEN_104 = GEN_802 == T_2550 ? GEN_1 : isJump_20;
  assign GEN_105 = GEN_803 == T_2550 ? GEN_1 : isJump_21;
  assign GEN_106 = GEN_804 == T_2550 ? GEN_1 : isJump_22;
  assign GEN_107 = GEN_805 == T_2550 ? GEN_1 : isJump_23;
  assign GEN_108 = GEN_806 == T_2550 ? GEN_1 : isJump_24;
  assign GEN_109 = GEN_807 == T_2550 ? GEN_1 : isJump_25;
  assign GEN_110 = GEN_808 == T_2550 ? GEN_1 : isJump_26;
  assign GEN_111 = GEN_809 == T_2550 ? GEN_1 : isJump_27;
  assign GEN_112 = GEN_810 == T_2550 ? GEN_1 : isJump_28;
  assign GEN_113 = GEN_811 == T_2550 ? GEN_1 : isJump_29;
  assign GEN_114 = GEN_812 == T_2550 ? GEN_1 : isJump_30;
  assign GEN_115 = GEN_813 == T_2550 ? GEN_1 : isJump_31;
  assign GEN_116 = 6'h20 == T_2550 ? GEN_1 : isJump_32;
  assign GEN_117 = 6'h21 == T_2550 ? GEN_1 : isJump_33;
  assign GEN_118 = 6'h22 == T_2550 ? GEN_1 : isJump_34;
  assign GEN_119 = 6'h23 == T_2550 ? GEN_1 : isJump_35;
  assign GEN_120 = 6'h24 == T_2550 ? GEN_1 : isJump_36;
  assign GEN_121 = 6'h25 == T_2550 ? GEN_1 : isJump_37;
  assign GEN_122 = 6'h26 == T_2550 ? GEN_1 : isJump_38;
  assign GEN_123 = 6'h27 == T_2550 ? GEN_1 : isJump_39;
  assign GEN_124 = 6'h28 == T_2550 ? GEN_1 : isJump_40;
  assign GEN_125 = 6'h29 == T_2550 ? GEN_1 : isJump_41;
  assign GEN_126 = 6'h2a == T_2550 ? GEN_1 : isJump_42;
  assign GEN_127 = 6'h2b == T_2550 ? GEN_1 : isJump_43;
  assign GEN_128 = 6'h2c == T_2550 ? GEN_1 : isJump_44;
  assign GEN_129 = 6'h2d == T_2550 ? GEN_1 : isJump_45;
  assign GEN_130 = 6'h2e == T_2550 ? GEN_1 : isJump_46;
  assign GEN_131 = 6'h2f == T_2550 ? GEN_1 : isJump_47;
  assign GEN_132 = 6'h30 == T_2550 ? GEN_1 : isJump_48;
  assign GEN_133 = 6'h31 == T_2550 ? GEN_1 : isJump_49;
  assign GEN_134 = 6'h32 == T_2550 ? GEN_1 : isJump_50;
  assign GEN_135 = 6'h33 == T_2550 ? GEN_1 : isJump_51;
  assign GEN_136 = 6'h34 == T_2550 ? GEN_1 : isJump_52;
  assign GEN_137 = 6'h35 == T_2550 ? GEN_1 : isJump_53;
  assign GEN_138 = 6'h36 == T_2550 ? GEN_1 : isJump_54;
  assign GEN_139 = 6'h37 == T_2550 ? GEN_1 : isJump_55;
  assign GEN_140 = 6'h38 == T_2550 ? GEN_1 : isJump_56;
  assign GEN_141 = 6'h39 == T_2550 ? GEN_1 : isJump_57;
  assign GEN_142 = 6'h3a == T_2550 ? GEN_1 : isJump_58;
  assign GEN_143 = 6'h3b == T_2550 ? GEN_1 : isJump_59;
  assign GEN_144 = 6'h3c == T_2550 ? GEN_1 : isJump_60;
  assign GEN_145 = 6'h3d == T_2550 ? GEN_1 : isJump_61;
  assign T_2881 = idxPageUpdateOH & 6'h15;
  assign T_2883 = T_2881 != GEN_581;
  assign T_2884 = T_2883 ? doIdxPageRepl : doTgtPageRepl;
  assign T_2887 = T_2883 ? T_1939 : T_1398;
  assign T_2888 = pageReplEn[0];
  assign T_2889 = T_2884 & T_2888;
  assign T_2892 = pageReplEn[2];
  assign T_2893 = T_2884 & T_2892;
  assign T_2896 = pageReplEn[4];
  assign T_2897 = T_2884 & T_2896;
  assign T_2900 = T_2883 ? doTgtPageRepl : doIdxPageRepl;
  assign T_2903 = T_2883 ? T_1398 : T_1939;
  assign T_2904 = pageReplEn[1];
  assign T_2905 = T_2900 & T_2904;
  assign T_2908 = pageReplEn[3];
  assign T_2909 = T_2900 & T_2908;
  assign T_2912 = pageReplEn[5];
  assign T_2913 = T_2900 & T_2912;
  assign T_2916 = pageValid | pageReplEn;
  assign GEN_176 = doPageRepl ? T_2916 : pageValid;
  assign GEN_239 = r_btb_update_valid ? T_2871 : {{2'd0}, idxValid};
  assign GEN_261 = r_btb_update_valid ? GEN_22 : useRAS_0;
  assign GEN_262 = r_btb_update_valid ? GEN_23 : useRAS_1;
  assign GEN_263 = r_btb_update_valid ? GEN_24 : useRAS_2;
  assign GEN_264 = r_btb_update_valid ? GEN_25 : useRAS_3;
  assign GEN_265 = r_btb_update_valid ? GEN_26 : useRAS_4;
  assign GEN_266 = r_btb_update_valid ? GEN_27 : useRAS_5;
  assign GEN_267 = r_btb_update_valid ? GEN_28 : useRAS_6;
  assign GEN_268 = r_btb_update_valid ? GEN_29 : useRAS_7;
  assign GEN_269 = r_btb_update_valid ? GEN_30 : useRAS_8;
  assign GEN_270 = r_btb_update_valid ? GEN_31 : useRAS_9;
  assign GEN_271 = r_btb_update_valid ? GEN_32 : useRAS_10;
  assign GEN_272 = r_btb_update_valid ? GEN_33 : useRAS_11;
  assign GEN_273 = r_btb_update_valid ? GEN_34 : useRAS_12;
  assign GEN_274 = r_btb_update_valid ? GEN_35 : useRAS_13;
  assign GEN_275 = r_btb_update_valid ? GEN_36 : useRAS_14;
  assign GEN_276 = r_btb_update_valid ? GEN_37 : useRAS_15;
  assign GEN_277 = r_btb_update_valid ? GEN_38 : useRAS_16;
  assign GEN_278 = r_btb_update_valid ? GEN_39 : useRAS_17;
  assign GEN_279 = r_btb_update_valid ? GEN_40 : useRAS_18;
  assign GEN_280 = r_btb_update_valid ? GEN_41 : useRAS_19;
  assign GEN_281 = r_btb_update_valid ? GEN_42 : useRAS_20;
  assign GEN_282 = r_btb_update_valid ? GEN_43 : useRAS_21;
  assign GEN_283 = r_btb_update_valid ? GEN_44 : useRAS_22;
  assign GEN_284 = r_btb_update_valid ? GEN_45 : useRAS_23;
  assign GEN_285 = r_btb_update_valid ? GEN_46 : useRAS_24;
  assign GEN_286 = r_btb_update_valid ? GEN_47 : useRAS_25;
  assign GEN_287 = r_btb_update_valid ? GEN_48 : useRAS_26;
  assign GEN_288 = r_btb_update_valid ? GEN_49 : useRAS_27;
  assign GEN_289 = r_btb_update_valid ? GEN_50 : useRAS_28;
  assign GEN_290 = r_btb_update_valid ? GEN_51 : useRAS_29;
  assign GEN_291 = r_btb_update_valid ? GEN_52 : useRAS_30;
  assign GEN_292 = r_btb_update_valid ? GEN_53 : useRAS_31;
  assign GEN_293 = r_btb_update_valid ? GEN_54 : useRAS_32;
  assign GEN_294 = r_btb_update_valid ? GEN_55 : useRAS_33;
  assign GEN_295 = r_btb_update_valid ? GEN_56 : useRAS_34;
  assign GEN_296 = r_btb_update_valid ? GEN_57 : useRAS_35;
  assign GEN_297 = r_btb_update_valid ? GEN_58 : useRAS_36;
  assign GEN_298 = r_btb_update_valid ? GEN_59 : useRAS_37;
  assign GEN_299 = r_btb_update_valid ? GEN_60 : useRAS_38;
  assign GEN_300 = r_btb_update_valid ? GEN_61 : useRAS_39;
  assign GEN_301 = r_btb_update_valid ? GEN_62 : useRAS_40;
  assign GEN_302 = r_btb_update_valid ? GEN_63 : useRAS_41;
  assign GEN_303 = r_btb_update_valid ? GEN_64 : useRAS_42;
  assign GEN_304 = r_btb_update_valid ? GEN_65 : useRAS_43;
  assign GEN_305 = r_btb_update_valid ? GEN_66 : useRAS_44;
  assign GEN_306 = r_btb_update_valid ? GEN_67 : useRAS_45;
  assign GEN_307 = r_btb_update_valid ? GEN_68 : useRAS_46;
  assign GEN_308 = r_btb_update_valid ? GEN_69 : useRAS_47;
  assign GEN_309 = r_btb_update_valid ? GEN_70 : useRAS_48;
  assign GEN_310 = r_btb_update_valid ? GEN_71 : useRAS_49;
  assign GEN_311 = r_btb_update_valid ? GEN_72 : useRAS_50;
  assign GEN_312 = r_btb_update_valid ? GEN_73 : useRAS_51;
  assign GEN_313 = r_btb_update_valid ? GEN_74 : useRAS_52;
  assign GEN_314 = r_btb_update_valid ? GEN_75 : useRAS_53;
  assign GEN_315 = r_btb_update_valid ? GEN_76 : useRAS_54;
  assign GEN_316 = r_btb_update_valid ? GEN_77 : useRAS_55;
  assign GEN_317 = r_btb_update_valid ? GEN_78 : useRAS_56;
  assign GEN_318 = r_btb_update_valid ? GEN_79 : useRAS_57;
  assign GEN_319 = r_btb_update_valid ? GEN_80 : useRAS_58;
  assign GEN_320 = r_btb_update_valid ? GEN_81 : useRAS_59;
  assign GEN_321 = r_btb_update_valid ? GEN_82 : useRAS_60;
  assign GEN_322 = r_btb_update_valid ? GEN_83 : useRAS_61;
  assign GEN_324 = r_btb_update_valid ? GEN_84 : isJump_0;
  assign GEN_325 = r_btb_update_valid ? GEN_85 : isJump_1;
  assign GEN_326 = r_btb_update_valid ? GEN_86 : isJump_2;
  assign GEN_327 = r_btb_update_valid ? GEN_87 : isJump_3;
  assign GEN_328 = r_btb_update_valid ? GEN_88 : isJump_4;
  assign GEN_329 = r_btb_update_valid ? GEN_89 : isJump_5;
  assign GEN_330 = r_btb_update_valid ? GEN_90 : isJump_6;
  assign GEN_331 = r_btb_update_valid ? GEN_91 : isJump_7;
  assign GEN_332 = r_btb_update_valid ? GEN_92 : isJump_8;
  assign GEN_333 = r_btb_update_valid ? GEN_93 : isJump_9;
  assign GEN_334 = r_btb_update_valid ? GEN_94 : isJump_10;
  assign GEN_335 = r_btb_update_valid ? GEN_95 : isJump_11;
  assign GEN_336 = r_btb_update_valid ? GEN_96 : isJump_12;
  assign GEN_337 = r_btb_update_valid ? GEN_97 : isJump_13;
  assign GEN_338 = r_btb_update_valid ? GEN_98 : isJump_14;
  assign GEN_339 = r_btb_update_valid ? GEN_99 : isJump_15;
  assign GEN_340 = r_btb_update_valid ? GEN_100 : isJump_16;
  assign GEN_341 = r_btb_update_valid ? GEN_101 : isJump_17;
  assign GEN_342 = r_btb_update_valid ? GEN_102 : isJump_18;
  assign GEN_343 = r_btb_update_valid ? GEN_103 : isJump_19;
  assign GEN_344 = r_btb_update_valid ? GEN_104 : isJump_20;
  assign GEN_345 = r_btb_update_valid ? GEN_105 : isJump_21;
  assign GEN_346 = r_btb_update_valid ? GEN_106 : isJump_22;
  assign GEN_347 = r_btb_update_valid ? GEN_107 : isJump_23;
  assign GEN_348 = r_btb_update_valid ? GEN_108 : isJump_24;
  assign GEN_349 = r_btb_update_valid ? GEN_109 : isJump_25;
  assign GEN_350 = r_btb_update_valid ? GEN_110 : isJump_26;
  assign GEN_351 = r_btb_update_valid ? GEN_111 : isJump_27;
  assign GEN_352 = r_btb_update_valid ? GEN_112 : isJump_28;
  assign GEN_353 = r_btb_update_valid ? GEN_113 : isJump_29;
  assign GEN_354 = r_btb_update_valid ? GEN_114 : isJump_30;
  assign GEN_355 = r_btb_update_valid ? GEN_115 : isJump_31;
  assign GEN_356 = r_btb_update_valid ? GEN_116 : isJump_32;
  assign GEN_357 = r_btb_update_valid ? GEN_117 : isJump_33;
  assign GEN_358 = r_btb_update_valid ? GEN_118 : isJump_34;
  assign GEN_359 = r_btb_update_valid ? GEN_119 : isJump_35;
  assign GEN_360 = r_btb_update_valid ? GEN_120 : isJump_36;
  assign GEN_361 = r_btb_update_valid ? GEN_121 : isJump_37;
  assign GEN_362 = r_btb_update_valid ? GEN_122 : isJump_38;
  assign GEN_363 = r_btb_update_valid ? GEN_123 : isJump_39;
  assign GEN_364 = r_btb_update_valid ? GEN_124 : isJump_40;
  assign GEN_365 = r_btb_update_valid ? GEN_125 : isJump_41;
  assign GEN_366 = r_btb_update_valid ? GEN_126 : isJump_42;
  assign GEN_367 = r_btb_update_valid ? GEN_127 : isJump_43;
  assign GEN_368 = r_btb_update_valid ? GEN_128 : isJump_44;
  assign GEN_369 = r_btb_update_valid ? GEN_129 : isJump_45;
  assign GEN_370 = r_btb_update_valid ? GEN_130 : isJump_46;
  assign GEN_371 = r_btb_update_valid ? GEN_131 : isJump_47;
  assign GEN_372 = r_btb_update_valid ? GEN_132 : isJump_48;
  assign GEN_373 = r_btb_update_valid ? GEN_133 : isJump_49;
  assign GEN_374 = r_btb_update_valid ? GEN_134 : isJump_50;
  assign GEN_375 = r_btb_update_valid ? GEN_135 : isJump_51;
  assign GEN_376 = r_btb_update_valid ? GEN_136 : isJump_52;
  assign GEN_377 = r_btb_update_valid ? GEN_137 : isJump_53;
  assign GEN_378 = r_btb_update_valid ? GEN_138 : isJump_54;
  assign GEN_379 = r_btb_update_valid ? GEN_139 : isJump_55;
  assign GEN_380 = r_btb_update_valid ? GEN_140 : isJump_56;
  assign GEN_381 = r_btb_update_valid ? GEN_141 : isJump_57;
  assign GEN_382 = r_btb_update_valid ? GEN_142 : isJump_58;
  assign GEN_383 = r_btb_update_valid ? GEN_143 : isJump_59;
  assign GEN_384 = r_btb_update_valid ? GEN_144 : isJump_60;
  assign GEN_385 = r_btb_update_valid ? GEN_145 : isJump_61;
  assign GEN_393 = r_btb_update_valid ? T_2889 : 1'h0;
  assign GEN_398 = r_btb_update_valid ? T_2893 : 1'h0;
  assign GEN_403 = r_btb_update_valid ? T_2897 : 1'h0;
  assign GEN_408 = r_btb_update_valid ? T_2905 : 1'h0;
  assign GEN_413 = r_btb_update_valid ? T_2909 : 1'h0;
  assign GEN_418 = r_btb_update_valid ? T_2913 : 1'h0;
  assign GEN_421 = r_btb_update_valid ? GEN_176 : pageValid;
  assign GEN_422 = io_invalidate ? {{63'd0}, 1'h0} : GEN_239;
  assign GEN_423 = io_invalidate ? {{5'd0}, 1'h0} : GEN_421;
  assign GEN_847 = {{61'd0}, 1'h0};
  assign T_2920 = hits != GEN_847;
  assign T_2921 = hits[0];
  assign T_2922 = hits[1];
  assign T_2923 = hits[2];
  assign T_2924 = hits[3];
  assign T_2925 = hits[4];
  assign T_2926 = hits[5];
  assign T_2927 = hits[6];
  assign T_2928 = hits[7];
  assign T_2929 = hits[8];
  assign T_2930 = hits[9];
  assign T_2931 = hits[10];
  assign T_2932 = hits[11];
  assign T_2933 = hits[12];
  assign T_2934 = hits[13];
  assign T_2935 = hits[14];
  assign T_2936 = hits[15];
  assign T_2937 = hits[16];
  assign T_2938 = hits[17];
  assign T_2939 = hits[18];
  assign T_2940 = hits[19];
  assign T_2941 = hits[20];
  assign T_2942 = hits[21];
  assign T_2943 = hits[22];
  assign T_2944 = hits[23];
  assign T_2945 = hits[24];
  assign T_2946 = hits[25];
  assign T_2947 = hits[26];
  assign T_2948 = hits[27];
  assign T_2949 = hits[28];
  assign T_2950 = hits[29];
  assign T_2951 = hits[30];
  assign T_2952 = hits[31];
  assign T_2953 = hits[32];
  assign T_2954 = hits[33];
  assign T_2955 = hits[34];
  assign T_2956 = hits[35];
  assign T_2957 = hits[36];
  assign T_2958 = hits[37];
  assign T_2959 = hits[38];
  assign T_2960 = hits[39];
  assign T_2961 = hits[40];
  assign T_2962 = hits[41];
  assign T_2963 = hits[42];
  assign T_2964 = hits[43];
  assign T_2965 = hits[44];
  assign T_2966 = hits[45];
  assign T_2967 = hits[46];
  assign T_2968 = hits[47];
  assign T_2969 = hits[48];
  assign T_2970 = hits[49];
  assign T_2971 = hits[50];
  assign T_2972 = hits[51];
  assign T_2973 = hits[52];
  assign T_2974 = hits[53];
  assign T_2975 = hits[54];
  assign T_2976 = hits[55];
  assign T_2977 = hits[56];
  assign T_2978 = hits[57];
  assign T_2979 = hits[58];
  assign T_2980 = hits[59];
  assign T_2981 = hits[60];
  assign T_2982 = hits[61];
  assign T_2984 = T_2921 ? T_891 : {{5'd0}, 1'h0};
  assign T_2986 = T_2922 ? T_896 : {{5'd0}, 1'h0};
  assign T_2988 = T_2923 ? T_901 : {{5'd0}, 1'h0};
  assign T_2990 = T_2924 ? T_906 : {{5'd0}, 1'h0};
  assign T_2992 = T_2925 ? T_911 : {{5'd0}, 1'h0};
  assign T_2994 = T_2926 ? T_916 : {{5'd0}, 1'h0};
  assign T_2996 = T_2927 ? T_921 : {{5'd0}, 1'h0};
  assign T_2998 = T_2928 ? T_926 : {{5'd0}, 1'h0};
  assign T_3000 = T_2929 ? T_931 : {{5'd0}, 1'h0};
  assign T_3002 = T_2930 ? T_936 : {{5'd0}, 1'h0};
  assign T_3004 = T_2931 ? T_941 : {{5'd0}, 1'h0};
  assign T_3006 = T_2932 ? T_946 : {{5'd0}, 1'h0};
  assign T_3008 = T_2933 ? T_951 : {{5'd0}, 1'h0};
  assign T_3010 = T_2934 ? T_956 : {{5'd0}, 1'h0};
  assign T_3012 = T_2935 ? T_961 : {{5'd0}, 1'h0};
  assign T_3014 = T_2936 ? T_966 : {{5'd0}, 1'h0};
  assign T_3016 = T_2937 ? T_971 : {{5'd0}, 1'h0};
  assign T_3018 = T_2938 ? T_976 : {{5'd0}, 1'h0};
  assign T_3020 = T_2939 ? T_981 : {{5'd0}, 1'h0};
  assign T_3022 = T_2940 ? T_986 : {{5'd0}, 1'h0};
  assign T_3024 = T_2941 ? T_991 : {{5'd0}, 1'h0};
  assign T_3026 = T_2942 ? T_996 : {{5'd0}, 1'h0};
  assign T_3028 = T_2943 ? T_1001 : {{5'd0}, 1'h0};
  assign T_3030 = T_2944 ? T_1006 : {{5'd0}, 1'h0};
  assign T_3032 = T_2945 ? T_1011 : {{5'd0}, 1'h0};
  assign T_3034 = T_2946 ? T_1016 : {{5'd0}, 1'h0};
  assign T_3036 = T_2947 ? T_1021 : {{5'd0}, 1'h0};
  assign T_3038 = T_2948 ? T_1026 : {{5'd0}, 1'h0};
  assign T_3040 = T_2949 ? T_1031 : {{5'd0}, 1'h0};
  assign T_3042 = T_2950 ? T_1036 : {{5'd0}, 1'h0};
  assign T_3044 = T_2951 ? T_1041 : {{5'd0}, 1'h0};
  assign T_3046 = T_2952 ? T_1046 : {{5'd0}, 1'h0};
  assign T_3048 = T_2953 ? T_1051 : {{5'd0}, 1'h0};
  assign T_3050 = T_2954 ? T_1056 : {{5'd0}, 1'h0};
  assign T_3052 = T_2955 ? T_1061 : {{5'd0}, 1'h0};
  assign T_3054 = T_2956 ? T_1066 : {{5'd0}, 1'h0};
  assign T_3056 = T_2957 ? T_1071 : {{5'd0}, 1'h0};
  assign T_3058 = T_2958 ? T_1076 : {{5'd0}, 1'h0};
  assign T_3060 = T_2959 ? T_1081 : {{5'd0}, 1'h0};
  assign T_3062 = T_2960 ? T_1086 : {{5'd0}, 1'h0};
  assign T_3064 = T_2961 ? T_1091 : {{5'd0}, 1'h0};
  assign T_3066 = T_2962 ? T_1096 : {{5'd0}, 1'h0};
  assign T_3068 = T_2963 ? T_1101 : {{5'd0}, 1'h0};
  assign T_3070 = T_2964 ? T_1106 : {{5'd0}, 1'h0};
  assign T_3072 = T_2965 ? T_1111 : {{5'd0}, 1'h0};
  assign T_3074 = T_2966 ? T_1116 : {{5'd0}, 1'h0};
  assign T_3076 = T_2967 ? T_1121 : {{5'd0}, 1'h0};
  assign T_3078 = T_2968 ? T_1126 : {{5'd0}, 1'h0};
  assign T_3080 = T_2969 ? T_1131 : {{5'd0}, 1'h0};
  assign T_3082 = T_2970 ? T_1136 : {{5'd0}, 1'h0};
  assign T_3084 = T_2971 ? T_1141 : {{5'd0}, 1'h0};
  assign T_3086 = T_2972 ? T_1146 : {{5'd0}, 1'h0};
  assign T_3088 = T_2973 ? T_1151 : {{5'd0}, 1'h0};
  assign T_3090 = T_2974 ? T_1156 : {{5'd0}, 1'h0};
  assign T_3092 = T_2975 ? T_1161 : {{5'd0}, 1'h0};
  assign T_3094 = T_2976 ? T_1166 : {{5'd0}, 1'h0};
  assign T_3096 = T_2977 ? T_1171 : {{5'd0}, 1'h0};
  assign T_3098 = T_2978 ? T_1176 : {{5'd0}, 1'h0};
  assign T_3100 = T_2979 ? T_1181 : {{5'd0}, 1'h0};
  assign T_3102 = T_2980 ? T_1186 : {{5'd0}, 1'h0};
  assign T_3104 = T_2981 ? T_1191 : {{5'd0}, 1'h0};
  assign T_3106 = T_2982 ? T_1196 : {{5'd0}, 1'h0};
  assign T_3108 = T_2984 | T_2986;
  assign T_3109 = T_3108 | T_2988;
  assign T_3110 = T_3109 | T_2990;
  assign T_3111 = T_3110 | T_2992;
  assign T_3112 = T_3111 | T_2994;
  assign T_3113 = T_3112 | T_2996;
  assign T_3114 = T_3113 | T_2998;
  assign T_3115 = T_3114 | T_3000;
  assign T_3116 = T_3115 | T_3002;
  assign T_3117 = T_3116 | T_3004;
  assign T_3118 = T_3117 | T_3006;
  assign T_3119 = T_3118 | T_3008;
  assign T_3120 = T_3119 | T_3010;
  assign T_3121 = T_3120 | T_3012;
  assign T_3122 = T_3121 | T_3014;
  assign T_3123 = T_3122 | T_3016;
  assign T_3124 = T_3123 | T_3018;
  assign T_3125 = T_3124 | T_3020;
  assign T_3126 = T_3125 | T_3022;
  assign T_3127 = T_3126 | T_3024;
  assign T_3128 = T_3127 | T_3026;
  assign T_3129 = T_3128 | T_3028;
  assign T_3130 = T_3129 | T_3030;
  assign T_3131 = T_3130 | T_3032;
  assign T_3132 = T_3131 | T_3034;
  assign T_3133 = T_3132 | T_3036;
  assign T_3134 = T_3133 | T_3038;
  assign T_3135 = T_3134 | T_3040;
  assign T_3136 = T_3135 | T_3042;
  assign T_3137 = T_3136 | T_3044;
  assign T_3138 = T_3137 | T_3046;
  assign T_3139 = T_3138 | T_3048;
  assign T_3140 = T_3139 | T_3050;
  assign T_3141 = T_3140 | T_3052;
  assign T_3142 = T_3141 | T_3054;
  assign T_3143 = T_3142 | T_3056;
  assign T_3144 = T_3143 | T_3058;
  assign T_3145 = T_3144 | T_3060;
  assign T_3146 = T_3145 | T_3062;
  assign T_3147 = T_3146 | T_3064;
  assign T_3148 = T_3147 | T_3066;
  assign T_3149 = T_3148 | T_3068;
  assign T_3150 = T_3149 | T_3070;
  assign T_3151 = T_3150 | T_3072;
  assign T_3152 = T_3151 | T_3074;
  assign T_3153 = T_3152 | T_3076;
  assign T_3154 = T_3153 | T_3078;
  assign T_3155 = T_3154 | T_3080;
  assign T_3156 = T_3155 | T_3082;
  assign T_3157 = T_3156 | T_3084;
  assign T_3158 = T_3157 | T_3086;
  assign T_3159 = T_3158 | T_3088;
  assign T_3160 = T_3159 | T_3090;
  assign T_3161 = T_3160 | T_3092;
  assign T_3162 = T_3161 | T_3094;
  assign T_3163 = T_3162 | T_3096;
  assign T_3164 = T_3163 | T_3098;
  assign T_3165 = T_3164 | T_3100;
  assign T_3166 = T_3165 | T_3102;
  assign T_3167 = T_3166 | T_3104;
  assign T_3168 = T_3167 | T_3106;
  assign T_3169 = T_3168;
  assign T_3170 = T_3169[0];
  assign T_3171 = T_3169[1];
  assign T_3172 = T_3169[2];
  assign T_3173 = T_3169[3];
  assign T_3174 = T_3169[4];
  assign T_3175 = T_3169[5];
  assign T_3189 = T_3170 ? pages_T_3177_data : {{26'd0}, 1'h0};
  assign T_3191 = T_3171 ? pages_T_3179_data : {{26'd0}, 1'h0};
  assign T_3193 = T_3172 ? pages_T_3181_data : {{26'd0}, 1'h0};
  assign T_3195 = T_3173 ? pages_T_3183_data : {{26'd0}, 1'h0};
  assign T_3197 = T_3174 ? pages_T_3185_data : {{26'd0}, 1'h0};
  assign T_3199 = T_3175 ? pages_T_3187_data : {{26'd0}, 1'h0};
  assign T_3201 = T_3189 | T_3191;
  assign T_3202 = T_3201 | T_3193;
  assign T_3203 = T_3202 | T_3195;
  assign T_3204 = T_3203 | T_3197;
  assign T_3205 = T_3204 | T_3199;
  assign T_3206 = T_3205;
  assign T_3394 = T_2921 ? tgts_T_3270_data : {{11'd0}, 1'h0};
  assign T_3396 = T_2922 ? tgts_T_3272_data : {{11'd0}, 1'h0};
  assign T_3398 = T_2923 ? tgts_T_3274_data : {{11'd0}, 1'h0};
  assign T_3400 = T_2924 ? tgts_T_3276_data : {{11'd0}, 1'h0};
  assign T_3402 = T_2925 ? tgts_T_3278_data : {{11'd0}, 1'h0};
  assign T_3404 = T_2926 ? tgts_T_3280_data : {{11'd0}, 1'h0};
  assign T_3406 = T_2927 ? tgts_T_3282_data : {{11'd0}, 1'h0};
  assign T_3408 = T_2928 ? tgts_T_3284_data : {{11'd0}, 1'h0};
  assign T_3410 = T_2929 ? tgts_T_3286_data : {{11'd0}, 1'h0};
  assign T_3412 = T_2930 ? tgts_T_3288_data : {{11'd0}, 1'h0};
  assign T_3414 = T_2931 ? tgts_T_3290_data : {{11'd0}, 1'h0};
  assign T_3416 = T_2932 ? tgts_T_3292_data : {{11'd0}, 1'h0};
  assign T_3418 = T_2933 ? tgts_T_3294_data : {{11'd0}, 1'h0};
  assign T_3420 = T_2934 ? tgts_T_3296_data : {{11'd0}, 1'h0};
  assign T_3422 = T_2935 ? tgts_T_3298_data : {{11'd0}, 1'h0};
  assign T_3424 = T_2936 ? tgts_T_3300_data : {{11'd0}, 1'h0};
  assign T_3426 = T_2937 ? tgts_T_3302_data : {{11'd0}, 1'h0};
  assign T_3428 = T_2938 ? tgts_T_3304_data : {{11'd0}, 1'h0};
  assign T_3430 = T_2939 ? tgts_T_3306_data : {{11'd0}, 1'h0};
  assign T_3432 = T_2940 ? tgts_T_3308_data : {{11'd0}, 1'h0};
  assign T_3434 = T_2941 ? tgts_T_3310_data : {{11'd0}, 1'h0};
  assign T_3436 = T_2942 ? tgts_T_3312_data : {{11'd0}, 1'h0};
  assign T_3438 = T_2943 ? tgts_T_3314_data : {{11'd0}, 1'h0};
  assign T_3440 = T_2944 ? tgts_T_3316_data : {{11'd0}, 1'h0};
  assign T_3442 = T_2945 ? tgts_T_3318_data : {{11'd0}, 1'h0};
  assign T_3444 = T_2946 ? tgts_T_3320_data : {{11'd0}, 1'h0};
  assign T_3446 = T_2947 ? tgts_T_3322_data : {{11'd0}, 1'h0};
  assign T_3448 = T_2948 ? tgts_T_3324_data : {{11'd0}, 1'h0};
  assign T_3450 = T_2949 ? tgts_T_3326_data : {{11'd0}, 1'h0};
  assign T_3452 = T_2950 ? tgts_T_3328_data : {{11'd0}, 1'h0};
  assign T_3454 = T_2951 ? tgts_T_3330_data : {{11'd0}, 1'h0};
  assign T_3456 = T_2952 ? tgts_T_3332_data : {{11'd0}, 1'h0};
  assign T_3458 = T_2953 ? tgts_T_3334_data : {{11'd0}, 1'h0};
  assign T_3460 = T_2954 ? tgts_T_3336_data : {{11'd0}, 1'h0};
  assign T_3462 = T_2955 ? tgts_T_3338_data : {{11'd0}, 1'h0};
  assign T_3464 = T_2956 ? tgts_T_3340_data : {{11'd0}, 1'h0};
  assign T_3466 = T_2957 ? tgts_T_3342_data : {{11'd0}, 1'h0};
  assign T_3468 = T_2958 ? tgts_T_3344_data : {{11'd0}, 1'h0};
  assign T_3470 = T_2959 ? tgts_T_3346_data : {{11'd0}, 1'h0};
  assign T_3472 = T_2960 ? tgts_T_3348_data : {{11'd0}, 1'h0};
  assign T_3474 = T_2961 ? tgts_T_3350_data : {{11'd0}, 1'h0};
  assign T_3476 = T_2962 ? tgts_T_3352_data : {{11'd0}, 1'h0};
  assign T_3478 = T_2963 ? tgts_T_3354_data : {{11'd0}, 1'h0};
  assign T_3480 = T_2964 ? tgts_T_3356_data : {{11'd0}, 1'h0};
  assign T_3482 = T_2965 ? tgts_T_3358_data : {{11'd0}, 1'h0};
  assign T_3484 = T_2966 ? tgts_T_3360_data : {{11'd0}, 1'h0};
  assign T_3486 = T_2967 ? tgts_T_3362_data : {{11'd0}, 1'h0};
  assign T_3488 = T_2968 ? tgts_T_3364_data : {{11'd0}, 1'h0};
  assign T_3490 = T_2969 ? tgts_T_3366_data : {{11'd0}, 1'h0};
  assign T_3492 = T_2970 ? tgts_T_3368_data : {{11'd0}, 1'h0};
  assign T_3494 = T_2971 ? tgts_T_3370_data : {{11'd0}, 1'h0};
  assign T_3496 = T_2972 ? tgts_T_3372_data : {{11'd0}, 1'h0};
  assign T_3498 = T_2973 ? tgts_T_3374_data : {{11'd0}, 1'h0};
  assign T_3500 = T_2974 ? tgts_T_3376_data : {{11'd0}, 1'h0};
  assign T_3502 = T_2975 ? tgts_T_3378_data : {{11'd0}, 1'h0};
  assign T_3504 = T_2976 ? tgts_T_3380_data : {{11'd0}, 1'h0};
  assign T_3506 = T_2977 ? tgts_T_3382_data : {{11'd0}, 1'h0};
  assign T_3508 = T_2978 ? tgts_T_3384_data : {{11'd0}, 1'h0};
  assign T_3510 = T_2979 ? tgts_T_3386_data : {{11'd0}, 1'h0};
  assign T_3512 = T_2980 ? tgts_T_3388_data : {{11'd0}, 1'h0};
  assign T_3514 = T_2981 ? tgts_T_3390_data : {{11'd0}, 1'h0};
  assign T_3516 = T_2982 ? tgts_T_3392_data : {{11'd0}, 1'h0};
  assign T_3518 = T_3394 | T_3396;
  assign T_3519 = T_3518 | T_3398;
  assign T_3520 = T_3519 | T_3400;
  assign T_3521 = T_3520 | T_3402;
  assign T_3522 = T_3521 | T_3404;
  assign T_3523 = T_3522 | T_3406;
  assign T_3524 = T_3523 | T_3408;
  assign T_3525 = T_3524 | T_3410;
  assign T_3526 = T_3525 | T_3412;
  assign T_3527 = T_3526 | T_3414;
  assign T_3528 = T_3527 | T_3416;
  assign T_3529 = T_3528 | T_3418;
  assign T_3530 = T_3529 | T_3420;
  assign T_3531 = T_3530 | T_3422;
  assign T_3532 = T_3531 | T_3424;
  assign T_3533 = T_3532 | T_3426;
  assign T_3534 = T_3533 | T_3428;
  assign T_3535 = T_3534 | T_3430;
  assign T_3536 = T_3535 | T_3432;
  assign T_3537 = T_3536 | T_3434;
  assign T_3538 = T_3537 | T_3436;
  assign T_3539 = T_3538 | T_3438;
  assign T_3540 = T_3539 | T_3440;
  assign T_3541 = T_3540 | T_3442;
  assign T_3542 = T_3541 | T_3444;
  assign T_3543 = T_3542 | T_3446;
  assign T_3544 = T_3543 | T_3448;
  assign T_3545 = T_3544 | T_3450;
  assign T_3546 = T_3545 | T_3452;
  assign T_3547 = T_3546 | T_3454;
  assign T_3548 = T_3547 | T_3456;
  assign T_3549 = T_3548 | T_3458;
  assign T_3550 = T_3549 | T_3460;
  assign T_3551 = T_3550 | T_3462;
  assign T_3552 = T_3551 | T_3464;
  assign T_3553 = T_3552 | T_3466;
  assign T_3554 = T_3553 | T_3468;
  assign T_3555 = T_3554 | T_3470;
  assign T_3556 = T_3555 | T_3472;
  assign T_3557 = T_3556 | T_3474;
  assign T_3558 = T_3557 | T_3476;
  assign T_3559 = T_3558 | T_3478;
  assign T_3560 = T_3559 | T_3480;
  assign T_3561 = T_3560 | T_3482;
  assign T_3562 = T_3561 | T_3484;
  assign T_3563 = T_3562 | T_3486;
  assign T_3564 = T_3563 | T_3488;
  assign T_3565 = T_3564 | T_3490;
  assign T_3566 = T_3565 | T_3492;
  assign T_3567 = T_3566 | T_3494;
  assign T_3568 = T_3567 | T_3496;
  assign T_3569 = T_3568 | T_3498;
  assign T_3570 = T_3569 | T_3500;
  assign T_3571 = T_3570 | T_3502;
  assign T_3572 = T_3571 | T_3504;
  assign T_3573 = T_3572 | T_3506;
  assign T_3574 = T_3573 | T_3508;
  assign T_3575 = T_3574 | T_3510;
  assign T_3576 = T_3575 | T_3512;
  assign T_3577 = T_3576 | T_3514;
  assign T_3578 = T_3577 | T_3516;
  assign T_3579 = T_3578;
  assign T_3580 = {T_3206,T_3579};
  assign T_3581 = hits[61:32];
  assign T_3582 = hits[31:0];
  assign GEN_848 = {{29'd0}, 1'h0};
  assign T_3584 = T_3581 != GEN_848;
  assign GEN_849 = {{2'd0}, T_3581};
  assign T_3585 = GEN_849 | T_3582;
  assign T_3586 = T_3585[31:16];
  assign T_3587 = T_3585[15:0];
  assign GEN_850 = {{15'd0}, 1'h0};
  assign T_3589 = T_3586 != GEN_850;
  assign T_3590 = T_3586 | T_3587;
  assign T_3591 = T_3590[15:8];
  assign T_3592 = T_3590[7:0];
  assign GEN_851 = {{7'd0}, 1'h0};
  assign T_3594 = T_3591 != GEN_851;
  assign T_3595 = T_3591 | T_3592;
  assign T_3596 = T_3595[7:4];
  assign T_3597 = T_3595[3:0];
  assign GEN_852 = {{3'd0}, 1'h0};
  assign T_3599 = T_3596 != GEN_852;
  assign T_3600 = T_3596 | T_3597;
  assign T_3601 = T_3600[3:2];
  assign T_3602 = T_3600[1:0];
  assign T_3604 = T_3601 != GEN_707;
  assign T_3605 = T_3601 | T_3602;
  assign T_3606 = T_3605[1];
  assign T_3607 = {T_3604,T_3606};
  assign T_3608 = {T_3599,T_3607};
  assign T_3609 = {T_3594,T_3608};
  assign T_3610 = {T_3589,T_3609};
  assign T_3611 = {T_3584,T_3610};
  assign T_3616_T_3942_addr = T_3941;
  assign T_3616_T_3942_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_3616_T_3942_data = T_3616[T_3616_T_3942_addr];
  `else
  assign T_3616_T_3942_data = T_3616_T_3942_addr >= 8'h80 ? $random : T_3616[T_3616_T_3942_addr];
  `endif
  assign T_3616_T_3949_data = T_3958;
  assign T_3616_T_3949_addr = T_3948;
  assign T_3616_T_3949_mask = T_3946;
  assign T_3616_T_3949_en = T_3946;
  assign T_3683 = T_2921 ? isJump_0 : 1'h0;
  assign T_3686 = T_2922 ? isJump_1 : 1'h0;
  assign T_3689 = T_2923 ? isJump_2 : 1'h0;
  assign T_3692 = T_2924 ? isJump_3 : 1'h0;
  assign T_3695 = T_2925 ? isJump_4 : 1'h0;
  assign T_3698 = T_2926 ? isJump_5 : 1'h0;
  assign T_3701 = T_2927 ? isJump_6 : 1'h0;
  assign T_3704 = T_2928 ? isJump_7 : 1'h0;
  assign T_3707 = T_2929 ? isJump_8 : 1'h0;
  assign T_3710 = T_2930 ? isJump_9 : 1'h0;
  assign T_3713 = T_2931 ? isJump_10 : 1'h0;
  assign T_3716 = T_2932 ? isJump_11 : 1'h0;
  assign T_3719 = T_2933 ? isJump_12 : 1'h0;
  assign T_3722 = T_2934 ? isJump_13 : 1'h0;
  assign T_3725 = T_2935 ? isJump_14 : 1'h0;
  assign T_3728 = T_2936 ? isJump_15 : 1'h0;
  assign T_3731 = T_2937 ? isJump_16 : 1'h0;
  assign T_3734 = T_2938 ? isJump_17 : 1'h0;
  assign T_3737 = T_2939 ? isJump_18 : 1'h0;
  assign T_3740 = T_2940 ? isJump_19 : 1'h0;
  assign T_3743 = T_2941 ? isJump_20 : 1'h0;
  assign T_3746 = T_2942 ? isJump_21 : 1'h0;
  assign T_3749 = T_2943 ? isJump_22 : 1'h0;
  assign T_3752 = T_2944 ? isJump_23 : 1'h0;
  assign T_3755 = T_2945 ? isJump_24 : 1'h0;
  assign T_3758 = T_2946 ? isJump_25 : 1'h0;
  assign T_3761 = T_2947 ? isJump_26 : 1'h0;
  assign T_3764 = T_2948 ? isJump_27 : 1'h0;
  assign T_3767 = T_2949 ? isJump_28 : 1'h0;
  assign T_3770 = T_2950 ? isJump_29 : 1'h0;
  assign T_3773 = T_2951 ? isJump_30 : 1'h0;
  assign T_3776 = T_2952 ? isJump_31 : 1'h0;
  assign T_3779 = T_2953 ? isJump_32 : 1'h0;
  assign T_3782 = T_2954 ? isJump_33 : 1'h0;
  assign T_3785 = T_2955 ? isJump_34 : 1'h0;
  assign T_3788 = T_2956 ? isJump_35 : 1'h0;
  assign T_3791 = T_2957 ? isJump_36 : 1'h0;
  assign T_3794 = T_2958 ? isJump_37 : 1'h0;
  assign T_3797 = T_2959 ? isJump_38 : 1'h0;
  assign T_3800 = T_2960 ? isJump_39 : 1'h0;
  assign T_3803 = T_2961 ? isJump_40 : 1'h0;
  assign T_3806 = T_2962 ? isJump_41 : 1'h0;
  assign T_3809 = T_2963 ? isJump_42 : 1'h0;
  assign T_3812 = T_2964 ? isJump_43 : 1'h0;
  assign T_3815 = T_2965 ? isJump_44 : 1'h0;
  assign T_3818 = T_2966 ? isJump_45 : 1'h0;
  assign T_3821 = T_2967 ? isJump_46 : 1'h0;
  assign T_3824 = T_2968 ? isJump_47 : 1'h0;
  assign T_3827 = T_2969 ? isJump_48 : 1'h0;
  assign T_3830 = T_2970 ? isJump_49 : 1'h0;
  assign T_3833 = T_2971 ? isJump_50 : 1'h0;
  assign T_3836 = T_2972 ? isJump_51 : 1'h0;
  assign T_3839 = T_2973 ? isJump_52 : 1'h0;
  assign T_3842 = T_2974 ? isJump_53 : 1'h0;
  assign T_3845 = T_2975 ? isJump_54 : 1'h0;
  assign T_3848 = T_2976 ? isJump_55 : 1'h0;
  assign T_3851 = T_2977 ? isJump_56 : 1'h0;
  assign T_3854 = T_2978 ? isJump_57 : 1'h0;
  assign T_3857 = T_2979 ? isJump_58 : 1'h0;
  assign T_3860 = T_2980 ? isJump_59 : 1'h0;
  assign T_3863 = T_2981 ? isJump_60 : 1'h0;
  assign T_3866 = T_2982 ? isJump_61 : 1'h0;
  assign T_3868 = T_3683 | T_3686;
  assign T_3869 = T_3868 | T_3689;
  assign T_3870 = T_3869 | T_3692;
  assign T_3871 = T_3870 | T_3695;
  assign T_3872 = T_3871 | T_3698;
  assign T_3873 = T_3872 | T_3701;
  assign T_3874 = T_3873 | T_3704;
  assign T_3875 = T_3874 | T_3707;
  assign T_3876 = T_3875 | T_3710;
  assign T_3877 = T_3876 | T_3713;
  assign T_3878 = T_3877 | T_3716;
  assign T_3879 = T_3878 | T_3719;
  assign T_3880 = T_3879 | T_3722;
  assign T_3881 = T_3880 | T_3725;
  assign T_3882 = T_3881 | T_3728;
  assign T_3883 = T_3882 | T_3731;
  assign T_3884 = T_3883 | T_3734;
  assign T_3885 = T_3884 | T_3737;
  assign T_3886 = T_3885 | T_3740;
  assign T_3887 = T_3886 | T_3743;
  assign T_3888 = T_3887 | T_3746;
  assign T_3889 = T_3888 | T_3749;
  assign T_3890 = T_3889 | T_3752;
  assign T_3891 = T_3890 | T_3755;
  assign T_3892 = T_3891 | T_3758;
  assign T_3893 = T_3892 | T_3761;
  assign T_3894 = T_3893 | T_3764;
  assign T_3895 = T_3894 | T_3767;
  assign T_3896 = T_3895 | T_3770;
  assign T_3897 = T_3896 | T_3773;
  assign T_3898 = T_3897 | T_3776;
  assign T_3899 = T_3898 | T_3779;
  assign T_3900 = T_3899 | T_3782;
  assign T_3901 = T_3900 | T_3785;
  assign T_3902 = T_3901 | T_3788;
  assign T_3903 = T_3902 | T_3791;
  assign T_3904 = T_3903 | T_3794;
  assign T_3905 = T_3904 | T_3797;
  assign T_3906 = T_3905 | T_3800;
  assign T_3907 = T_3906 | T_3803;
  assign T_3908 = T_3907 | T_3806;
  assign T_3909 = T_3908 | T_3809;
  assign T_3910 = T_3909 | T_3812;
  assign T_3911 = T_3910 | T_3815;
  assign T_3912 = T_3911 | T_3818;
  assign T_3913 = T_3912 | T_3821;
  assign T_3914 = T_3913 | T_3824;
  assign T_3915 = T_3914 | T_3827;
  assign T_3916 = T_3915 | T_3830;
  assign T_3917 = T_3916 | T_3833;
  assign T_3918 = T_3917 | T_3836;
  assign T_3919 = T_3918 | T_3839;
  assign T_3920 = T_3919 | T_3842;
  assign T_3921 = T_3920 | T_3845;
  assign T_3922 = T_3921 | T_3848;
  assign T_3923 = T_3922 | T_3851;
  assign T_3924 = T_3923 | T_3854;
  assign T_3925 = T_3924 | T_3857;
  assign T_3926 = T_3925 | T_3860;
  assign T_3927 = T_3926 | T_3863;
  assign T_3928 = T_3927 | T_3866;
  assign T_3929 = T_3928;
  assign T_3931 = T_3929 == 1'h0;
  assign T_3932 = io_req_valid & io_resp_valid;
  assign T_3933 = T_3932 & T_3931;
  assign T_3937_history = T_3618;
  assign T_3937_value = T_3616_T_3942_data;
  assign T_3940 = io_req_bits_addr[8:2];
  assign T_3941 = T_3940 ^ T_3618;
  assign T_3943 = T_3937_value[0];
  assign T_3944 = T_3618[6:1];
  assign T_3945 = {T_3943,T_3944};
  assign GEN_424 = T_3933 ? T_3945 : T_3618;
  assign T_3946 = io_bht_update_valid & io_bht_update_bits_prediction_valid;
  assign T_3947 = io_bht_update_bits_pc[8:2];
  assign T_3948 = T_3947 ^ io_bht_update_bits_prediction_bits_bht_history;
  assign T_3950 = io_bht_update_bits_prediction_bits_bht_value[1];
  assign T_3951 = io_bht_update_bits_prediction_bits_bht_value[0];
  assign T_3952 = T_3950 & T_3951;
  assign T_3955 = T_3950 | T_3951;
  assign T_3956 = T_3955 & io_bht_update_bits_taken;
  assign T_3957 = T_3952 | T_3956;
  assign T_3958 = {io_bht_update_bits_taken,T_3957};
  assign T_3959 = io_bht_update_bits_prediction_bits_bht_history[6:1];
  assign T_3960 = {io_bht_update_bits_taken,T_3959};
  assign GEN_425 = io_bht_update_bits_mispredict ? T_3960 : GEN_424;
  assign GEN_431 = T_3946 ? GEN_425 : GEN_424;
  assign T_3963 = T_3943 == 1'h0;
  assign T_3964 = T_3963 & T_3931;
  assign GEN_432 = T_3964 ? 1'h0 : io_resp_valid;
  assign T_4042 = T_2921 ? useRAS_0 : 1'h0;
  assign T_4045 = T_2922 ? useRAS_1 : 1'h0;
  assign T_4048 = T_2923 ? useRAS_2 : 1'h0;
  assign T_4051 = T_2924 ? useRAS_3 : 1'h0;
  assign T_4054 = T_2925 ? useRAS_4 : 1'h0;
  assign T_4057 = T_2926 ? useRAS_5 : 1'h0;
  assign T_4060 = T_2927 ? useRAS_6 : 1'h0;
  assign T_4063 = T_2928 ? useRAS_7 : 1'h0;
  assign T_4066 = T_2929 ? useRAS_8 : 1'h0;
  assign T_4069 = T_2930 ? useRAS_9 : 1'h0;
  assign T_4072 = T_2931 ? useRAS_10 : 1'h0;
  assign T_4075 = T_2932 ? useRAS_11 : 1'h0;
  assign T_4078 = T_2933 ? useRAS_12 : 1'h0;
  assign T_4081 = T_2934 ? useRAS_13 : 1'h0;
  assign T_4084 = T_2935 ? useRAS_14 : 1'h0;
  assign T_4087 = T_2936 ? useRAS_15 : 1'h0;
  assign T_4090 = T_2937 ? useRAS_16 : 1'h0;
  assign T_4093 = T_2938 ? useRAS_17 : 1'h0;
  assign T_4096 = T_2939 ? useRAS_18 : 1'h0;
  assign T_4099 = T_2940 ? useRAS_19 : 1'h0;
  assign T_4102 = T_2941 ? useRAS_20 : 1'h0;
  assign T_4105 = T_2942 ? useRAS_21 : 1'h0;
  assign T_4108 = T_2943 ? useRAS_22 : 1'h0;
  assign T_4111 = T_2944 ? useRAS_23 : 1'h0;
  assign T_4114 = T_2945 ? useRAS_24 : 1'h0;
  assign T_4117 = T_2946 ? useRAS_25 : 1'h0;
  assign T_4120 = T_2947 ? useRAS_26 : 1'h0;
  assign T_4123 = T_2948 ? useRAS_27 : 1'h0;
  assign T_4126 = T_2949 ? useRAS_28 : 1'h0;
  assign T_4129 = T_2950 ? useRAS_29 : 1'h0;
  assign T_4132 = T_2951 ? useRAS_30 : 1'h0;
  assign T_4135 = T_2952 ? useRAS_31 : 1'h0;
  assign T_4138 = T_2953 ? useRAS_32 : 1'h0;
  assign T_4141 = T_2954 ? useRAS_33 : 1'h0;
  assign T_4144 = T_2955 ? useRAS_34 : 1'h0;
  assign T_4147 = T_2956 ? useRAS_35 : 1'h0;
  assign T_4150 = T_2957 ? useRAS_36 : 1'h0;
  assign T_4153 = T_2958 ? useRAS_37 : 1'h0;
  assign T_4156 = T_2959 ? useRAS_38 : 1'h0;
  assign T_4159 = T_2960 ? useRAS_39 : 1'h0;
  assign T_4162 = T_2961 ? useRAS_40 : 1'h0;
  assign T_4165 = T_2962 ? useRAS_41 : 1'h0;
  assign T_4168 = T_2963 ? useRAS_42 : 1'h0;
  assign T_4171 = T_2964 ? useRAS_43 : 1'h0;
  assign T_4174 = T_2965 ? useRAS_44 : 1'h0;
  assign T_4177 = T_2966 ? useRAS_45 : 1'h0;
  assign T_4180 = T_2967 ? useRAS_46 : 1'h0;
  assign T_4183 = T_2968 ? useRAS_47 : 1'h0;
  assign T_4186 = T_2969 ? useRAS_48 : 1'h0;
  assign T_4189 = T_2970 ? useRAS_49 : 1'h0;
  assign T_4192 = T_2971 ? useRAS_50 : 1'h0;
  assign T_4195 = T_2972 ? useRAS_51 : 1'h0;
  assign T_4198 = T_2973 ? useRAS_52 : 1'h0;
  assign T_4201 = T_2974 ? useRAS_53 : 1'h0;
  assign T_4204 = T_2975 ? useRAS_54 : 1'h0;
  assign T_4207 = T_2976 ? useRAS_55 : 1'h0;
  assign T_4210 = T_2977 ? useRAS_56 : 1'h0;
  assign T_4213 = T_2978 ? useRAS_57 : 1'h0;
  assign T_4216 = T_2979 ? useRAS_58 : 1'h0;
  assign T_4219 = T_2980 ? useRAS_59 : 1'h0;
  assign T_4222 = T_2981 ? useRAS_60 : 1'h0;
  assign T_4225 = T_2982 ? useRAS_61 : 1'h0;
  assign T_4227 = T_4042 | T_4045;
  assign T_4228 = T_4227 | T_4048;
  assign T_4229 = T_4228 | T_4051;
  assign T_4230 = T_4229 | T_4054;
  assign T_4231 = T_4230 | T_4057;
  assign T_4232 = T_4231 | T_4060;
  assign T_4233 = T_4232 | T_4063;
  assign T_4234 = T_4233 | T_4066;
  assign T_4235 = T_4234 | T_4069;
  assign T_4236 = T_4235 | T_4072;
  assign T_4237 = T_4236 | T_4075;
  assign T_4238 = T_4237 | T_4078;
  assign T_4239 = T_4238 | T_4081;
  assign T_4240 = T_4239 | T_4084;
  assign T_4241 = T_4240 | T_4087;
  assign T_4242 = T_4241 | T_4090;
  assign T_4243 = T_4242 | T_4093;
  assign T_4244 = T_4243 | T_4096;
  assign T_4245 = T_4244 | T_4099;
  assign T_4246 = T_4245 | T_4102;
  assign T_4247 = T_4246 | T_4105;
  assign T_4248 = T_4247 | T_4108;
  assign T_4249 = T_4248 | T_4111;
  assign T_4250 = T_4249 | T_4114;
  assign T_4251 = T_4250 | T_4117;
  assign T_4252 = T_4251 | T_4120;
  assign T_4253 = T_4252 | T_4123;
  assign T_4254 = T_4253 | T_4126;
  assign T_4255 = T_4254 | T_4129;
  assign T_4256 = T_4255 | T_4132;
  assign T_4257 = T_4256 | T_4135;
  assign T_4258 = T_4257 | T_4138;
  assign T_4259 = T_4258 | T_4141;
  assign T_4260 = T_4259 | T_4144;
  assign T_4261 = T_4260 | T_4147;
  assign T_4262 = T_4261 | T_4150;
  assign T_4263 = T_4262 | T_4153;
  assign T_4264 = T_4263 | T_4156;
  assign T_4265 = T_4264 | T_4159;
  assign T_4266 = T_4265 | T_4162;
  assign T_4267 = T_4266 | T_4165;
  assign T_4268 = T_4267 | T_4168;
  assign T_4269 = T_4268 | T_4171;
  assign T_4270 = T_4269 | T_4174;
  assign T_4271 = T_4270 | T_4177;
  assign T_4272 = T_4271 | T_4180;
  assign T_4273 = T_4272 | T_4183;
  assign T_4274 = T_4273 | T_4186;
  assign T_4275 = T_4274 | T_4189;
  assign T_4276 = T_4275 | T_4192;
  assign T_4277 = T_4276 | T_4195;
  assign T_4278 = T_4277 | T_4198;
  assign T_4279 = T_4278 | T_4201;
  assign T_4280 = T_4279 | T_4204;
  assign T_4281 = T_4280 | T_4207;
  assign T_4282 = T_4281 | T_4210;
  assign T_4283 = T_4282 | T_4213;
  assign T_4284 = T_4283 | T_4216;
  assign T_4285 = T_4284 | T_4219;
  assign T_4286 = T_4285 | T_4222;
  assign T_4287 = T_4286 | T_4225;
  assign T_4288 = T_4287;
  assign T_4290 = T_3967 == GEN_707;
  assign T_4292 = T_4290 == 1'h0;
  assign T_4293 = T_4292 & T_4288;
  assign GEN_2 = GEN_433;
  assign GEN_433 = T_3969 ? T_3976_1 : T_3976_0;
  assign GEN_435 = T_4293 ? GEN_2 : T_3580;
  assign T_4295 = T_3967 < 2'h2;
  assign GEN_855 = {{1'd0}, 1'h1};
  assign T_4297 = T_3967 + GEN_855;
  assign T_4298 = T_4297[1:0];
  assign GEN_436 = T_4295 ? T_4298 : T_3967;
  assign T_4304 = T_3969 + 1'h1;
  assign T_4305 = T_4304[0:0];
  assign GEN_3 = io_ras_update_bits_returnAddr;
  assign GEN_437 = 1'h0 == T_4305 ? GEN_3 : T_3976_0;
  assign GEN_438 = T_4305 ? GEN_3 : T_3976_1;
  assign GEN_439 = T_4288 ? io_ras_update_bits_returnAddr : GEN_435;
  assign GEN_440 = io_ras_update_bits_isCall ? GEN_436 : T_3967;
  assign GEN_442 = io_ras_update_bits_isCall ? GEN_437 : T_3976_0;
  assign GEN_443 = io_ras_update_bits_isCall ? GEN_438 : T_3976_1;
  assign GEN_444 = io_ras_update_bits_isCall ? T_4305 : T_3969;
  assign GEN_445 = io_ras_update_bits_isCall ? GEN_439 : GEN_435;
  assign T_4308 = io_ras_update_bits_isReturn & io_ras_update_bits_prediction_valid;
  assign T_4310 = io_ras_update_bits_isCall == 1'h0;
  assign T_4311 = T_4310 & T_4308;
  assign T_4317 = T_3967 - GEN_855;
  assign T_4318 = T_4317[1:0];
  assign T_4324 = T_3969 - 1'h1;
  assign T_4325 = T_4324[0:0];
  assign GEN_446 = T_4292 ? T_4318 : GEN_440;
  assign GEN_447 = T_4292 ? T_4325 : GEN_444;
  assign GEN_448 = T_4311 ? GEN_446 : GEN_440;
  assign GEN_449 = T_4311 ? GEN_447 : GEN_444;
  assign GEN_450 = io_ras_update_valid ? GEN_448 : T_3967;
  assign GEN_452 = io_ras_update_valid ? GEN_442 : T_3976_0;
  assign GEN_453 = io_ras_update_valid ? GEN_443 : T_3976_1;
  assign GEN_454 = io_ras_update_valid ? GEN_449 : T_3969;
  assign GEN_455 = io_ras_update_valid ? GEN_445 : GEN_435;
  assign GEN_456 = io_invalidate ? {{1'd0}, 1'h0} : GEN_450;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_146 = {2{$random}};
  idxValid = GEN_146[61:0];
  GEN_147 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    idxs[initvar] = GEN_147[11:0];
  GEN_148 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    idxPages[initvar] = GEN_148[2:0];
  GEN_149 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    tgts[initvar] = GEN_149[11:0];
  GEN_150 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    tgtPages[initvar] = GEN_150[2:0];
  GEN_151 = {1{$random}};
  for (initvar = 0; initvar < 6; initvar = initvar+1)
    pages[initvar] = GEN_151[26:0];
  GEN_152 = {1{$random}};
  pageValid = GEN_152[5:0];
  GEN_153 = {1{$random}};
  useRAS_0 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  useRAS_1 = GEN_154[0:0];
  GEN_155 = {1{$random}};
  useRAS_2 = GEN_155[0:0];
  GEN_156 = {1{$random}};
  useRAS_3 = GEN_156[0:0];
  GEN_157 = {1{$random}};
  useRAS_4 = GEN_157[0:0];
  GEN_158 = {1{$random}};
  useRAS_5 = GEN_158[0:0];
  GEN_159 = {1{$random}};
  useRAS_6 = GEN_159[0:0];
  GEN_160 = {1{$random}};
  useRAS_7 = GEN_160[0:0];
  GEN_161 = {1{$random}};
  useRAS_8 = GEN_161[0:0];
  GEN_162 = {1{$random}};
  useRAS_9 = GEN_162[0:0];
  GEN_163 = {1{$random}};
  useRAS_10 = GEN_163[0:0];
  GEN_164 = {1{$random}};
  useRAS_11 = GEN_164[0:0];
  GEN_165 = {1{$random}};
  useRAS_12 = GEN_165[0:0];
  GEN_166 = {1{$random}};
  useRAS_13 = GEN_166[0:0];
  GEN_167 = {1{$random}};
  useRAS_14 = GEN_167[0:0];
  GEN_168 = {1{$random}};
  useRAS_15 = GEN_168[0:0];
  GEN_169 = {1{$random}};
  useRAS_16 = GEN_169[0:0];
  GEN_170 = {1{$random}};
  useRAS_17 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  useRAS_18 = GEN_171[0:0];
  GEN_172 = {1{$random}};
  useRAS_19 = GEN_172[0:0];
  GEN_173 = {1{$random}};
  useRAS_20 = GEN_173[0:0];
  GEN_174 = {1{$random}};
  useRAS_21 = GEN_174[0:0];
  GEN_175 = {1{$random}};
  useRAS_22 = GEN_175[0:0];
  GEN_177 = {1{$random}};
  useRAS_23 = GEN_177[0:0];
  GEN_178 = {1{$random}};
  useRAS_24 = GEN_178[0:0];
  GEN_179 = {1{$random}};
  useRAS_25 = GEN_179[0:0];
  GEN_180 = {1{$random}};
  useRAS_26 = GEN_180[0:0];
  GEN_181 = {1{$random}};
  useRAS_27 = GEN_181[0:0];
  GEN_182 = {1{$random}};
  useRAS_28 = GEN_182[0:0];
  GEN_183 = {1{$random}};
  useRAS_29 = GEN_183[0:0];
  GEN_184 = {1{$random}};
  useRAS_30 = GEN_184[0:0];
  GEN_185 = {1{$random}};
  useRAS_31 = GEN_185[0:0];
  GEN_186 = {1{$random}};
  useRAS_32 = GEN_186[0:0];
  GEN_187 = {1{$random}};
  useRAS_33 = GEN_187[0:0];
  GEN_188 = {1{$random}};
  useRAS_34 = GEN_188[0:0];
  GEN_189 = {1{$random}};
  useRAS_35 = GEN_189[0:0];
  GEN_190 = {1{$random}};
  useRAS_36 = GEN_190[0:0];
  GEN_191 = {1{$random}};
  useRAS_37 = GEN_191[0:0];
  GEN_192 = {1{$random}};
  useRAS_38 = GEN_192[0:0];
  GEN_193 = {1{$random}};
  useRAS_39 = GEN_193[0:0];
  GEN_194 = {1{$random}};
  useRAS_40 = GEN_194[0:0];
  GEN_195 = {1{$random}};
  useRAS_41 = GEN_195[0:0];
  GEN_196 = {1{$random}};
  useRAS_42 = GEN_196[0:0];
  GEN_197 = {1{$random}};
  useRAS_43 = GEN_197[0:0];
  GEN_198 = {1{$random}};
  useRAS_44 = GEN_198[0:0];
  GEN_199 = {1{$random}};
  useRAS_45 = GEN_199[0:0];
  GEN_200 = {1{$random}};
  useRAS_46 = GEN_200[0:0];
  GEN_201 = {1{$random}};
  useRAS_47 = GEN_201[0:0];
  GEN_202 = {1{$random}};
  useRAS_48 = GEN_202[0:0];
  GEN_203 = {1{$random}};
  useRAS_49 = GEN_203[0:0];
  GEN_204 = {1{$random}};
  useRAS_50 = GEN_204[0:0];
  GEN_205 = {1{$random}};
  useRAS_51 = GEN_205[0:0];
  GEN_206 = {1{$random}};
  useRAS_52 = GEN_206[0:0];
  GEN_207 = {1{$random}};
  useRAS_53 = GEN_207[0:0];
  GEN_208 = {1{$random}};
  useRAS_54 = GEN_208[0:0];
  GEN_209 = {1{$random}};
  useRAS_55 = GEN_209[0:0];
  GEN_210 = {1{$random}};
  useRAS_56 = GEN_210[0:0];
  GEN_211 = {1{$random}};
  useRAS_57 = GEN_211[0:0];
  GEN_212 = {1{$random}};
  useRAS_58 = GEN_212[0:0];
  GEN_213 = {1{$random}};
  useRAS_59 = GEN_213[0:0];
  GEN_214 = {1{$random}};
  useRAS_60 = GEN_214[0:0];
  GEN_215 = {1{$random}};
  useRAS_61 = GEN_215[0:0];
  GEN_216 = {1{$random}};
  isJump_0 = GEN_216[0:0];
  GEN_217 = {1{$random}};
  isJump_1 = GEN_217[0:0];
  GEN_218 = {1{$random}};
  isJump_2 = GEN_218[0:0];
  GEN_219 = {1{$random}};
  isJump_3 = GEN_219[0:0];
  GEN_220 = {1{$random}};
  isJump_4 = GEN_220[0:0];
  GEN_221 = {1{$random}};
  isJump_5 = GEN_221[0:0];
  GEN_222 = {1{$random}};
  isJump_6 = GEN_222[0:0];
  GEN_223 = {1{$random}};
  isJump_7 = GEN_223[0:0];
  GEN_224 = {1{$random}};
  isJump_8 = GEN_224[0:0];
  GEN_225 = {1{$random}};
  isJump_9 = GEN_225[0:0];
  GEN_226 = {1{$random}};
  isJump_10 = GEN_226[0:0];
  GEN_227 = {1{$random}};
  isJump_11 = GEN_227[0:0];
  GEN_228 = {1{$random}};
  isJump_12 = GEN_228[0:0];
  GEN_229 = {1{$random}};
  isJump_13 = GEN_229[0:0];
  GEN_230 = {1{$random}};
  isJump_14 = GEN_230[0:0];
  GEN_231 = {1{$random}};
  isJump_15 = GEN_231[0:0];
  GEN_232 = {1{$random}};
  isJump_16 = GEN_232[0:0];
  GEN_233 = {1{$random}};
  isJump_17 = GEN_233[0:0];
  GEN_234 = {1{$random}};
  isJump_18 = GEN_234[0:0];
  GEN_235 = {1{$random}};
  isJump_19 = GEN_235[0:0];
  GEN_236 = {1{$random}};
  isJump_20 = GEN_236[0:0];
  GEN_237 = {1{$random}};
  isJump_21 = GEN_237[0:0];
  GEN_238 = {1{$random}};
  isJump_22 = GEN_238[0:0];
  GEN_240 = {1{$random}};
  isJump_23 = GEN_240[0:0];
  GEN_241 = {1{$random}};
  isJump_24 = GEN_241[0:0];
  GEN_242 = {1{$random}};
  isJump_25 = GEN_242[0:0];
  GEN_243 = {1{$random}};
  isJump_26 = GEN_243[0:0];
  GEN_244 = {1{$random}};
  isJump_27 = GEN_244[0:0];
  GEN_245 = {1{$random}};
  isJump_28 = GEN_245[0:0];
  GEN_246 = {1{$random}};
  isJump_29 = GEN_246[0:0];
  GEN_247 = {1{$random}};
  isJump_30 = GEN_247[0:0];
  GEN_248 = {1{$random}};
  isJump_31 = GEN_248[0:0];
  GEN_249 = {1{$random}};
  isJump_32 = GEN_249[0:0];
  GEN_250 = {1{$random}};
  isJump_33 = GEN_250[0:0];
  GEN_251 = {1{$random}};
  isJump_34 = GEN_251[0:0];
  GEN_252 = {1{$random}};
  isJump_35 = GEN_252[0:0];
  GEN_253 = {1{$random}};
  isJump_36 = GEN_253[0:0];
  GEN_254 = {1{$random}};
  isJump_37 = GEN_254[0:0];
  GEN_255 = {1{$random}};
  isJump_38 = GEN_255[0:0];
  GEN_256 = {1{$random}};
  isJump_39 = GEN_256[0:0];
  GEN_257 = {1{$random}};
  isJump_40 = GEN_257[0:0];
  GEN_258 = {1{$random}};
  isJump_41 = GEN_258[0:0];
  GEN_259 = {1{$random}};
  isJump_42 = GEN_259[0:0];
  GEN_260 = {1{$random}};
  isJump_43 = GEN_260[0:0];
  GEN_323 = {1{$random}};
  isJump_44 = GEN_323[0:0];
  GEN_386 = {1{$random}};
  isJump_45 = GEN_386[0:0];
  GEN_387 = {1{$random}};
  isJump_46 = GEN_387[0:0];
  GEN_388 = {1{$random}};
  isJump_47 = GEN_388[0:0];
  GEN_389 = {1{$random}};
  isJump_48 = GEN_389[0:0];
  GEN_390 = {1{$random}};
  isJump_49 = GEN_390[0:0];
  GEN_391 = {1{$random}};
  isJump_50 = GEN_391[0:0];
  GEN_392 = {1{$random}};
  isJump_51 = GEN_392[0:0];
  GEN_394 = {1{$random}};
  isJump_52 = GEN_394[0:0];
  GEN_395 = {1{$random}};
  isJump_53 = GEN_395[0:0];
  GEN_396 = {1{$random}};
  isJump_54 = GEN_396[0:0];
  GEN_397 = {1{$random}};
  isJump_55 = GEN_397[0:0];
  GEN_399 = {1{$random}};
  isJump_56 = GEN_399[0:0];
  GEN_400 = {1{$random}};
  isJump_57 = GEN_400[0:0];
  GEN_401 = {1{$random}};
  isJump_58 = GEN_401[0:0];
  GEN_402 = {1{$random}};
  isJump_59 = GEN_402[0:0];
  GEN_404 = {1{$random}};
  isJump_60 = GEN_404[0:0];
  GEN_405 = {1{$random}};
  isJump_61 = GEN_405[0:0];
  GEN_406 = {1{$random}};
  for (initvar = 0; initvar < 62; initvar = initvar+1)
    brIdx[initvar] = GEN_406[0:0];
  GEN_407 = {1{$random}};
  T_1215 = GEN_407[0:0];
  GEN_409 = {1{$random}};
  T_1216_prediction_valid = GEN_409[0:0];
  GEN_410 = {1{$random}};
  T_1216_prediction_bits_taken = GEN_410[0:0];
  GEN_411 = {1{$random}};
  T_1216_prediction_bits_mask = GEN_411[0:0];
  GEN_412 = {1{$random}};
  T_1216_prediction_bits_bridx = GEN_412[0:0];
  GEN_414 = {2{$random}};
  T_1216_prediction_bits_target = GEN_414[38:0];
  GEN_415 = {1{$random}};
  T_1216_prediction_bits_entry = GEN_415[5:0];
  GEN_416 = {1{$random}};
  T_1216_prediction_bits_bht_history = GEN_416[6:0];
  GEN_417 = {1{$random}};
  T_1216_prediction_bits_bht_value = GEN_417[1:0];
  GEN_419 = {2{$random}};
  T_1216_pc = GEN_419[38:0];
  GEN_420 = {2{$random}};
  T_1216_target = GEN_420[38:0];
  GEN_426 = {1{$random}};
  T_1216_taken = GEN_426[0:0];
  GEN_427 = {1{$random}};
  T_1216_isJump = GEN_427[0:0];
  GEN_428 = {1{$random}};
  T_1216_isReturn = GEN_428[0:0];
  GEN_429 = {2{$random}};
  T_1216_br_pc = GEN_429[38:0];
  GEN_430 = {1{$random}};
  nextRepl = GEN_430[5:0];
  GEN_434 = {1{$random}};
  T_2536 = GEN_434[2:0];
  GEN_441 = {1{$random}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    T_3616[initvar] = GEN_441[1:0];
  GEN_451 = {1{$random}};
  T_3618 = GEN_451[6:0];
  GEN_458 = {1{$random}};
  T_3967 = GEN_458[1:0];
  GEN_459 = {1{$random}};
  T_3969 = GEN_459[0:0];
  GEN_460 = {2{$random}};
  T_3976_0 = GEN_460[38:0];
  GEN_461 = {2{$random}};
  T_3976_1 = GEN_461[38:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      idxValid <= 62'h0;
    end else begin
      idxValid <= GEN_422[61:0];
    end
    if(idxs_T_2872_en & idxs_T_2872_mask) begin
      idxs[idxs_T_2872_addr] <= idxs_T_2872_data;
    end
    if(idxPages_T_2874_en & idxPages_T_2874_mask) begin
      idxPages[idxPages_T_2874_addr] <= idxPages_T_2874_data;
    end
    if(tgts_T_2873_en & tgts_T_2873_mask) begin
      tgts[tgts_T_2873_addr] <= tgts_T_2873_data;
    end
    if(tgtPages_T_2875_en & tgtPages_T_2875_mask) begin
      tgtPages[tgtPages_T_2875_addr] <= tgtPages_T_2875_data;
    end
    if(pages_T_2891_en & pages_T_2891_mask) begin
      pages[pages_T_2891_addr] <= pages_T_2891_data;
    end
    if(pages_T_2895_en & pages_T_2895_mask) begin
      pages[pages_T_2895_addr] <= pages_T_2895_data;
    end
    if(pages_T_2899_en & pages_T_2899_mask) begin
      pages[pages_T_2899_addr] <= pages_T_2899_data;
    end
    if(pages_T_2907_en & pages_T_2907_mask) begin
      pages[pages_T_2907_addr] <= pages_T_2907_data;
    end
    if(pages_T_2911_en & pages_T_2911_mask) begin
      pages[pages_T_2911_addr] <= pages_T_2911_data;
    end
    if(pages_T_2915_en & pages_T_2915_mask) begin
      pages[pages_T_2915_addr] <= pages_T_2915_data;
    end
    if(reset) begin
      pageValid <= 6'h0;
    end else begin
      pageValid <= GEN_423;
    end
    if(1'h0) begin
    end else begin
      useRAS_0 <= GEN_261;
    end
    if(1'h0) begin
    end else begin
      useRAS_1 <= GEN_262;
    end
    if(1'h0) begin
    end else begin
      useRAS_2 <= GEN_263;
    end
    if(1'h0) begin
    end else begin
      useRAS_3 <= GEN_264;
    end
    if(1'h0) begin
    end else begin
      useRAS_4 <= GEN_265;
    end
    if(1'h0) begin
    end else begin
      useRAS_5 <= GEN_266;
    end
    if(1'h0) begin
    end else begin
      useRAS_6 <= GEN_267;
    end
    if(1'h0) begin
    end else begin
      useRAS_7 <= GEN_268;
    end
    if(1'h0) begin
    end else begin
      useRAS_8 <= GEN_269;
    end
    if(1'h0) begin
    end else begin
      useRAS_9 <= GEN_270;
    end
    if(1'h0) begin
    end else begin
      useRAS_10 <= GEN_271;
    end
    if(1'h0) begin
    end else begin
      useRAS_11 <= GEN_272;
    end
    if(1'h0) begin
    end else begin
      useRAS_12 <= GEN_273;
    end
    if(1'h0) begin
    end else begin
      useRAS_13 <= GEN_274;
    end
    if(1'h0) begin
    end else begin
      useRAS_14 <= GEN_275;
    end
    if(1'h0) begin
    end else begin
      useRAS_15 <= GEN_276;
    end
    if(1'h0) begin
    end else begin
      useRAS_16 <= GEN_277;
    end
    if(1'h0) begin
    end else begin
      useRAS_17 <= GEN_278;
    end
    if(1'h0) begin
    end else begin
      useRAS_18 <= GEN_279;
    end
    if(1'h0) begin
    end else begin
      useRAS_19 <= GEN_280;
    end
    if(1'h0) begin
    end else begin
      useRAS_20 <= GEN_281;
    end
    if(1'h0) begin
    end else begin
      useRAS_21 <= GEN_282;
    end
    if(1'h0) begin
    end else begin
      useRAS_22 <= GEN_283;
    end
    if(1'h0) begin
    end else begin
      useRAS_23 <= GEN_284;
    end
    if(1'h0) begin
    end else begin
      useRAS_24 <= GEN_285;
    end
    if(1'h0) begin
    end else begin
      useRAS_25 <= GEN_286;
    end
    if(1'h0) begin
    end else begin
      useRAS_26 <= GEN_287;
    end
    if(1'h0) begin
    end else begin
      useRAS_27 <= GEN_288;
    end
    if(1'h0) begin
    end else begin
      useRAS_28 <= GEN_289;
    end
    if(1'h0) begin
    end else begin
      useRAS_29 <= GEN_290;
    end
    if(1'h0) begin
    end else begin
      useRAS_30 <= GEN_291;
    end
    if(1'h0) begin
    end else begin
      useRAS_31 <= GEN_292;
    end
    if(1'h0) begin
    end else begin
      useRAS_32 <= GEN_293;
    end
    if(1'h0) begin
    end else begin
      useRAS_33 <= GEN_294;
    end
    if(1'h0) begin
    end else begin
      useRAS_34 <= GEN_295;
    end
    if(1'h0) begin
    end else begin
      useRAS_35 <= GEN_296;
    end
    if(1'h0) begin
    end else begin
      useRAS_36 <= GEN_297;
    end
    if(1'h0) begin
    end else begin
      useRAS_37 <= GEN_298;
    end
    if(1'h0) begin
    end else begin
      useRAS_38 <= GEN_299;
    end
    if(1'h0) begin
    end else begin
      useRAS_39 <= GEN_300;
    end
    if(1'h0) begin
    end else begin
      useRAS_40 <= GEN_301;
    end
    if(1'h0) begin
    end else begin
      useRAS_41 <= GEN_302;
    end
    if(1'h0) begin
    end else begin
      useRAS_42 <= GEN_303;
    end
    if(1'h0) begin
    end else begin
      useRAS_43 <= GEN_304;
    end
    if(1'h0) begin
    end else begin
      useRAS_44 <= GEN_305;
    end
    if(1'h0) begin
    end else begin
      useRAS_45 <= GEN_306;
    end
    if(1'h0) begin
    end else begin
      useRAS_46 <= GEN_307;
    end
    if(1'h0) begin
    end else begin
      useRAS_47 <= GEN_308;
    end
    if(1'h0) begin
    end else begin
      useRAS_48 <= GEN_309;
    end
    if(1'h0) begin
    end else begin
      useRAS_49 <= GEN_310;
    end
    if(1'h0) begin
    end else begin
      useRAS_50 <= GEN_311;
    end
    if(1'h0) begin
    end else begin
      useRAS_51 <= GEN_312;
    end
    if(1'h0) begin
    end else begin
      useRAS_52 <= GEN_313;
    end
    if(1'h0) begin
    end else begin
      useRAS_53 <= GEN_314;
    end
    if(1'h0) begin
    end else begin
      useRAS_54 <= GEN_315;
    end
    if(1'h0) begin
    end else begin
      useRAS_55 <= GEN_316;
    end
    if(1'h0) begin
    end else begin
      useRAS_56 <= GEN_317;
    end
    if(1'h0) begin
    end else begin
      useRAS_57 <= GEN_318;
    end
    if(1'h0) begin
    end else begin
      useRAS_58 <= GEN_319;
    end
    if(1'h0) begin
    end else begin
      useRAS_59 <= GEN_320;
    end
    if(1'h0) begin
    end else begin
      useRAS_60 <= GEN_321;
    end
    if(1'h0) begin
    end else begin
      useRAS_61 <= GEN_322;
    end
    if(1'h0) begin
    end else begin
      isJump_0 <= GEN_324;
    end
    if(1'h0) begin
    end else begin
      isJump_1 <= GEN_325;
    end
    if(1'h0) begin
    end else begin
      isJump_2 <= GEN_326;
    end
    if(1'h0) begin
    end else begin
      isJump_3 <= GEN_327;
    end
    if(1'h0) begin
    end else begin
      isJump_4 <= GEN_328;
    end
    if(1'h0) begin
    end else begin
      isJump_5 <= GEN_329;
    end
    if(1'h0) begin
    end else begin
      isJump_6 <= GEN_330;
    end
    if(1'h0) begin
    end else begin
      isJump_7 <= GEN_331;
    end
    if(1'h0) begin
    end else begin
      isJump_8 <= GEN_332;
    end
    if(1'h0) begin
    end else begin
      isJump_9 <= GEN_333;
    end
    if(1'h0) begin
    end else begin
      isJump_10 <= GEN_334;
    end
    if(1'h0) begin
    end else begin
      isJump_11 <= GEN_335;
    end
    if(1'h0) begin
    end else begin
      isJump_12 <= GEN_336;
    end
    if(1'h0) begin
    end else begin
      isJump_13 <= GEN_337;
    end
    if(1'h0) begin
    end else begin
      isJump_14 <= GEN_338;
    end
    if(1'h0) begin
    end else begin
      isJump_15 <= GEN_339;
    end
    if(1'h0) begin
    end else begin
      isJump_16 <= GEN_340;
    end
    if(1'h0) begin
    end else begin
      isJump_17 <= GEN_341;
    end
    if(1'h0) begin
    end else begin
      isJump_18 <= GEN_342;
    end
    if(1'h0) begin
    end else begin
      isJump_19 <= GEN_343;
    end
    if(1'h0) begin
    end else begin
      isJump_20 <= GEN_344;
    end
    if(1'h0) begin
    end else begin
      isJump_21 <= GEN_345;
    end
    if(1'h0) begin
    end else begin
      isJump_22 <= GEN_346;
    end
    if(1'h0) begin
    end else begin
      isJump_23 <= GEN_347;
    end
    if(1'h0) begin
    end else begin
      isJump_24 <= GEN_348;
    end
    if(1'h0) begin
    end else begin
      isJump_25 <= GEN_349;
    end
    if(1'h0) begin
    end else begin
      isJump_26 <= GEN_350;
    end
    if(1'h0) begin
    end else begin
      isJump_27 <= GEN_351;
    end
    if(1'h0) begin
    end else begin
      isJump_28 <= GEN_352;
    end
    if(1'h0) begin
    end else begin
      isJump_29 <= GEN_353;
    end
    if(1'h0) begin
    end else begin
      isJump_30 <= GEN_354;
    end
    if(1'h0) begin
    end else begin
      isJump_31 <= GEN_355;
    end
    if(1'h0) begin
    end else begin
      isJump_32 <= GEN_356;
    end
    if(1'h0) begin
    end else begin
      isJump_33 <= GEN_357;
    end
    if(1'h0) begin
    end else begin
      isJump_34 <= GEN_358;
    end
    if(1'h0) begin
    end else begin
      isJump_35 <= GEN_359;
    end
    if(1'h0) begin
    end else begin
      isJump_36 <= GEN_360;
    end
    if(1'h0) begin
    end else begin
      isJump_37 <= GEN_361;
    end
    if(1'h0) begin
    end else begin
      isJump_38 <= GEN_362;
    end
    if(1'h0) begin
    end else begin
      isJump_39 <= GEN_363;
    end
    if(1'h0) begin
    end else begin
      isJump_40 <= GEN_364;
    end
    if(1'h0) begin
    end else begin
      isJump_41 <= GEN_365;
    end
    if(1'h0) begin
    end else begin
      isJump_42 <= GEN_366;
    end
    if(1'h0) begin
    end else begin
      isJump_43 <= GEN_367;
    end
    if(1'h0) begin
    end else begin
      isJump_44 <= GEN_368;
    end
    if(1'h0) begin
    end else begin
      isJump_45 <= GEN_369;
    end
    if(1'h0) begin
    end else begin
      isJump_46 <= GEN_370;
    end
    if(1'h0) begin
    end else begin
      isJump_47 <= GEN_371;
    end
    if(1'h0) begin
    end else begin
      isJump_48 <= GEN_372;
    end
    if(1'h0) begin
    end else begin
      isJump_49 <= GEN_373;
    end
    if(1'h0) begin
    end else begin
      isJump_50 <= GEN_374;
    end
    if(1'h0) begin
    end else begin
      isJump_51 <= GEN_375;
    end
    if(1'h0) begin
    end else begin
      isJump_52 <= GEN_376;
    end
    if(1'h0) begin
    end else begin
      isJump_53 <= GEN_377;
    end
    if(1'h0) begin
    end else begin
      isJump_54 <= GEN_378;
    end
    if(1'h0) begin
    end else begin
      isJump_55 <= GEN_379;
    end
    if(1'h0) begin
    end else begin
      isJump_56 <= GEN_380;
    end
    if(1'h0) begin
    end else begin
      isJump_57 <= GEN_381;
    end
    if(1'h0) begin
    end else begin
      isJump_58 <= GEN_382;
    end
    if(1'h0) begin
    end else begin
      isJump_59 <= GEN_383;
    end
    if(1'h0) begin
    end else begin
      isJump_60 <= GEN_384;
    end
    if(1'h0) begin
    end else begin
      isJump_61 <= GEN_385;
    end
    if(brIdx_T_2876_en & brIdx_T_2876_mask) begin
      brIdx[brIdx_T_2876_addr] <= brIdx_T_2876_data;
    end
    if(reset) begin
      T_1215 <= 1'h0;
    end else begin
      T_1215 <= io_btb_update_valid;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_valid <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_taken <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_mask <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_bridx <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_target <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_entry <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_bht_history <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      T_1216_prediction_bits_bht_value <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      T_1216_pc <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      T_1216_target <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      T_1216_taken <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      T_1216_isJump <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_1216_isReturn <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      T_1216_br_pc <= GEN_17;
    end
    if(reset) begin
      nextRepl <= 6'h0;
    end else begin
      nextRepl <= GEN_19;
    end
    if(reset) begin
      T_2536 <= 3'h0;
    end else begin
      T_2536 <= GEN_21;
    end
    if(T_3616_T_3949_en & T_3616_T_3949_mask) begin
      T_3616[T_3616_T_3949_addr] <= T_3616_T_3949_data;
    end
    if(1'h0) begin
    end else begin
      T_3618 <= GEN_431;
    end
    if(reset) begin
      T_3967 <= 2'h0;
    end else begin
      T_3967 <= GEN_456;
    end
    if(reset) begin
      T_3969 <= 1'h0;
    end else begin
      T_3969 <= GEN_454;
    end
    if(1'h0) begin
    end else begin
      T_3976_0 <= GEN_452;
    end
    if(1'h0) begin
    end else begin
      T_3976_1 <= GEN_453;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (r_btb_update_valid & T_2549) begin
          $fwrite(32'h80000002,"Assertion failed: BTB request != I$ target\n    at btb.scala:202 assert(io.req.bits.addr === r_btb_update.bits.target, \"BTB request != I$ target\")\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (r_btb_update_valid & T_2549) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module Queue_66(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [31:0] io_enq_bits_data,
  input  [63:0] io_enq_bits_datablock,
  input   io_deq_ready,
  output  io_deq_valid,
  output [31:0] io_deq_bits_data,
  output [63:0] io_deq_bits_datablock,
  output  io_count
);
  reg [31:0] ram_data [0:0];
  reg [31:0] GEN_0;
  wire [31:0] ram_data_T_744_data;
  wire  ram_data_T_744_addr;
  wire  ram_data_T_744_en;
  wire [31:0] ram_data_T_665_data;
  wire  ram_data_T_665_addr;
  wire  ram_data_T_665_mask;
  wire  ram_data_T_665_en;
  reg [63:0] ram_datablock [0:0];
  reg [63:0] GEN_1;
  wire [63:0] ram_datablock_T_744_data;
  wire  ram_datablock_T_744_addr;
  wire  ram_datablock_T_744_en;
  wire [63:0] ram_datablock_T_665_data;
  wire  ram_datablock_T_665_addr;
  wire  ram_datablock_T_665_mask;
  wire  ram_datablock_T_665_en;
  reg  maybe_full;
  reg [31:0] GEN_2;
  wire  T_662;
  wire  T_663;
  wire  do_enq;
  wire  T_664;
  wire  do_deq;
  wire  T_739;
  wire  GEN_7;
  wire  T_741;
  wire  GEN_8;
  wire [1:0] T_817;
  wire  ptr_diff;
  wire [1:0] T_819;
  assign io_enq_ready = GEN_8;
  assign io_deq_valid = T_741;
  assign io_deq_bits_data = ram_data_T_744_data;
  assign io_deq_bits_datablock = ram_datablock_T_744_data;
  assign io_count = T_819[0];
  assign ram_data_T_744_addr = 1'h0;
  assign ram_data_T_744_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_data_T_744_data = ram_data[ram_data_T_744_addr];
  `else
  assign ram_data_T_744_data = ram_data_T_744_addr >= 1'h1 ? $random : ram_data[ram_data_T_744_addr];
  `endif
  assign ram_data_T_665_data = io_enq_bits_data;
  assign ram_data_T_665_addr = 1'h0;
  assign ram_data_T_665_mask = do_enq;
  assign ram_data_T_665_en = do_enq;
  assign ram_datablock_T_744_addr = 1'h0;
  assign ram_datablock_T_744_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_datablock_T_744_data = ram_datablock[ram_datablock_T_744_addr];
  `else
  assign ram_datablock_T_744_data = ram_datablock_T_744_addr >= 1'h1 ? $random : ram_datablock[ram_datablock_T_744_addr];
  `endif
  assign ram_datablock_T_665_data = io_enq_bits_datablock;
  assign ram_datablock_T_665_addr = 1'h0;
  assign ram_datablock_T_665_mask = do_enq;
  assign ram_datablock_T_665_en = do_enq;
  assign T_662 = maybe_full == 1'h0;
  assign T_663 = io_enq_ready & io_enq_valid;
  assign do_enq = T_663;
  assign T_664 = io_deq_ready & io_deq_valid;
  assign do_deq = T_664;
  assign T_739 = do_enq != do_deq;
  assign GEN_7 = T_739 ? do_enq : maybe_full;
  assign T_741 = T_662 == 1'h0;
  assign GEN_8 = io_deq_ready ? 1'h1 : T_662;
  assign T_817 = 1'h0 - 1'h0;
  assign ptr_diff = T_817[0:0];
  assign T_819 = {maybe_full,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_data[initvar] = GEN_0[31:0];
  GEN_1 = {2{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_datablock[initvar] = GEN_1[63:0];
  GEN_2 = {1{$random}};
  maybe_full = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_data_T_665_en & ram_data_T_665_mask) begin
      ram_data[ram_data_T_665_addr] <= ram_data_T_665_data;
    end
    if(ram_datablock_T_665_en & ram_datablock_T_665_mask) begin
      ram_datablock[ram_datablock_T_665_addr] <= ram_datablock_T_665_data;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_7;
    end
  end
endmodule
module Frontend(
  input   clk,
  input   reset,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_pc,
  input   io_cpu_resp_ready,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_data_0,
  output  io_cpu_resp_bits_mask,
  output  io_cpu_resp_bits_xcpt_if,
  output  io_cpu_btb_resp_valid,
  output  io_cpu_btb_resp_bits_taken,
  output  io_cpu_btb_resp_bits_mask,
  output  io_cpu_btb_resp_bits_bridx,
  output [38:0] io_cpu_btb_resp_bits_target,
  output [5:0] io_cpu_btb_resp_bits_entry,
  output [6:0] io_cpu_btb_resp_bits_bht_history,
  output [1:0] io_cpu_btb_resp_bits_bht_value,
  input   io_cpu_btb_update_valid,
  input   io_cpu_btb_update_bits_prediction_valid,
  input   io_cpu_btb_update_bits_prediction_bits_taken,
  input   io_cpu_btb_update_bits_prediction_bits_mask,
  input   io_cpu_btb_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_btb_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_btb_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_btb_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_btb_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_btb_update_bits_pc,
  input  [38:0] io_cpu_btb_update_bits_target,
  input   io_cpu_btb_update_bits_taken,
  input   io_cpu_btb_update_bits_isJump,
  input   io_cpu_btb_update_bits_isReturn,
  input  [38:0] io_cpu_btb_update_bits_br_pc,
  input   io_cpu_bht_update_valid,
  input   io_cpu_bht_update_bits_prediction_valid,
  input   io_cpu_bht_update_bits_prediction_bits_taken,
  input   io_cpu_bht_update_bits_prediction_bits_mask,
  input   io_cpu_bht_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_bht_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_bht_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_bht_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_bht_update_bits_prediction_bits_bht_value,
  input  [38:0] io_cpu_bht_update_bits_pc,
  input   io_cpu_bht_update_bits_taken,
  input   io_cpu_bht_update_bits_mispredict,
  input   io_cpu_ras_update_valid,
  input   io_cpu_ras_update_bits_isCall,
  input   io_cpu_ras_update_bits_isReturn,
  input  [38:0] io_cpu_ras_update_bits_returnAddr,
  input   io_cpu_ras_update_bits_prediction_valid,
  input   io_cpu_ras_update_bits_prediction_bits_taken,
  input   io_cpu_ras_update_bits_prediction_bits_mask,
  input   io_cpu_ras_update_bits_prediction_bits_bridx,
  input  [38:0] io_cpu_ras_update_bits_prediction_bits_target,
  input  [5:0] io_cpu_ras_update_bits_prediction_bits_entry,
  input  [6:0] io_cpu_ras_update_bits_prediction_bits_bht_history,
  input  [1:0] io_cpu_ras_update_bits_prediction_bits_bht_value,
  input   io_cpu_flush_icache,
  input   io_cpu_flush_tlb,
  output [39:0] io_cpu_npc,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_ptw_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data
);
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_req_valid;
  wire [38:0] icache_io_req_bits_addr;
  wire [19:0] icache_io_s1_ppn;
  wire  icache_io_s1_kill;
  wire  icache_io_resp_ready;
  wire  icache_io_resp_valid;
  wire [31:0] icache_io_resp_bits_data;
  wire [63:0] icache_io_resp_bits_datablock;
  wire  icache_io_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  tlb_clk;
  wire  tlb_reset;
  wire  tlb_io_req_ready;
  wire  tlb_io_req_valid;
  wire [6:0] tlb_io_req_bits_asid;
  wire [27:0] tlb_io_req_bits_vpn;
  wire  tlb_io_req_bits_passthrough;
  wire  tlb_io_req_bits_instruction;
  wire  tlb_io_req_bits_store;
  wire  tlb_io_resp_miss;
  wire [19:0] tlb_io_resp_ppn;
  wire  tlb_io_resp_xcpt_ld;
  wire  tlb_io_resp_xcpt_st;
  wire  tlb_io_resp_xcpt_if;
  wire [7:0] tlb_io_resp_hit_idx;
  wire  tlb_io_ptw_req_ready;
  wire  tlb_io_ptw_req_valid;
  wire [26:0] tlb_io_ptw_req_bits_addr;
  wire [1:0] tlb_io_ptw_req_bits_prv;
  wire  tlb_io_ptw_req_bits_store;
  wire  tlb_io_ptw_req_bits_fetch;
  wire  tlb_io_ptw_resp_valid;
  wire [19:0] tlb_io_ptw_resp_bits_pte_ppn;
  wire [2:0] tlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  tlb_io_ptw_resp_bits_pte_d;
  wire  tlb_io_ptw_resp_bits_pte_r;
  wire [3:0] tlb_io_ptw_resp_bits_pte_typ;
  wire  tlb_io_ptw_resp_bits_pte_v;
  wire  tlb_io_ptw_status_debug;
  wire [1:0] tlb_io_ptw_status_prv;
  wire  tlb_io_ptw_status_sd;
  wire [30:0] tlb_io_ptw_status_zero3;
  wire  tlb_io_ptw_status_sd_rv32;
  wire [1:0] tlb_io_ptw_status_zero2;
  wire [4:0] tlb_io_ptw_status_vm;
  wire [4:0] tlb_io_ptw_status_zero1;
  wire  tlb_io_ptw_status_pum;
  wire  tlb_io_ptw_status_mprv;
  wire [1:0] tlb_io_ptw_status_xs;
  wire [1:0] tlb_io_ptw_status_fs;
  wire [1:0] tlb_io_ptw_status_mpp;
  wire [1:0] tlb_io_ptw_status_hpp;
  wire  tlb_io_ptw_status_spp;
  wire  tlb_io_ptw_status_mpie;
  wire  tlb_io_ptw_status_hpie;
  wire  tlb_io_ptw_status_spie;
  wire  tlb_io_ptw_status_upie;
  wire  tlb_io_ptw_status_mie;
  wire  tlb_io_ptw_status_hie;
  wire  tlb_io_ptw_status_sie;
  wire  tlb_io_ptw_status_uie;
  wire  tlb_io_ptw_invalidate;
  reg [39:0] s1_pc_;
  reg [63:0] GEN_10;
  wire [39:0] T_1296;
  wire [39:0] GEN_21;
  wire [39:0] T_1298;
  wire [39:0] s1_pc;
  reg  s1_same_block;
  reg [31:0] GEN_22;
  reg  s2_valid;
  reg [31:0] GEN_28;
  reg [39:0] s2_pc;
  reg [63:0] GEN_29;
  reg  s2_btb_resp_valid;
  reg [31:0] GEN_30;
  reg  s2_btb_resp_bits_taken;
  reg [31:0] GEN_31;
  reg  s2_btb_resp_bits_mask;
  reg [31:0] GEN_32;
  reg  s2_btb_resp_bits_bridx;
  reg [31:0] GEN_33;
  reg [38:0] s2_btb_resp_bits_target;
  reg [63:0] GEN_34;
  reg [5:0] s2_btb_resp_bits_entry;
  reg [31:0] GEN_35;
  reg [6:0] s2_btb_resp_bits_bht_history;
  reg [31:0] GEN_36;
  reg [1:0] s2_btb_resp_bits_bht_value;
  reg [31:0] GEN_37;
  reg  s2_xcpt_if;
  reg [31:0] GEN_38;
  wire  s2_resp_valid;
  wire [63:0] s2_resp_data;
  wire [39:0] T_1323;
  wire [39:0] T_1325;
  wire [39:0] T_1326;
  wire [39:0] GEN_23;
  wire [40:0] T_1328;
  wire [39:0] ntpc_0;
  wire  T_1329;
  wire  T_1330;
  wire  T_1331;
  wire [40:0] ntpc;
  wire [40:0] predicted_npc;
  wire  T_1333;
  wire  icmiss;
  wire [40:0] npc;
  wire  T_1335;
  wire  T_1337;
  wire  T_1338;
  wire [40:0] GEN_24;
  wire [40:0] T_1340;
  wire [39:0] GEN_25;
  wire [39:0] T_1342;
  wire [40:0] GEN_26;
  wire  T_1343;
  wire  T_1344;
  wire  s0_same_block;
  wire  T_1346;
  wire  stall;
  wire  T_1348;
  wire  T_1350;
  wire  T_1351;
  wire [39:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire [40:0] GEN_3;
  wire  GEN_4;
  wire [39:0] GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire [40:0] GEN_8;
  wire  GEN_9;
  wire  BTB_1358_clk;
  wire  BTB_1358_reset;
  wire  BTB_1358_io_req_valid;
  wire [38:0] BTB_1358_io_req_bits_addr;
  wire  BTB_1358_io_resp_valid;
  wire  BTB_1358_io_resp_bits_taken;
  wire  BTB_1358_io_resp_bits_mask;
  wire  BTB_1358_io_resp_bits_bridx;
  wire [38:0] BTB_1358_io_resp_bits_target;
  wire [5:0] BTB_1358_io_resp_bits_entry;
  wire [6:0] BTB_1358_io_resp_bits_bht_history;
  wire [1:0] BTB_1358_io_resp_bits_bht_value;
  wire  BTB_1358_io_btb_update_valid;
  wire  BTB_1358_io_btb_update_bits_prediction_valid;
  wire  BTB_1358_io_btb_update_bits_prediction_bits_taken;
  wire  BTB_1358_io_btb_update_bits_prediction_bits_mask;
  wire  BTB_1358_io_btb_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1358_io_btb_update_bits_prediction_bits_target;
  wire [5:0] BTB_1358_io_btb_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1358_io_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1358_io_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1358_io_btb_update_bits_pc;
  wire [38:0] BTB_1358_io_btb_update_bits_target;
  wire  BTB_1358_io_btb_update_bits_taken;
  wire  BTB_1358_io_btb_update_bits_isJump;
  wire  BTB_1358_io_btb_update_bits_isReturn;
  wire [38:0] BTB_1358_io_btb_update_bits_br_pc;
  wire  BTB_1358_io_bht_update_valid;
  wire  BTB_1358_io_bht_update_bits_prediction_valid;
  wire  BTB_1358_io_bht_update_bits_prediction_bits_taken;
  wire  BTB_1358_io_bht_update_bits_prediction_bits_mask;
  wire  BTB_1358_io_bht_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1358_io_bht_update_bits_prediction_bits_target;
  wire [5:0] BTB_1358_io_bht_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1358_io_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1358_io_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] BTB_1358_io_bht_update_bits_pc;
  wire  BTB_1358_io_bht_update_bits_taken;
  wire  BTB_1358_io_bht_update_bits_mispredict;
  wire  BTB_1358_io_ras_update_valid;
  wire  BTB_1358_io_ras_update_bits_isCall;
  wire  BTB_1358_io_ras_update_bits_isReturn;
  wire [38:0] BTB_1358_io_ras_update_bits_returnAddr;
  wire  BTB_1358_io_ras_update_bits_prediction_valid;
  wire  BTB_1358_io_ras_update_bits_prediction_bits_taken;
  wire  BTB_1358_io_ras_update_bits_prediction_bits_mask;
  wire  BTB_1358_io_ras_update_bits_prediction_bits_bridx;
  wire [38:0] BTB_1358_io_ras_update_bits_prediction_bits_target;
  wire [5:0] BTB_1358_io_ras_update_bits_prediction_bits_entry;
  wire [6:0] BTB_1358_io_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] BTB_1358_io_ras_update_bits_prediction_bits_bht_value;
  wire  BTB_1358_io_invalidate;
  wire  T_1360;
  wire  T_1365;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire [38:0] GEN_15;
  wire [5:0] GEN_16;
  wire [6:0] GEN_17;
  wire [1:0] GEN_18;
  wire  T_1367;
  wire [39:0] T_1368;
  wire [40:0] GEN_19;
  wire  GEN_20;
  wire [27:0] T_1375;
  wire  T_1383;
  wire  T_1384;
  wire  T_1385;
  wire  T_1386;
  wire  T_1387;
  wire  T_1388;
  wire  T_1389;
  wire  T_1390;
  wire [40:0] T_1391;
  wire  Queue_66_1464_clk;
  wire  Queue_66_1464_reset;
  wire  Queue_66_1464_io_enq_ready;
  wire  Queue_66_1464_io_enq_valid;
  wire [31:0] Queue_66_1464_io_enq_bits_data;
  wire [63:0] Queue_66_1464_io_enq_bits_datablock;
  wire  Queue_66_1464_io_deq_ready;
  wire  Queue_66_1464_io_deq_valid;
  wire [31:0] Queue_66_1464_io_deq_bits_data;
  wire [63:0] Queue_66_1464_io_deq_bits_datablock;
  wire  Queue_66_1464_io_count;
  wire  T_1468;
  wire  T_1469;
  wire  T_1470;
  wire [5:0] GEN_27;
  wire [5:0] T_1471;
  wire [63:0] fetch_data;
  wire [31:0] T_1472;
  ICache icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_req_valid(icache_io_req_valid),
    .io_req_bits_addr(icache_io_req_bits_addr),
    .io_s1_ppn(icache_io_s1_ppn),
    .io_s1_kill(icache_io_s1_kill),
    .io_resp_ready(icache_io_resp_ready),
    .io_resp_valid(icache_io_resp_valid),
    .io_resp_bits_data(icache_io_resp_bits_data),
    .io_resp_bits_datablock(icache_io_resp_bits_datablock),
    .io_invalidate(icache_io_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  TLB tlb (
    .clk(tlb_clk),
    .reset(tlb_reset),
    .io_req_ready(tlb_io_req_ready),
    .io_req_valid(tlb_io_req_valid),
    .io_req_bits_asid(tlb_io_req_bits_asid),
    .io_req_bits_vpn(tlb_io_req_bits_vpn),
    .io_req_bits_passthrough(tlb_io_req_bits_passthrough),
    .io_req_bits_instruction(tlb_io_req_bits_instruction),
    .io_req_bits_store(tlb_io_req_bits_store),
    .io_resp_miss(tlb_io_resp_miss),
    .io_resp_ppn(tlb_io_resp_ppn),
    .io_resp_xcpt_ld(tlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(tlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(tlb_io_resp_xcpt_if),
    .io_resp_hit_idx(tlb_io_resp_hit_idx),
    .io_ptw_req_ready(tlb_io_ptw_req_ready),
    .io_ptw_req_valid(tlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(tlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(tlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(tlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(tlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(tlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(tlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(tlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(tlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(tlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(tlb_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(tlb_io_ptw_resp_bits_pte_v),
    .io_ptw_status_debug(tlb_io_ptw_status_debug),
    .io_ptw_status_prv(tlb_io_ptw_status_prv),
    .io_ptw_status_sd(tlb_io_ptw_status_sd),
    .io_ptw_status_zero3(tlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(tlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(tlb_io_ptw_status_zero2),
    .io_ptw_status_vm(tlb_io_ptw_status_vm),
    .io_ptw_status_zero1(tlb_io_ptw_status_zero1),
    .io_ptw_status_pum(tlb_io_ptw_status_pum),
    .io_ptw_status_mprv(tlb_io_ptw_status_mprv),
    .io_ptw_status_xs(tlb_io_ptw_status_xs),
    .io_ptw_status_fs(tlb_io_ptw_status_fs),
    .io_ptw_status_mpp(tlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(tlb_io_ptw_status_hpp),
    .io_ptw_status_spp(tlb_io_ptw_status_spp),
    .io_ptw_status_mpie(tlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(tlb_io_ptw_status_hpie),
    .io_ptw_status_spie(tlb_io_ptw_status_spie),
    .io_ptw_status_upie(tlb_io_ptw_status_upie),
    .io_ptw_status_mie(tlb_io_ptw_status_mie),
    .io_ptw_status_hie(tlb_io_ptw_status_hie),
    .io_ptw_status_sie(tlb_io_ptw_status_sie),
    .io_ptw_status_uie(tlb_io_ptw_status_uie),
    .io_ptw_invalidate(tlb_io_ptw_invalidate)
  );
  BTB BTB_1358 (
    .clk(BTB_1358_clk),
    .reset(BTB_1358_reset),
    .io_req_valid(BTB_1358_io_req_valid),
    .io_req_bits_addr(BTB_1358_io_req_bits_addr),
    .io_resp_valid(BTB_1358_io_resp_valid),
    .io_resp_bits_taken(BTB_1358_io_resp_bits_taken),
    .io_resp_bits_mask(BTB_1358_io_resp_bits_mask),
    .io_resp_bits_bridx(BTB_1358_io_resp_bits_bridx),
    .io_resp_bits_target(BTB_1358_io_resp_bits_target),
    .io_resp_bits_entry(BTB_1358_io_resp_bits_entry),
    .io_resp_bits_bht_history(BTB_1358_io_resp_bits_bht_history),
    .io_resp_bits_bht_value(BTB_1358_io_resp_bits_bht_value),
    .io_btb_update_valid(BTB_1358_io_btb_update_valid),
    .io_btb_update_bits_prediction_valid(BTB_1358_io_btb_update_bits_prediction_valid),
    .io_btb_update_bits_prediction_bits_taken(BTB_1358_io_btb_update_bits_prediction_bits_taken),
    .io_btb_update_bits_prediction_bits_mask(BTB_1358_io_btb_update_bits_prediction_bits_mask),
    .io_btb_update_bits_prediction_bits_bridx(BTB_1358_io_btb_update_bits_prediction_bits_bridx),
    .io_btb_update_bits_prediction_bits_target(BTB_1358_io_btb_update_bits_prediction_bits_target),
    .io_btb_update_bits_prediction_bits_entry(BTB_1358_io_btb_update_bits_prediction_bits_entry),
    .io_btb_update_bits_prediction_bits_bht_history(BTB_1358_io_btb_update_bits_prediction_bits_bht_history),
    .io_btb_update_bits_prediction_bits_bht_value(BTB_1358_io_btb_update_bits_prediction_bits_bht_value),
    .io_btb_update_bits_pc(BTB_1358_io_btb_update_bits_pc),
    .io_btb_update_bits_target(BTB_1358_io_btb_update_bits_target),
    .io_btb_update_bits_taken(BTB_1358_io_btb_update_bits_taken),
    .io_btb_update_bits_isJump(BTB_1358_io_btb_update_bits_isJump),
    .io_btb_update_bits_isReturn(BTB_1358_io_btb_update_bits_isReturn),
    .io_btb_update_bits_br_pc(BTB_1358_io_btb_update_bits_br_pc),
    .io_bht_update_valid(BTB_1358_io_bht_update_valid),
    .io_bht_update_bits_prediction_valid(BTB_1358_io_bht_update_bits_prediction_valid),
    .io_bht_update_bits_prediction_bits_taken(BTB_1358_io_bht_update_bits_prediction_bits_taken),
    .io_bht_update_bits_prediction_bits_mask(BTB_1358_io_bht_update_bits_prediction_bits_mask),
    .io_bht_update_bits_prediction_bits_bridx(BTB_1358_io_bht_update_bits_prediction_bits_bridx),
    .io_bht_update_bits_prediction_bits_target(BTB_1358_io_bht_update_bits_prediction_bits_target),
    .io_bht_update_bits_prediction_bits_entry(BTB_1358_io_bht_update_bits_prediction_bits_entry),
    .io_bht_update_bits_prediction_bits_bht_history(BTB_1358_io_bht_update_bits_prediction_bits_bht_history),
    .io_bht_update_bits_prediction_bits_bht_value(BTB_1358_io_bht_update_bits_prediction_bits_bht_value),
    .io_bht_update_bits_pc(BTB_1358_io_bht_update_bits_pc),
    .io_bht_update_bits_taken(BTB_1358_io_bht_update_bits_taken),
    .io_bht_update_bits_mispredict(BTB_1358_io_bht_update_bits_mispredict),
    .io_ras_update_valid(BTB_1358_io_ras_update_valid),
    .io_ras_update_bits_isCall(BTB_1358_io_ras_update_bits_isCall),
    .io_ras_update_bits_isReturn(BTB_1358_io_ras_update_bits_isReturn),
    .io_ras_update_bits_returnAddr(BTB_1358_io_ras_update_bits_returnAddr),
    .io_ras_update_bits_prediction_valid(BTB_1358_io_ras_update_bits_prediction_valid),
    .io_ras_update_bits_prediction_bits_taken(BTB_1358_io_ras_update_bits_prediction_bits_taken),
    .io_ras_update_bits_prediction_bits_mask(BTB_1358_io_ras_update_bits_prediction_bits_mask),
    .io_ras_update_bits_prediction_bits_bridx(BTB_1358_io_ras_update_bits_prediction_bits_bridx),
    .io_ras_update_bits_prediction_bits_target(BTB_1358_io_ras_update_bits_prediction_bits_target),
    .io_ras_update_bits_prediction_bits_entry(BTB_1358_io_ras_update_bits_prediction_bits_entry),
    .io_ras_update_bits_prediction_bits_bht_history(BTB_1358_io_ras_update_bits_prediction_bits_bht_history),
    .io_ras_update_bits_prediction_bits_bht_value(BTB_1358_io_ras_update_bits_prediction_bits_bht_value),
    .io_invalidate(BTB_1358_io_invalidate)
  );
  Queue_66 Queue_66_1464 (
    .clk(Queue_66_1464_clk),
    .reset(Queue_66_1464_reset),
    .io_enq_ready(Queue_66_1464_io_enq_ready),
    .io_enq_valid(Queue_66_1464_io_enq_valid),
    .io_enq_bits_data(Queue_66_1464_io_enq_bits_data),
    .io_enq_bits_datablock(Queue_66_1464_io_enq_bits_datablock),
    .io_deq_ready(Queue_66_1464_io_deq_ready),
    .io_deq_valid(Queue_66_1464_io_deq_valid),
    .io_deq_bits_data(Queue_66_1464_io_deq_bits_data),
    .io_deq_bits_datablock(Queue_66_1464_io_deq_bits_datablock),
    .io_count(Queue_66_1464_io_count)
  );
  assign io_cpu_resp_valid = T_1390;
  assign io_cpu_resp_bits_pc = s2_pc;
  assign io_cpu_resp_bits_data_0 = T_1472;
  assign io_cpu_resp_bits_mask = 1'h1;
  assign io_cpu_resp_bits_xcpt_if = s2_xcpt_if;
  assign io_cpu_btb_resp_valid = s2_btb_resp_valid;
  assign io_cpu_btb_resp_bits_taken = s2_btb_resp_bits_taken;
  assign io_cpu_btb_resp_bits_mask = s2_btb_resp_bits_mask;
  assign io_cpu_btb_resp_bits_bridx = s2_btb_resp_bits_bridx;
  assign io_cpu_btb_resp_bits_target = s2_btb_resp_bits_target;
  assign io_cpu_btb_resp_bits_entry = s2_btb_resp_bits_entry;
  assign io_cpu_btb_resp_bits_bht_history = s2_btb_resp_bits_bht_history;
  assign io_cpu_btb_resp_bits_bht_value = s2_btb_resp_bits_bht_value;
  assign io_cpu_npc = T_1391[39:0];
  assign io_ptw_req_valid = tlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = tlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_prv = tlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_store = tlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = tlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = icache_io_mem_acquire_valid;
  assign io_mem_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign io_mem_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign io_mem_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign io_mem_grant_ready = icache_io_mem_grant_ready;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_req_valid = T_1384;
  assign icache_io_req_bits_addr = io_cpu_npc[38:0];
  assign icache_io_s1_ppn = tlb_io_resp_ppn;
  assign icache_io_s1_kill = T_1388;
  assign icache_io_resp_ready = Queue_66_1464_io_enq_ready;
  assign icache_io_invalidate = io_cpu_flush_icache;
  assign icache_io_mem_acquire_ready = io_mem_acquire_ready;
  assign icache_io_mem_grant_valid = io_mem_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign tlb_clk = clk;
  assign tlb_reset = reset;
  assign tlb_io_req_valid = T_1365;
  assign tlb_io_req_bits_asid = {{6'd0}, 1'h0};
  assign tlb_io_req_bits_vpn = T_1375;
  assign tlb_io_req_bits_passthrough = 1'h0;
  assign tlb_io_req_bits_instruction = 1'h1;
  assign tlb_io_req_bits_store = 1'h0;
  assign tlb_io_ptw_req_ready = io_ptw_req_ready;
  assign tlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign tlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign tlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign tlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign tlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign tlb_io_ptw_resp_bits_pte_typ = io_ptw_resp_bits_pte_typ;
  assign tlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign tlb_io_ptw_status_debug = io_ptw_status_debug;
  assign tlb_io_ptw_status_prv = io_ptw_status_prv;
  assign tlb_io_ptw_status_sd = io_ptw_status_sd;
  assign tlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign tlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign tlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign tlb_io_ptw_status_vm = io_ptw_status_vm;
  assign tlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign tlb_io_ptw_status_pum = io_ptw_status_pum;
  assign tlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign tlb_io_ptw_status_xs = io_ptw_status_xs;
  assign tlb_io_ptw_status_fs = io_ptw_status_fs;
  assign tlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign tlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign tlb_io_ptw_status_spp = io_ptw_status_spp;
  assign tlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign tlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign tlb_io_ptw_status_spie = io_ptw_status_spie;
  assign tlb_io_ptw_status_upie = io_ptw_status_upie;
  assign tlb_io_ptw_status_mie = io_ptw_status_mie;
  assign tlb_io_ptw_status_hie = io_ptw_status_hie;
  assign tlb_io_ptw_status_sie = io_ptw_status_sie;
  assign tlb_io_ptw_status_uie = io_ptw_status_uie;
  assign tlb_io_ptw_invalidate = io_ptw_invalidate;
  assign T_1296 = ~ s1_pc_;
  assign GEN_21 = {{38'd0}, 2'h3};
  assign T_1298 = T_1296 | GEN_21;
  assign s1_pc = ~ T_1298;
  assign s2_resp_valid = Queue_66_1464_io_deq_valid;
  assign s2_resp_data = Queue_66_1464_io_deq_bits_datablock;
  assign T_1323 = ~ s1_pc;
  assign T_1325 = T_1323 | GEN_21;
  assign T_1326 = ~ T_1325;
  assign GEN_23 = {{37'd0}, 3'h4};
  assign T_1328 = T_1326 + GEN_23;
  assign ntpc_0 = T_1328[39:0];
  assign T_1329 = s1_pc[38];
  assign T_1330 = ntpc_0[38];
  assign T_1331 = T_1329 & T_1330;
  assign ntpc = {T_1331,ntpc_0};
  assign predicted_npc = GEN_19;
  assign T_1333 = s2_resp_valid == 1'h0;
  assign icmiss = s2_valid & T_1333;
  assign npc = icmiss ? {{1'd0}, s2_pc} : predicted_npc;
  assign T_1335 = icmiss == 1'h0;
  assign T_1337 = io_cpu_req_valid == 1'h0;
  assign T_1338 = T_1335 & T_1337;
  assign GEN_24 = {{37'd0}, 4'h8};
  assign T_1340 = ntpc & GEN_24;
  assign GEN_25 = {{36'd0}, 4'h8};
  assign T_1342 = s1_pc & GEN_25;
  assign GEN_26 = {{1'd0}, T_1342};
  assign T_1343 = T_1340 == GEN_26;
  assign T_1344 = T_1338 & T_1343;
  assign s0_same_block = GEN_20;
  assign T_1346 = io_cpu_resp_ready == 1'h0;
  assign stall = io_cpu_resp_valid & T_1346;
  assign T_1348 = stall == 1'h0;
  assign T_1350 = tlb_io_resp_miss == 1'h0;
  assign T_1351 = s0_same_block & T_1350;
  assign GEN_0 = T_1335 ? s1_pc : s2_pc;
  assign GEN_1 = T_1335 ? tlb_io_resp_xcpt_if : s2_xcpt_if;
  assign GEN_2 = T_1348 ? T_1351 : s1_same_block;
  assign GEN_3 = T_1348 ? npc : {{1'd0}, s1_pc_};
  assign GEN_4 = T_1348 ? T_1335 : s2_valid;
  assign GEN_5 = T_1348 ? GEN_0 : s2_pc;
  assign GEN_6 = T_1348 ? GEN_1 : s2_xcpt_if;
  assign GEN_7 = io_cpu_req_valid ? 1'h0 : GEN_2;
  assign GEN_8 = io_cpu_req_valid ? {{1'd0}, io_cpu_req_bits_pc} : GEN_3;
  assign GEN_9 = io_cpu_req_valid ? 1'h0 : GEN_4;
  assign BTB_1358_clk = clk;
  assign BTB_1358_reset = reset;
  assign BTB_1358_io_req_valid = T_1365;
  assign BTB_1358_io_req_bits_addr = s1_pc[38:0];
  assign BTB_1358_io_btb_update_valid = io_cpu_btb_update_valid;
  assign BTB_1358_io_btb_update_bits_prediction_valid = io_cpu_btb_update_bits_prediction_valid;
  assign BTB_1358_io_btb_update_bits_prediction_bits_taken = io_cpu_btb_update_bits_prediction_bits_taken;
  assign BTB_1358_io_btb_update_bits_prediction_bits_mask = io_cpu_btb_update_bits_prediction_bits_mask;
  assign BTB_1358_io_btb_update_bits_prediction_bits_bridx = io_cpu_btb_update_bits_prediction_bits_bridx;
  assign BTB_1358_io_btb_update_bits_prediction_bits_target = io_cpu_btb_update_bits_prediction_bits_target;
  assign BTB_1358_io_btb_update_bits_prediction_bits_entry = io_cpu_btb_update_bits_prediction_bits_entry;
  assign BTB_1358_io_btb_update_bits_prediction_bits_bht_history = io_cpu_btb_update_bits_prediction_bits_bht_history;
  assign BTB_1358_io_btb_update_bits_prediction_bits_bht_value = io_cpu_btb_update_bits_prediction_bits_bht_value;
  assign BTB_1358_io_btb_update_bits_pc = io_cpu_btb_update_bits_pc;
  assign BTB_1358_io_btb_update_bits_target = io_cpu_btb_update_bits_target;
  assign BTB_1358_io_btb_update_bits_taken = io_cpu_btb_update_bits_taken;
  assign BTB_1358_io_btb_update_bits_isJump = io_cpu_btb_update_bits_isJump;
  assign BTB_1358_io_btb_update_bits_isReturn = io_cpu_btb_update_bits_isReturn;
  assign BTB_1358_io_btb_update_bits_br_pc = io_cpu_btb_update_bits_br_pc;
  assign BTB_1358_io_bht_update_valid = io_cpu_bht_update_valid;
  assign BTB_1358_io_bht_update_bits_prediction_valid = io_cpu_bht_update_bits_prediction_valid;
  assign BTB_1358_io_bht_update_bits_prediction_bits_taken = io_cpu_bht_update_bits_prediction_bits_taken;
  assign BTB_1358_io_bht_update_bits_prediction_bits_mask = io_cpu_bht_update_bits_prediction_bits_mask;
  assign BTB_1358_io_bht_update_bits_prediction_bits_bridx = io_cpu_bht_update_bits_prediction_bits_bridx;
  assign BTB_1358_io_bht_update_bits_prediction_bits_target = io_cpu_bht_update_bits_prediction_bits_target;
  assign BTB_1358_io_bht_update_bits_prediction_bits_entry = io_cpu_bht_update_bits_prediction_bits_entry;
  assign BTB_1358_io_bht_update_bits_prediction_bits_bht_history = io_cpu_bht_update_bits_prediction_bits_bht_history;
  assign BTB_1358_io_bht_update_bits_prediction_bits_bht_value = io_cpu_bht_update_bits_prediction_bits_bht_value;
  assign BTB_1358_io_bht_update_bits_pc = io_cpu_bht_update_bits_pc;
  assign BTB_1358_io_bht_update_bits_taken = io_cpu_bht_update_bits_taken;
  assign BTB_1358_io_bht_update_bits_mispredict = io_cpu_bht_update_bits_mispredict;
  assign BTB_1358_io_ras_update_valid = io_cpu_ras_update_valid;
  assign BTB_1358_io_ras_update_bits_isCall = io_cpu_ras_update_bits_isCall;
  assign BTB_1358_io_ras_update_bits_isReturn = io_cpu_ras_update_bits_isReturn;
  assign BTB_1358_io_ras_update_bits_returnAddr = io_cpu_ras_update_bits_returnAddr;
  assign BTB_1358_io_ras_update_bits_prediction_valid = io_cpu_ras_update_bits_prediction_valid;
  assign BTB_1358_io_ras_update_bits_prediction_bits_taken = io_cpu_ras_update_bits_prediction_bits_taken;
  assign BTB_1358_io_ras_update_bits_prediction_bits_mask = io_cpu_ras_update_bits_prediction_bits_mask;
  assign BTB_1358_io_ras_update_bits_prediction_bits_bridx = io_cpu_ras_update_bits_prediction_bits_bridx;
  assign BTB_1358_io_ras_update_bits_prediction_bits_target = io_cpu_ras_update_bits_prediction_bits_target;
  assign BTB_1358_io_ras_update_bits_prediction_bits_entry = io_cpu_ras_update_bits_prediction_bits_entry;
  assign BTB_1358_io_ras_update_bits_prediction_bits_bht_history = io_cpu_ras_update_bits_prediction_bits_bht_history;
  assign BTB_1358_io_ras_update_bits_prediction_bits_bht_value = io_cpu_ras_update_bits_prediction_bits_bht_value;
  assign BTB_1358_io_invalidate = T_1360;
  assign T_1360 = io_cpu_flush_icache | io_cpu_flush_tlb;
  assign T_1365 = T_1348 & T_1335;
  assign GEN_11 = T_1365 ? BTB_1358_io_resp_valid : s2_btb_resp_valid;
  assign GEN_12 = T_1365 ? BTB_1358_io_resp_bits_taken : s2_btb_resp_bits_taken;
  assign GEN_13 = T_1365 ? BTB_1358_io_resp_bits_mask : s2_btb_resp_bits_mask;
  assign GEN_14 = T_1365 ? BTB_1358_io_resp_bits_bridx : s2_btb_resp_bits_bridx;
  assign GEN_15 = T_1365 ? BTB_1358_io_resp_bits_target : s2_btb_resp_bits_target;
  assign GEN_16 = T_1365 ? BTB_1358_io_resp_bits_entry : s2_btb_resp_bits_entry;
  assign GEN_17 = T_1365 ? BTB_1358_io_resp_bits_bht_history : s2_btb_resp_bits_bht_history;
  assign GEN_18 = T_1365 ? BTB_1358_io_resp_bits_bht_value : s2_btb_resp_bits_bht_value;
  assign T_1367 = BTB_1358_io_resp_bits_target[38];
  assign T_1368 = {T_1367,BTB_1358_io_resp_bits_target};
  assign GEN_19 = BTB_1358_io_resp_bits_taken ? {{1'd0}, T_1368} : ntpc;
  assign GEN_20 = BTB_1358_io_resp_bits_taken ? 1'h0 : T_1344;
  assign T_1375 = s1_pc[39:12];
  assign T_1383 = s0_same_block == 1'h0;
  assign T_1384 = T_1348 & T_1383;
  assign T_1385 = io_cpu_req_valid | tlb_io_resp_miss;
  assign T_1386 = T_1385 | tlb_io_resp_xcpt_if;
  assign T_1387 = T_1386 | icmiss;
  assign T_1388 = T_1387 | io_cpu_flush_tlb;
  assign T_1389 = s2_xcpt_if | s2_resp_valid;
  assign T_1390 = s2_valid & T_1389;
  assign T_1391 = io_cpu_req_valid ? {{1'd0}, io_cpu_req_bits_pc} : npc;
  assign Queue_66_1464_clk = clk;
  assign Queue_66_1464_reset = reset;
  assign Queue_66_1464_io_enq_valid = icache_io_resp_valid;
  assign Queue_66_1464_io_enq_bits_data = icache_io_resp_bits_data;
  assign Queue_66_1464_io_enq_bits_datablock = icache_io_resp_bits_datablock;
  assign Queue_66_1464_io_deq_ready = T_1469;
  assign T_1468 = s1_same_block == 1'h0;
  assign T_1469 = T_1348 & T_1468;
  assign T_1470 = s2_pc[2];
  assign GEN_27 = {{5'd0}, T_1470};
  assign T_1471 = GEN_27 << 5;
  assign fetch_data = s2_resp_data >> T_1471;
  assign T_1472 = fetch_data[31:0];
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_10 = {2{$random}};
  s1_pc_ = GEN_10[39:0];
  GEN_22 = {1{$random}};
  s1_same_block = GEN_22[0:0];
  GEN_28 = {1{$random}};
  s2_valid = GEN_28[0:0];
  GEN_29 = {2{$random}};
  s2_pc = GEN_29[39:0];
  GEN_30 = {1{$random}};
  s2_btb_resp_valid = GEN_30[0:0];
  GEN_31 = {1{$random}};
  s2_btb_resp_bits_taken = GEN_31[0:0];
  GEN_32 = {1{$random}};
  s2_btb_resp_bits_mask = GEN_32[0:0];
  GEN_33 = {1{$random}};
  s2_btb_resp_bits_bridx = GEN_33[0:0];
  GEN_34 = {2{$random}};
  s2_btb_resp_bits_target = GEN_34[38:0];
  GEN_35 = {1{$random}};
  s2_btb_resp_bits_entry = GEN_35[5:0];
  GEN_36 = {1{$random}};
  s2_btb_resp_bits_bht_history = GEN_36[6:0];
  GEN_37 = {1{$random}};
  s2_btb_resp_bits_bht_value = GEN_37[1:0];
  GEN_38 = {1{$random}};
  s2_xcpt_if = GEN_38[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      s1_pc_ <= GEN_8[39:0];
    end
    if(1'h0) begin
    end else begin
      s1_same_block <= GEN_7;
    end
    if(reset) begin
      s2_valid <= 1'h1;
    end else begin
      s2_valid <= GEN_9;
    end
    if(reset) begin
      s2_pc <= {{27'd0}, 13'h1000};
    end else begin
      s2_pc <= GEN_5;
    end
    if(reset) begin
      s2_btb_resp_valid <= 1'h0;
    end else begin
      s2_btb_resp_valid <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_taken <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_mask <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_bridx <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_target <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_entry <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_bht_history <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      s2_btb_resp_bits_bht_value <= GEN_18;
    end
    if(reset) begin
      s2_xcpt_if <= 1'h0;
    end else begin
      s2_xcpt_if <= GEN_6;
    end
  end
endmodule
module WritebackUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [2:0] io_req_bits_addr_beat,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_req_bits_voluntary,
  input  [2:0] io_req_bits_r_type,
  input  [63:0] io_req_bits_data,
  input  [3:0] io_req_bits_way_en,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_data_req_ready,
  output  io_data_req_valid,
  output [3:0] io_data_req_bits_way_en,
  output [11:0] io_data_req_bits_addr,
  input  [63:0] io_data_resp,
  input   io_release_ready,
  output  io_release_valid,
  output [2:0] io_release_bits_addr_beat,
  output [25:0] io_release_bits_addr_block,
  output [1:0] io_release_bits_client_xact_id,
  output  io_release_bits_voluntary,
  output [2:0] io_release_bits_r_type,
  output [63:0] io_release_bits_data
);
  reg  active;
  reg [31:0] GEN_6;
  reg  r1_data_req_fired;
  reg [31:0] GEN_7;
  reg  r2_data_req_fired;
  reg [31:0] GEN_8;
  reg [3:0] data_req_cnt;
  reg [31:0] GEN_10;
  wire  T_748;
  reg [2:0] beat_cnt;
  reg [31:0] GEN_33;
  wire [2:0] GEN_29;
  wire [3:0] T_753;
  wire [2:0] T_754;
  wire [2:0] GEN_0;
  reg [2:0] req_addr_beat;
  reg [31:0] GEN_34;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_35;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_36;
  reg  req_voluntary;
  reg [31:0] GEN_37;
  reg [2:0] req_r_type;
  reg [31:0] GEN_38;
  reg [63:0] req_data;
  reg [63:0] GEN_39;
  reg [3:0] req_way_en;
  reg [31:0] GEN_40;
  wire  T_864;
  wire  T_865;
  wire  T_866;
  wire [3:0] GEN_30;
  wire [4:0] T_869;
  wire [3:0] T_870;
  wire [3:0] GEN_2;
  wire  T_872;
  wire [1:0] T_879;
  wire [3:0] GEN_31;
  wire [4:0] T_880;
  wire [3:0] T_881;
  wire  GEN_3;
  wire  GEN_4;
  wire [3:0] GEN_5;
  wire  T_885;
  wire  T_887;
  wire  T_890;
  wire  GEN_9;
  wire  GEN_11;
  wire  GEN_12;
  wire [3:0] GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [3:0] GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  T_891;
  wire  GEN_20;
  wire [3:0] GEN_21;
  wire [2:0] GEN_22;
  wire [25:0] GEN_23;
  wire [1:0] GEN_24;
  wire  GEN_25;
  wire [2:0] GEN_26;
  wire [63:0] GEN_27;
  wire [3:0] GEN_28;
  wire  T_895;
  wire [5:0] req_idx;
  wire  fire;
  wire [19:0] T_898;
  wire [2:0] T_899;
  wire [8:0] T_900;
  wire [11:0] GEN_32;
  wire [11:0] T_901;
  reg [3:0] GEN_1;
  reg [31:0] GEN_41;
  assign io_req_ready = T_895;
  assign io_meta_read_valid = fire;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_1;
  assign io_meta_read_bits_tag = T_898;
  assign io_data_req_valid = fire;
  assign io_data_req_bits_way_en = req_way_en;
  assign io_data_req_bits_addr = T_901;
  assign io_release_valid = GEN_18;
  assign io_release_bits_addr_beat = beat_cnt;
  assign io_release_bits_addr_block = req_addr_block;
  assign io_release_bits_client_xact_id = req_client_xact_id;
  assign io_release_bits_voluntary = req_voluntary;
  assign io_release_bits_r_type = req_r_type;
  assign io_release_bits_data = io_data_resp;
  assign T_748 = io_release_ready & io_release_valid;
  assign GEN_29 = {{2'd0}, 1'h1};
  assign T_753 = beat_cnt + GEN_29;
  assign T_754 = T_753[2:0];
  assign GEN_0 = T_748 ? T_754 : beat_cnt;
  assign T_864 = io_data_req_ready & io_data_req_valid;
  assign T_865 = io_meta_read_ready & io_meta_read_valid;
  assign T_866 = T_864 & T_865;
  assign GEN_30 = {{3'd0}, 1'h1};
  assign T_869 = data_req_cnt + GEN_30;
  assign T_870 = T_869[3:0];
  assign GEN_2 = T_866 ? T_870 : data_req_cnt;
  assign T_872 = io_release_ready == 1'h0;
  assign T_879 = r1_data_req_fired ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_31 = {{2'd0}, T_879};
  assign T_880 = data_req_cnt - GEN_31;
  assign T_881 = T_880[3:0];
  assign GEN_3 = T_872 ? 1'h0 : T_866;
  assign GEN_4 = T_872 ? 1'h0 : r1_data_req_fired;
  assign GEN_5 = T_872 ? T_881 : GEN_2;
  assign T_885 = r1_data_req_fired == 1'h0;
  assign T_887 = data_req_cnt < 4'h8;
  assign T_890 = T_887 | T_872;
  assign GEN_9 = T_885 ? T_890 : active;
  assign GEN_11 = r2_data_req_fired ? GEN_3 : T_866;
  assign GEN_12 = r2_data_req_fired ? GEN_4 : r1_data_req_fired;
  assign GEN_13 = r2_data_req_fired ? GEN_5 : GEN_2;
  assign GEN_14 = r2_data_req_fired ? GEN_9 : active;
  assign GEN_15 = active ? GEN_11 : r1_data_req_fired;
  assign GEN_16 = active ? GEN_12 : r2_data_req_fired;
  assign GEN_17 = active ? GEN_13 : data_req_cnt;
  assign GEN_18 = active ? r2_data_req_fired : 1'h0;
  assign GEN_19 = active ? GEN_14 : active;
  assign T_891 = io_req_ready & io_req_valid;
  assign GEN_20 = T_891 ? 1'h1 : GEN_19;
  assign GEN_21 = T_891 ? {{3'd0}, 1'h0} : GEN_17;
  assign GEN_22 = T_891 ? io_req_bits_addr_beat : req_addr_beat;
  assign GEN_23 = T_891 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_24 = T_891 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign GEN_25 = T_891 ? io_req_bits_voluntary : req_voluntary;
  assign GEN_26 = T_891 ? io_req_bits_r_type : req_r_type;
  assign GEN_27 = T_891 ? io_req_bits_data : req_data;
  assign GEN_28 = T_891 ? io_req_bits_way_en : req_way_en;
  assign T_895 = active == 1'h0;
  assign req_idx = req_addr_block[5:0];
  assign fire = active & T_887;
  assign T_898 = req_addr_block[25:6];
  assign T_899 = data_req_cnt[2:0];
  assign T_900 = {req_idx,T_899};
  assign GEN_32 = {{3'd0}, T_900};
  assign T_901 = GEN_32 << 3;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_6 = {1{$random}};
  active = GEN_6[0:0];
  GEN_7 = {1{$random}};
  r1_data_req_fired = GEN_7[0:0];
  GEN_8 = {1{$random}};
  r2_data_req_fired = GEN_8[0:0];
  GEN_10 = {1{$random}};
  data_req_cnt = GEN_10[3:0];
  GEN_33 = {1{$random}};
  beat_cnt = GEN_33[2:0];
  GEN_34 = {1{$random}};
  req_addr_beat = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_addr_block = GEN_35[25:0];
  GEN_36 = {1{$random}};
  req_client_xact_id = GEN_36[1:0];
  GEN_37 = {1{$random}};
  req_voluntary = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_r_type = GEN_38[2:0];
  GEN_39 = {2{$random}};
  req_data = GEN_39[63:0];
  GEN_40 = {1{$random}};
  req_way_en = GEN_40[3:0];
  GEN_41 = {1{$random}};
  GEN_1 = GEN_41[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      active <= 1'h0;
    end else begin
      active <= GEN_20;
    end
    if(reset) begin
      r1_data_req_fired <= 1'h0;
    end else begin
      r1_data_req_fired <= GEN_15;
    end
    if(reset) begin
      r2_data_req_fired <= 1'h0;
    end else begin
      r2_data_req_fired <= GEN_16;
    end
    if(reset) begin
      data_req_cnt <= 4'h0;
    end else begin
      data_req_cnt <= GEN_21;
    end
    if(reset) begin
      beat_cnt <= 3'h0;
    end else begin
      beat_cnt <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      req_addr_beat <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      req_addr_block <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      req_client_xact_id <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      req_voluntary <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      req_r_type <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      req_data <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      req_way_en <= GEN_28;
    end
  end
endmodule
module ProbeUnit(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [25:0] io_req_bits_addr_block,
  input  [1:0] io_req_bits_p_type,
  input  [1:0] io_req_bits_client_xact_id,
  input   io_rep_ready,
  output  io_rep_valid,
  output [2:0] io_rep_bits_addr_beat,
  output [25:0] io_rep_bits_addr_block,
  output [1:0] io_rep_bits_client_xact_id,
  output  io_rep_bits_voluntary,
  output [2:0] io_rep_bits_r_type,
  output [63:0] io_rep_bits_data,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  input  [3:0] io_way_en,
  input   io_mshr_rdy,
  input  [1:0] io_block_state_state
);
  reg [3:0] state;
  reg [31:0] GEN_17;
  reg [1:0] old_coh_state;
  reg [31:0] GEN_18;
  reg [3:0] way_en;
  reg [31:0] GEN_19;
  reg [25:0] req_addr_block;
  reg [31:0] GEN_20;
  reg [1:0] req_p_type;
  reg [31:0] GEN_21;
  reg [1:0] req_client_xact_id;
  reg [31:0] GEN_22;
  wire [3:0] GEN_16;
  wire  tag_matches;
  wire [1:0] miss_coh_state;
  wire [1:0] reply_coh_state;
  wire [1:0] T_1256_0;
  wire  T_1258;
  wire [2:0] T_1261;
  wire [1:0] T_1275_0;
  wire  T_1277;
  wire [2:0] T_1281;
  wire [1:0] T_1294_0;
  wire  T_1296;
  wire [2:0] T_1301;
  wire  T_1308;
  wire [2:0] T_1309;
  wire  T_1310;
  wire [2:0] T_1311;
  wire  T_1312;
  wire [2:0] T_1313;
  wire [2:0] reply_addr_beat;
  wire [25:0] reply_addr_block;
  wire [1:0] reply_client_xact_id;
  wire  reply_voluntary;
  wire [2:0] reply_r_type;
  wire [63:0] reply_data;
  wire  T_1374;
  wire  T_1375;
  wire  T_1377;
  wire [2:0] T_1383_0;
  wire [2:0] T_1383_1;
  wire [2:0] T_1383_2;
  wire  T_1385;
  wire  T_1386;
  wire  T_1387;
  wire  T_1390;
  wire  T_1391;
  wire  T_1393;
  wire  T_1394;
  wire  T_1395;
  wire  T_1397;
  wire  T_1398;
  wire [19:0] T_1399;
  wire  T_1400;
  wire [1:0] T_1405;
  wire [1:0] T_1407;
  wire [1:0] T_1433_state;
  wire  T_1458;
  wire  T_1459;
  wire [3:0] GEN_0;
  wire [25:0] GEN_1;
  wire [1:0] GEN_2;
  wire [1:0] GEN_3;
  wire  T_1460;
  wire [3:0] GEN_4;
  wire  T_1461;
  wire [3:0] GEN_5;
  wire  T_1462;
  wire  T_1464;
  wire [3:0] GEN_6;
  wire [3:0] GEN_7;
  wire [1:0] GEN_8;
  wire [3:0] GEN_9;
  wire  T_1465;
  wire [1:0] T_1471_0;
  wire  T_1473;
  wire  T_1476;
  wire [3:0] T_1477;
  wire [3:0] GEN_11;
  wire  T_1479;
  wire [3:0] T_1480;
  wire [3:0] GEN_12;
  wire  T_1481;
  wire [3:0] GEN_13;
  wire  T_1482;
  wire  T_1483;
  wire [3:0] GEN_14;
  wire  T_1484;
  wire [3:0] GEN_15;
  reg [3:0] GEN_10;
  reg [31:0] GEN_23;
  assign io_req_ready = T_1374;
  assign io_rep_valid = T_1375;
  assign io_rep_bits_addr_beat = reply_addr_beat;
  assign io_rep_bits_addr_block = reply_addr_block;
  assign io_rep_bits_client_xact_id = reply_client_xact_id;
  assign io_rep_bits_voluntary = reply_voluntary;
  assign io_rep_bits_r_type = reply_r_type;
  assign io_rep_bits_data = reply_data;
  assign io_meta_read_valid = T_1398;
  assign io_meta_read_bits_idx = req_addr_block[5:0];
  assign io_meta_read_bits_way_en = GEN_10;
  assign io_meta_read_bits_tag = T_1399;
  assign io_meta_write_valid = T_1400;
  assign io_meta_write_bits_idx = req_addr_block[5:0];
  assign io_meta_write_bits_way_en = way_en;
  assign io_meta_write_bits_data_tag = T_1399;
  assign io_meta_write_bits_data_coh_state = T_1433_state;
  assign io_wb_req_valid = T_1458;
  assign io_wb_req_bits_addr_beat = reply_addr_beat;
  assign io_wb_req_bits_addr_block = reply_addr_block;
  assign io_wb_req_bits_client_xact_id = reply_client_xact_id;
  assign io_wb_req_bits_voluntary = reply_voluntary;
  assign io_wb_req_bits_r_type = reply_r_type;
  assign io_wb_req_bits_data = reply_data;
  assign io_wb_req_bits_way_en = way_en;
  assign GEN_16 = {{3'd0}, 1'h0};
  assign tag_matches = way_en != GEN_16;
  assign miss_coh_state = {{1'd0}, 1'h0};
  assign reply_coh_state = tag_matches ? old_coh_state : miss_coh_state;
  assign T_1256_0 = 2'h3;
  assign T_1258 = T_1256_0 == reply_coh_state;
  assign T_1261 = T_1258 ? 3'h0 : 3'h3;
  assign T_1275_0 = 2'h3;
  assign T_1277 = T_1275_0 == reply_coh_state;
  assign T_1281 = T_1277 ? 3'h1 : 3'h4;
  assign T_1294_0 = 2'h3;
  assign T_1296 = T_1294_0 == reply_coh_state;
  assign T_1301 = T_1296 ? 3'h2 : 3'h5;
  assign T_1308 = 2'h2 == req_p_type;
  assign T_1309 = T_1308 ? T_1301 : 3'h3;
  assign T_1310 = 2'h1 == req_p_type;
  assign T_1311 = T_1310 ? T_1281 : T_1309;
  assign T_1312 = 2'h0 == req_p_type;
  assign T_1313 = T_1312 ? T_1261 : T_1311;
  assign reply_addr_beat = {{2'd0}, 1'h0};
  assign reply_addr_block = req_addr_block;
  assign reply_client_xact_id = {{1'd0}, 1'h0};
  assign reply_voluntary = 1'h0;
  assign reply_r_type = T_1313;
  assign reply_data = {{63'd0}, 1'h0};
  assign T_1374 = state == 4'h0;
  assign T_1375 = state == 4'h5;
  assign T_1377 = io_rep_valid == 1'h0;
  assign T_1383_0 = 3'h0;
  assign T_1383_1 = 3'h1;
  assign T_1383_2 = 3'h2;
  assign T_1385 = T_1383_0 == io_rep_bits_r_type;
  assign T_1386 = T_1383_1 == io_rep_bits_r_type;
  assign T_1387 = T_1383_2 == io_rep_bits_r_type;
  assign T_1390 = T_1385 | T_1386;
  assign T_1391 = T_1390 | T_1387;
  assign T_1393 = T_1391 == 1'h0;
  assign T_1394 = T_1377 | T_1393;
  assign T_1395 = T_1394 | reset;
  assign T_1397 = T_1395 == 1'h0;
  assign T_1398 = state == 4'h1;
  assign T_1399 = req_addr_block[25:6];
  assign T_1400 = state == 4'h8;
  assign T_1405 = T_1310 ? 2'h1 : old_coh_state;
  assign T_1407 = T_1312 ? 2'h0 : T_1405;
  assign T_1433_state = T_1407;
  assign T_1458 = state == 4'h6;
  assign T_1459 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1459 ? 4'h1 : state;
  assign GEN_1 = T_1459 ? io_req_bits_addr_block : req_addr_block;
  assign GEN_2 = T_1459 ? io_req_bits_p_type : req_p_type;
  assign GEN_3 = T_1459 ? io_req_bits_client_xact_id : req_client_xact_id;
  assign T_1460 = io_meta_read_ready & io_meta_read_valid;
  assign GEN_4 = T_1460 ? 4'h2 : GEN_0;
  assign T_1461 = state == 4'h2;
  assign GEN_5 = T_1461 ? 4'h3 : GEN_4;
  assign T_1462 = state == 4'h3;
  assign T_1464 = io_mshr_rdy == 1'h0;
  assign GEN_6 = T_1464 ? 4'h1 : 4'h4;
  assign GEN_7 = T_1462 ? GEN_6 : GEN_5;
  assign GEN_8 = T_1462 ? io_block_state_state : old_coh_state;
  assign GEN_9 = T_1462 ? io_way_en : way_en;
  assign T_1465 = state == 4'h4;
  assign T_1471_0 = 2'h3;
  assign T_1473 = T_1471_0 == old_coh_state;
  assign T_1476 = tag_matches & T_1473;
  assign T_1477 = T_1476 ? 4'h6 : 4'h5;
  assign GEN_11 = T_1465 ? T_1477 : GEN_7;
  assign T_1479 = T_1375 & io_rep_ready;
  assign T_1480 = tag_matches ? 4'h8 : 4'h0;
  assign GEN_12 = T_1479 ? T_1480 : GEN_11;
  assign T_1481 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_13 = T_1481 ? 4'h7 : GEN_12;
  assign T_1482 = state == 4'h7;
  assign T_1483 = T_1482 & io_wb_req_ready;
  assign GEN_14 = T_1483 ? 4'h8 : GEN_13;
  assign T_1484 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_15 = T_1484 ? 4'h0 : GEN_14;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_17 = {1{$random}};
  state = GEN_17[3:0];
  GEN_18 = {1{$random}};
  old_coh_state = GEN_18[1:0];
  GEN_19 = {1{$random}};
  way_en = GEN_19[3:0];
  GEN_20 = {1{$random}};
  req_addr_block = GEN_20[25:0];
  GEN_21 = {1{$random}};
  req_p_type = GEN_21[1:0];
  GEN_22 = {1{$random}};
  req_client_xact_id = GEN_22[1:0];
  GEN_23 = {1{$random}};
  GEN_10 = GEN_23[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      state <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      old_coh_state <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      way_en <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      req_addr_block <= GEN_1;
    end
    if(1'h0) begin
    end else begin
      req_p_type <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      req_client_xact_id <= GEN_3;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1397) begin
          $fwrite(32'h80000002,"Assertion failed: ProbeUnit should not send releases with data\n    at nbdcache.scala:669 assert(!io.rep.valid || !io.rep.bits.hasData(),\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1397) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module Arbiter_67(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_tag,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_tag,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_tag,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire  T_630;
  wire  T_632;
  wire  T_634;
  wire  T_635;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_632;
  assign io_out_valid = T_635;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_tag = GEN_3;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign T_630 = io_in_0_valid == 1'h0;
  assign T_632 = T_630 & io_out_ready;
  assign T_634 = T_630 == 1'h0;
  assign T_635 = T_634 | io_in_1_valid;
endmodule
module Arbiter_68(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  input  [19:0] io_in_0_bits_data_tag,
  input  [1:0] io_in_0_bits_data_coh_state,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  input  [19:0] io_in_1_bits_data_tag,
  input  [1:0] io_in_1_bits_data_coh_state,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [19:0] io_out_bits_data_tag,
  output [1:0] io_out_bits_data_coh_state,
  output  io_chosen
);
  wire  GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [19:0] GEN_3;
  wire [1:0] GEN_4;
  wire  T_2720;
  wire  T_2722;
  wire  T_2724;
  wire  T_2725;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2722;
  assign io_out_valid = T_2725;
  assign io_out_bits_idx = GEN_1;
  assign io_out_bits_way_en = GEN_2;
  assign io_out_bits_data_tag = GEN_3;
  assign io_out_bits_data_coh_state = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_idx : io_in_1_bits_idx;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data_coh_state : io_in_1_bits_data_coh_state;
  assign T_2720 = io_in_0_valid == 1'h0;
  assign T_2722 = T_2720 & io_out_ready;
  assign T_2724 = T_2720 == 1'h0;
  assign T_2725 = T_2724 | io_in_1_valid;
endmodule
module LockingArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input  [2:0] io_in_0_bits_addr_beat,
  input   io_in_0_bits_is_builtin_type,
  input  [2:0] io_in_0_bits_a_type,
  input  [11:0] io_in_0_bits_union,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input  [2:0] io_in_1_bits_addr_beat,
  input   io_in_1_bits_is_builtin_type,
  input  [2:0] io_in_1_bits_a_type,
  input  [11:0] io_in_1_bits_union,
  input  [63:0] io_in_1_bits_data,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [25:0] io_in_2_bits_addr_block,
  input  [1:0] io_in_2_bits_client_xact_id,
  input  [2:0] io_in_2_bits_addr_beat,
  input   io_in_2_bits_is_builtin_type,
  input  [2:0] io_in_2_bits_a_type,
  input  [11:0] io_in_2_bits_union,
  input  [63:0] io_in_2_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_addr_beat,
  output  io_out_bits_is_builtin_type,
  output [2:0] io_out_bits_a_type,
  output [11:0] io_out_bits_union,
  output [63:0] io_out_bits_data,
  output [1:0] io_chosen
);
  wire [1:0] choice;
  wire  GEN_0;
  wire [1:0] GEN_29;
  wire  GEN_8;
  wire  GEN_9;
  wire [25:0] GEN_1;
  wire [25:0] GEN_10;
  wire [25:0] GEN_11;
  wire [1:0] GEN_2;
  wire [1:0] GEN_12;
  wire [1:0] GEN_13;
  wire [2:0] GEN_3;
  wire [2:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_4;
  wire  GEN_16;
  wire  GEN_17;
  wire [2:0] GEN_5;
  wire [2:0] GEN_18;
  wire [2:0] GEN_19;
  wire [11:0] GEN_6;
  wire [11:0] GEN_20;
  wire [11:0] GEN_21;
  wire [63:0] GEN_7;
  wire [63:0] GEN_22;
  wire [63:0] GEN_23;
  reg [2:0] T_972;
  reg [31:0] GEN_30;
  reg [1:0] T_974;
  reg [31:0] GEN_31;
  wire [2:0] GEN_37;
  wire  T_976;
  wire [2:0] T_985_0;
  wire  T_987;
  wire  T_990;
  wire  T_991;
  wire  T_992;
  wire [2:0] GEN_38;
  wire [3:0] T_996;
  wire [2:0] T_997;
  wire [1:0] GEN_24;
  wire [2:0] GEN_25;
  wire [1:0] GEN_26;
  wire  T_999;
  wire  T_1001;
  wire  T_1003;
  wire [1:0] GEN_39;
  wire  T_1005;
  wire  T_1006;
  wire  T_1007;
  wire  T_1009;
  wire  T_1010;
  wire  T_1011;
  wire  T_1013;
  wire  T_1014;
  wire  T_1015;
  wire [1:0] GEN_27;
  wire [1:0] GEN_28;
  assign io_in_0_ready = T_1007;
  assign io_in_1_ready = T_1011;
  assign io_in_2_ready = T_1015;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_block = GEN_1;
  assign io_out_bits_client_xact_id = GEN_2;
  assign io_out_bits_addr_beat = GEN_3;
  assign io_out_bits_is_builtin_type = GEN_4;
  assign io_out_bits_a_type = GEN_5;
  assign io_out_bits_union = GEN_6;
  assign io_out_bits_data = GEN_7;
  assign io_chosen = GEN_26;
  assign choice = GEN_28;
  assign GEN_0 = GEN_9;
  assign GEN_29 = {{1'd0}, 1'h1};
  assign GEN_8 = GEN_29 == io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_9 = 2'h2 == io_chosen ? io_in_2_valid : GEN_8;
  assign GEN_1 = GEN_11;
  assign GEN_10 = GEN_29 == io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_11 = 2'h2 == io_chosen ? io_in_2_bits_addr_block : GEN_10;
  assign GEN_2 = GEN_13;
  assign GEN_12 = GEN_29 == io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_13 = 2'h2 == io_chosen ? io_in_2_bits_client_xact_id : GEN_12;
  assign GEN_3 = GEN_15;
  assign GEN_14 = GEN_29 == io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_15 = 2'h2 == io_chosen ? io_in_2_bits_addr_beat : GEN_14;
  assign GEN_4 = GEN_17;
  assign GEN_16 = GEN_29 == io_chosen ? io_in_1_bits_is_builtin_type : io_in_0_bits_is_builtin_type;
  assign GEN_17 = 2'h2 == io_chosen ? io_in_2_bits_is_builtin_type : GEN_16;
  assign GEN_5 = GEN_19;
  assign GEN_18 = GEN_29 == io_chosen ? io_in_1_bits_a_type : io_in_0_bits_a_type;
  assign GEN_19 = 2'h2 == io_chosen ? io_in_2_bits_a_type : GEN_18;
  assign GEN_6 = GEN_21;
  assign GEN_20 = GEN_29 == io_chosen ? io_in_1_bits_union : io_in_0_bits_union;
  assign GEN_21 = 2'h2 == io_chosen ? io_in_2_bits_union : GEN_20;
  assign GEN_7 = GEN_23;
  assign GEN_22 = GEN_29 == io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_23 = 2'h2 == io_chosen ? io_in_2_bits_data : GEN_22;
  assign GEN_37 = {{2'd0}, 1'h0};
  assign T_976 = T_972 != GEN_37;
  assign T_985_0 = 3'h3;
  assign T_987 = T_985_0 == io_out_bits_a_type;
  assign T_990 = io_out_bits_is_builtin_type & T_987;
  assign T_991 = io_out_ready & io_out_valid;
  assign T_992 = T_991 & T_990;
  assign GEN_38 = {{2'd0}, 1'h1};
  assign T_996 = T_972 + GEN_38;
  assign T_997 = T_996[2:0];
  assign GEN_24 = T_992 ? io_chosen : T_974;
  assign GEN_25 = T_992 ? T_997 : T_972;
  assign GEN_26 = T_976 ? T_974 : choice;
  assign T_999 = io_in_0_valid | io_in_1_valid;
  assign T_1001 = io_in_0_valid == 1'h0;
  assign T_1003 = T_999 == 1'h0;
  assign GEN_39 = {{1'd0}, 1'h0};
  assign T_1005 = T_974 == GEN_39;
  assign T_1006 = T_976 ? T_1005 : 1'h1;
  assign T_1007 = T_1006 & io_out_ready;
  assign T_1009 = T_974 == GEN_29;
  assign T_1010 = T_976 ? T_1009 : T_1001;
  assign T_1011 = T_1010 & io_out_ready;
  assign T_1013 = T_974 == 2'h2;
  assign T_1014 = T_976 ? T_1013 : T_1003;
  assign T_1015 = T_1014 & io_out_ready;
  assign GEN_27 = io_in_1_valid ? {{1'd0}, 1'h1} : 2'h2;
  assign GEN_28 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_27;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  T_972 = GEN_30[2:0];
  GEN_31 = {1{$random}};
  T_974 = GEN_31[1:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_972 <= 3'h0;
    end else begin
      T_972 <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      T_974 <= GEN_24;
    end
  end
endmodule
module Arbiter_69(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_manager_xact_id,
  input   io_in_0_bits_manager_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_manager_xact_id,
  input   io_in_1_bits_manager_id,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [2:0] io_in_2_bits_manager_xact_id,
  input   io_in_2_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_manager_id,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [2:0] GEN_1;
  wire  GEN_2;
  wire [1:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire  T_716;
  wire  T_718;
  wire  T_720;
  wire  T_722;
  wire  T_723;
  wire  T_725;
  wire  T_726;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_722;
  assign io_in_2_ready = T_723;
  assign io_out_valid = T_726;
  assign io_out_bits_manager_xact_id = GEN_4;
  assign io_out_bits_manager_id = GEN_5;
  assign io_chosen = GEN_3;
  assign GEN_0 = io_in_1_valid ? {{1'd0}, 1'h1} : 2'h2;
  assign GEN_1 = io_in_1_valid ? io_in_1_bits_manager_xact_id : io_in_2_bits_manager_xact_id;
  assign GEN_2 = io_in_1_valid ? io_in_1_bits_manager_id : io_in_2_bits_manager_id;
  assign GEN_3 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_0;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_manager_xact_id : GEN_1;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_manager_id : GEN_2;
  assign T_716 = io_in_0_valid | io_in_1_valid;
  assign T_718 = io_in_0_valid == 1'h0;
  assign T_720 = T_716 == 1'h0;
  assign T_722 = T_718 & io_out_ready;
  assign T_723 = T_720 & io_out_ready;
  assign T_725 = T_720 == 1'h0;
  assign T_726 = T_725 | io_in_2_valid;
endmodule
module Arbiter_70(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input  [3:0] io_in_1_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output [3:0] io_out_bits_way_en,
  output  io_chosen
);
  wire  GEN_0;
  wire [2:0] GEN_1;
  wire [25:0] GEN_2;
  wire [1:0] GEN_3;
  wire  GEN_4;
  wire [2:0] GEN_5;
  wire [63:0] GEN_6;
  wire [3:0] GEN_7;
  wire  T_1224;
  wire  T_1226;
  wire  T_1228;
  wire  T_1229;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1226;
  assign io_out_valid = T_1229;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_out_bits_way_en = GEN_7;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr_beat : io_in_1_bits_addr_beat;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr_block : io_in_1_bits_addr_block;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_client_xact_id : io_in_1_bits_client_xact_id;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_voluntary : io_in_1_bits_voluntary;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_r_type : io_in_1_bits_r_type;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign T_1224 = io_in_0_valid == 1'h0;
  assign T_1226 = T_1224 & io_out_ready;
  assign T_1228 = T_1224 == 1'h0;
  assign T_1229 = T_1228 | io_in_1_valid;
endmodule
module Arbiter_71(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [8:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input   io_in_0_bits_phys,
  input  [4:0] io_in_0_bits_sdq_id,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [39:0] io_in_1_bits_addr,
  input  [8:0] io_in_1_bits_tag,
  input  [4:0] io_in_1_bits_cmd,
  input  [2:0] io_in_1_bits_typ,
  input   io_in_1_bits_phys,
  input  [4:0] io_in_1_bits_sdq_id,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [8:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output  io_out_bits_phys,
  output [4:0] io_out_bits_sdq_id,
  output  io_chosen
);
  wire  GEN_0;
  wire [39:0] GEN_1;
  wire [8:0] GEN_2;
  wire [4:0] GEN_3;
  wire [2:0] GEN_4;
  wire  GEN_5;
  wire [4:0] GEN_6;
  wire  T_1708;
  wire  T_1710;
  wire  T_1712;
  wire  T_1713;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1710;
  assign io_out_valid = T_1713;
  assign io_out_bits_addr = GEN_1;
  assign io_out_bits_tag = GEN_2;
  assign io_out_bits_cmd = GEN_3;
  assign io_out_bits_typ = GEN_4;
  assign io_out_bits_phys = GEN_5;
  assign io_out_bits_sdq_id = GEN_6;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_typ : io_in_1_bits_typ;
  assign GEN_5 = io_in_0_valid ? io_in_0_bits_phys : io_in_1_bits_phys;
  assign GEN_6 = io_in_0_valid ? io_in_0_bits_sdq_id : io_in_1_bits_sdq_id;
  assign T_1708 = io_in_0_valid == 1'h0;
  assign T_1710 = T_1708 & io_out_ready;
  assign T_1712 = T_1708 == 1'h0;
  assign T_1713 = T_1712 | io_in_1_valid;
endmodule
module Arbiter_72(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_in_1_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  wire  GEN_0;
  wire  GEN_1;
  wire  T_58;
  wire  T_60;
  wire  T_62;
  wire  T_63;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_60;
  assign io_out_valid = T_63;
  assign io_out_bits = GEN_1;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits : io_in_1_bits;
  assign T_58 = io_in_0_valid == 1'h0;
  assign T_60 = T_58 & io_out_ready;
  assign T_62 = T_58 == 1'h0;
  assign T_63 = T_62 | io_in_1_valid;
endmodule
module Queue_73(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [39:0] io_enq_bits_addr,
  input  [8:0] io_enq_bits_tag,
  input  [4:0] io_enq_bits_cmd,
  input  [2:0] io_enq_bits_typ,
  input   io_enq_bits_phys,
  input  [4:0] io_enq_bits_sdq_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [39:0] io_deq_bits_addr,
  output [8:0] io_deq_bits_tag,
  output [4:0] io_deq_bits_cmd,
  output [2:0] io_deq_bits_typ,
  output  io_deq_bits_phys,
  output [4:0] io_deq_bits_sdq_id,
  output [4:0] io_count
);
  reg [39:0] ram_addr [0:15];
  reg [63:0] GEN_0;
  wire [39:0] ram_addr_T_794_data;
  wire [3:0] ram_addr_T_794_addr;
  wire  ram_addr_T_794_en;
  wire [39:0] ram_addr_T_703_data;
  wire [3:0] ram_addr_T_703_addr;
  wire  ram_addr_T_703_mask;
  wire  ram_addr_T_703_en;
  reg [8:0] ram_tag [0:15];
  reg [31:0] GEN_1;
  wire [8:0] ram_tag_T_794_data;
  wire [3:0] ram_tag_T_794_addr;
  wire  ram_tag_T_794_en;
  wire [8:0] ram_tag_T_703_data;
  wire [3:0] ram_tag_T_703_addr;
  wire  ram_tag_T_703_mask;
  wire  ram_tag_T_703_en;
  reg [4:0] ram_cmd [0:15];
  reg [31:0] GEN_2;
  wire [4:0] ram_cmd_T_794_data;
  wire [3:0] ram_cmd_T_794_addr;
  wire  ram_cmd_T_794_en;
  wire [4:0] ram_cmd_T_703_data;
  wire [3:0] ram_cmd_T_703_addr;
  wire  ram_cmd_T_703_mask;
  wire  ram_cmd_T_703_en;
  reg [2:0] ram_typ [0:15];
  reg [31:0] GEN_3;
  wire [2:0] ram_typ_T_794_data;
  wire [3:0] ram_typ_T_794_addr;
  wire  ram_typ_T_794_en;
  wire [2:0] ram_typ_T_703_data;
  wire [3:0] ram_typ_T_703_addr;
  wire  ram_typ_T_703_mask;
  wire  ram_typ_T_703_en;
  reg  ram_phys [0:15];
  reg [31:0] GEN_4;
  wire  ram_phys_T_794_data;
  wire [3:0] ram_phys_T_794_addr;
  wire  ram_phys_T_794_en;
  wire  ram_phys_T_703_data;
  wire [3:0] ram_phys_T_703_addr;
  wire  ram_phys_T_703_mask;
  wire  ram_phys_T_703_en;
  reg [4:0] ram_sdq_id [0:15];
  reg [31:0] GEN_5;
  wire [4:0] ram_sdq_id_T_794_data;
  wire [3:0] ram_sdq_id_T_794_addr;
  wire  ram_sdq_id_T_794_en;
  wire [4:0] ram_sdq_id_T_703_data;
  wire [3:0] ram_sdq_id_T_703_addr;
  wire  ram_sdq_id_T_703_mask;
  wire  ram_sdq_id_T_703_en;
  reg [3:0] T_695;
  reg [31:0] GEN_6;
  reg [3:0] T_697;
  reg [31:0] GEN_7;
  reg  maybe_full;
  reg [31:0] GEN_8;
  wire  ptr_match;
  wire  T_700;
  wire  empty;
  wire  full;
  wire  T_701;
  wire  do_enq;
  wire  T_702;
  wire  do_deq;
  wire [3:0] GEN_18;
  wire [4:0] T_782;
  wire [3:0] T_783;
  wire [3:0] GEN_15;
  wire [4:0] T_787;
  wire [3:0] T_788;
  wire [3:0] GEN_16;
  wire  T_789;
  wire  GEN_17;
  wire  T_791;
  wire  T_793;
  wire [4:0] T_870;
  wire [3:0] ptr_diff;
  wire  T_871;
  wire [4:0] T_872;
  assign io_enq_ready = T_793;
  assign io_deq_valid = T_791;
  assign io_deq_bits_addr = ram_addr_T_794_data;
  assign io_deq_bits_tag = ram_tag_T_794_data;
  assign io_deq_bits_cmd = ram_cmd_T_794_data;
  assign io_deq_bits_typ = ram_typ_T_794_data;
  assign io_deq_bits_phys = ram_phys_T_794_data;
  assign io_deq_bits_sdq_id = ram_sdq_id_T_794_data;
  assign io_count = T_872;
  assign ram_addr_T_794_addr = T_697;
  assign ram_addr_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_addr_T_794_data = ram_addr[ram_addr_T_794_addr];
  `else
  assign ram_addr_T_794_data = ram_addr_T_794_addr >= 5'h10 ? $random : ram_addr[ram_addr_T_794_addr];
  `endif
  assign ram_addr_T_703_data = io_enq_bits_addr;
  assign ram_addr_T_703_addr = T_695;
  assign ram_addr_T_703_mask = do_enq;
  assign ram_addr_T_703_en = do_enq;
  assign ram_tag_T_794_addr = T_697;
  assign ram_tag_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_tag_T_794_data = ram_tag[ram_tag_T_794_addr];
  `else
  assign ram_tag_T_794_data = ram_tag_T_794_addr >= 5'h10 ? $random : ram_tag[ram_tag_T_794_addr];
  `endif
  assign ram_tag_T_703_data = io_enq_bits_tag;
  assign ram_tag_T_703_addr = T_695;
  assign ram_tag_T_703_mask = do_enq;
  assign ram_tag_T_703_en = do_enq;
  assign ram_cmd_T_794_addr = T_697;
  assign ram_cmd_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_cmd_T_794_data = ram_cmd[ram_cmd_T_794_addr];
  `else
  assign ram_cmd_T_794_data = ram_cmd_T_794_addr >= 5'h10 ? $random : ram_cmd[ram_cmd_T_794_addr];
  `endif
  assign ram_cmd_T_703_data = io_enq_bits_cmd;
  assign ram_cmd_T_703_addr = T_695;
  assign ram_cmd_T_703_mask = do_enq;
  assign ram_cmd_T_703_en = do_enq;
  assign ram_typ_T_794_addr = T_697;
  assign ram_typ_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_typ_T_794_data = ram_typ[ram_typ_T_794_addr];
  `else
  assign ram_typ_T_794_data = ram_typ_T_794_addr >= 5'h10 ? $random : ram_typ[ram_typ_T_794_addr];
  `endif
  assign ram_typ_T_703_data = io_enq_bits_typ;
  assign ram_typ_T_703_addr = T_695;
  assign ram_typ_T_703_mask = do_enq;
  assign ram_typ_T_703_en = do_enq;
  assign ram_phys_T_794_addr = T_697;
  assign ram_phys_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_phys_T_794_data = ram_phys[ram_phys_T_794_addr];
  `else
  assign ram_phys_T_794_data = ram_phys_T_794_addr >= 5'h10 ? $random : ram_phys[ram_phys_T_794_addr];
  `endif
  assign ram_phys_T_703_data = io_enq_bits_phys;
  assign ram_phys_T_703_addr = T_695;
  assign ram_phys_T_703_mask = do_enq;
  assign ram_phys_T_703_en = do_enq;
  assign ram_sdq_id_T_794_addr = T_697;
  assign ram_sdq_id_T_794_en = 1'h1;
  `ifdef SYNTHESIS
  assign ram_sdq_id_T_794_data = ram_sdq_id[ram_sdq_id_T_794_addr];
  `else
  assign ram_sdq_id_T_794_data = ram_sdq_id_T_794_addr >= 5'h10 ? $random : ram_sdq_id[ram_sdq_id_T_794_addr];
  `endif
  assign ram_sdq_id_T_703_data = io_enq_bits_sdq_id;
  assign ram_sdq_id_T_703_addr = T_695;
  assign ram_sdq_id_T_703_mask = do_enq;
  assign ram_sdq_id_T_703_en = do_enq;
  assign ptr_match = T_695 == T_697;
  assign T_700 = maybe_full == 1'h0;
  assign empty = ptr_match & T_700;
  assign full = ptr_match & maybe_full;
  assign T_701 = io_enq_ready & io_enq_valid;
  assign do_enq = T_701;
  assign T_702 = io_deq_ready & io_deq_valid;
  assign do_deq = T_702;
  assign GEN_18 = {{3'd0}, 1'h1};
  assign T_782 = T_695 + GEN_18;
  assign T_783 = T_782[3:0];
  assign GEN_15 = do_enq ? T_783 : T_695;
  assign T_787 = T_697 + GEN_18;
  assign T_788 = T_787[3:0];
  assign GEN_16 = do_deq ? T_788 : T_697;
  assign T_789 = do_enq != do_deq;
  assign GEN_17 = T_789 ? do_enq : maybe_full;
  assign T_791 = empty == 1'h0;
  assign T_793 = full == 1'h0;
  assign T_870 = T_695 - T_697;
  assign ptr_diff = T_870[3:0];
  assign T_871 = maybe_full & ptr_match;
  assign T_872 = {T_871,ptr_diff};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {2{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_addr[initvar] = GEN_0[39:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_tag[initvar] = GEN_1[8:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_cmd[initvar] = GEN_2[4:0];
  GEN_3 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_typ[initvar] = GEN_3[2:0];
  GEN_4 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_phys[initvar] = GEN_4[0:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram_sdq_id[initvar] = GEN_5[4:0];
  GEN_6 = {1{$random}};
  T_695 = GEN_6[3:0];
  GEN_7 = {1{$random}};
  T_697 = GEN_7[3:0];
  GEN_8 = {1{$random}};
  maybe_full = GEN_8[0:0];
  end
`endif
  always @(posedge clk) begin
    if(ram_addr_T_703_en & ram_addr_T_703_mask) begin
      ram_addr[ram_addr_T_703_addr] <= ram_addr_T_703_data;
    end
    if(ram_tag_T_703_en & ram_tag_T_703_mask) begin
      ram_tag[ram_tag_T_703_addr] <= ram_tag_T_703_data;
    end
    if(ram_cmd_T_703_en & ram_cmd_T_703_mask) begin
      ram_cmd[ram_cmd_T_703_addr] <= ram_cmd_T_703_data;
    end
    if(ram_typ_T_703_en & ram_typ_T_703_mask) begin
      ram_typ[ram_typ_T_703_addr] <= ram_typ_T_703_data;
    end
    if(ram_phys_T_703_en & ram_phys_T_703_mask) begin
      ram_phys[ram_phys_T_703_addr] <= ram_phys_T_703_data;
    end
    if(ram_sdq_id_T_703_en & ram_sdq_id_T_703_mask) begin
      ram_sdq_id[ram_sdq_id_T_703_addr] <= ram_sdq_id_T_703_data;
    end
    if(reset) begin
      T_695 <= 4'h0;
    end else begin
      T_695 <= GEN_15;
    end
    if(reset) begin
      T_697 <= 4'h0;
    end else begin
      T_697 <= GEN_16;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else begin
      maybe_full <= GEN_17;
    end
  end
endmodule
module FinishQueue_74(
  input   clk,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input  [2:0] io_enq_bits_manager_xact_id,
  input   io_enq_bits_manager_id,
  input   io_deq_ready,
  output  io_deq_valid,
  output [2:0] io_deq_bits_manager_xact_id,
  output  io_deq_bits_manager_id,
  output  io_count
);
  reg [2:0] T_244_manager_xact_id [0:0];
  reg [31:0] GEN_0;
  wire [2:0] T_244_manager_xact_id_T_291_data;
  wire  T_244_manager_xact_id_T_291_addr;
  wire  T_244_manager_xact_id_T_291_en;
  wire [2:0] T_244_manager_xact_id_T_258_data;
  wire  T_244_manager_xact_id_T_258_addr;
  wire  T_244_manager_xact_id_T_258_mask;
  wire  T_244_manager_xact_id_T_258_en;
  reg  T_244_manager_id [0:0];
  reg [31:0] GEN_1;
  wire  T_244_manager_id_T_291_data;
  wire  T_244_manager_id_T_291_addr;
  wire  T_244_manager_id_T_291_en;
  wire  T_244_manager_id_T_258_data;
  wire  T_244_manager_id_T_258_addr;
  wire  T_244_manager_id_T_258_mask;
  wire  T_244_manager_id_T_258_en;
  reg  T_248;
  reg [31:0] GEN_2;
  wire  T_251;
  wire  T_254;
  wire  T_255;
  wire  T_256;
  wire  T_257;
  wire  T_286;
  wire  GEN_7;
  wire  T_288;
  wire [1:0] T_317;
  wire  T_318;
  wire [1:0] T_320;
  assign io_enq_ready = T_251;
  assign io_deq_valid = T_288;
  assign io_deq_bits_manager_xact_id = T_244_manager_xact_id_T_291_data;
  assign io_deq_bits_manager_id = T_244_manager_id_T_291_data;
  assign io_count = T_320[0];
  assign T_244_manager_xact_id_T_291_addr = 1'h0;
  assign T_244_manager_xact_id_T_291_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_xact_id_T_291_data = T_244_manager_xact_id[T_244_manager_xact_id_T_291_addr];
  `else
  assign T_244_manager_xact_id_T_291_data = T_244_manager_xact_id_T_291_addr >= 1'h1 ? $random : T_244_manager_xact_id[T_244_manager_xact_id_T_291_addr];
  `endif
  assign T_244_manager_xact_id_T_258_data = io_enq_bits_manager_xact_id;
  assign T_244_manager_xact_id_T_258_addr = 1'h0;
  assign T_244_manager_xact_id_T_258_mask = T_255;
  assign T_244_manager_xact_id_T_258_en = T_255;
  assign T_244_manager_id_T_291_addr = 1'h0;
  assign T_244_manager_id_T_291_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_244_manager_id_T_291_data = T_244_manager_id[T_244_manager_id_T_291_addr];
  `else
  assign T_244_manager_id_T_291_data = T_244_manager_id_T_291_addr >= 1'h1 ? $random : T_244_manager_id[T_244_manager_id_T_291_addr];
  `endif
  assign T_244_manager_id_T_258_data = io_enq_bits_manager_id;
  assign T_244_manager_id_T_258_addr = 1'h0;
  assign T_244_manager_id_T_258_mask = T_255;
  assign T_244_manager_id_T_258_en = T_255;
  assign T_251 = T_248 == 1'h0;
  assign T_254 = io_enq_ready & io_enq_valid;
  assign T_255 = T_254;
  assign T_256 = io_deq_ready & io_deq_valid;
  assign T_257 = T_256;
  assign T_286 = T_255 != T_257;
  assign GEN_7 = T_286 ? T_255 : T_248;
  assign T_288 = T_251 == 1'h0;
  assign T_317 = 1'h0 - 1'h0;
  assign T_318 = T_317[0:0];
  assign T_320 = {T_248,T_318};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_0 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    T_244_manager_xact_id[initvar] = GEN_0[2:0];
  GEN_1 = {1{$random}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    T_244_manager_id[initvar] = GEN_1[0:0];
  GEN_2 = {1{$random}};
  T_248 = GEN_2[0:0];
  end
`endif
  always @(posedge clk) begin
    if(T_244_manager_xact_id_T_258_en & T_244_manager_xact_id_T_258_mask) begin
      T_244_manager_xact_id[T_244_manager_xact_id_T_258_addr] <= T_244_manager_xact_id_T_258_data;
    end
    if(T_244_manager_id_T_258_en & T_244_manager_id_T_258_mask) begin
      T_244_manager_id[T_244_manager_id_T_258_addr] <= T_244_manager_id_T_258_data;
    end
    if(reset) begin
      T_248 <= 1'h0;
    end else begin
      T_248 <= GEN_7;
    end
  end
endmodule
module MSHR(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_16;
  wire [1:0] T_1875_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_17;
  reg [39:0] req_addr;
  reg [63:0] GEN_18;
  reg [8:0] req_tag;
  reg [31:0] GEN_19;
  reg [4:0] req_cmd;
  reg [31:0] GEN_22;
  reg [2:0] req_typ;
  reg [31:0] GEN_34;
  reg  req_phys;
  reg [31:0] GEN_35;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_36;
  reg  req_tag_match;
  reg [31:0] GEN_37;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_38;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_41;
  reg [3:0] req_way_en;
  reg [31:0] GEN_57;
  wire [5:0] req_idx;
  wire [5:0] T_2271;
  wire  idx_match;
  wire  T_2272;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2278;
  wire  T_2279;
  wire  T_2280;
  wire  T_2281;
  wire  T_2282;
  wire  T_2283;
  wire  T_2284;
  wire  T_2285;
  wire  T_2286;
  wire  T_2287;
  wire  T_2288;
  wire  T_2289;
  wire  T_2290;
  wire  T_2291;
  wire  T_2292;
  wire  T_2293;
  wire  T_2295;
  wire  cmd_requires_second_acquire;
  wire [3:0] states_before_refill_0;
  wire [3:0] states_before_refill_1;
  wire [3:0] states_before_refill_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire [3:0] T_2314_0;
  wire [3:0] T_2314_1;
  wire  T_2316;
  wire  T_2317;
  wire  T_2320;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  sec_rdy;
  wire [2:0] T_2332_0;
  wire [3:0] GEN_46;
  wire  T_2334;
  wire [1:0] T_2342_0;
  wire [1:0] T_2342_1;
  wire [3:0] GEN_47;
  wire  T_2344;
  wire [3:0] GEN_48;
  wire  T_2345;
  wire  T_2348;
  wire  T_2349;
  wire  T_2350;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_58;
  wire  T_2353;
  wire [2:0] GEN_49;
  wire [3:0] T_2355;
  wire [2:0] T_2356;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2358;
  wire  T_2359;
  wire  refill_done;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [8:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [8:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire  T_2439;
  wire  T_2441;
  wire  T_2443;
  wire  T_2444;
  wire  T_2445;
  wire  T_2446;
  wire  T_2447;
  wire  T_2448;
  wire [1:0] T_2456;
  wire [3:0] GEN_50;
  wire  T_2457;
  wire [1:0] T_2458;
  wire [3:0] GEN_51;
  wire  T_2459;
  wire [1:0] T_2460;
  wire [3:0] GEN_52;
  wire  T_2461;
  wire [1:0] T_2462;
  wire [1:0] T_2463;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2520;
  wire [1:0] coh_on_hit_state;
  wire  T_2572;
  wire  T_2573;
  wire [3:0] GEN_1;
  wire  T_2574;
  wire [3:0] GEN_2;
  wire  T_2575;
  wire  T_2576;
  wire [3:0] GEN_3;
  wire  T_2577;
  wire  T_2578;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2579;
  wire [3:0] GEN_6;
  wire  T_2580;
  wire  T_2581;
  wire [3:0] GEN_7;
  wire  T_2582;
  wire  T_2583;
  wire [3:0] GEN_8;
  wire  T_2584;
  wire [3:0] GEN_9;
  wire  T_2589;
  wire [4:0] GEN_10;
  wire [4:0] GEN_11;
  wire [1:0] T_2607_0;
  wire [1:0] T_2607_1;
  wire  T_2609;
  wire  T_2610;
  wire  T_2613;
  wire [1:0] T_2619_0;
  wire [1:0] T_2619_1;
  wire [1:0] T_2619_2;
  wire  T_2621;
  wire  T_2622;
  wire  T_2623;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire [3:0] GEN_12;
  wire [1:0] GEN_13;
  wire  T_2630;
  wire [3:0] GEN_14;
  wire [3:0] GEN_20;
  wire [1:0] GEN_21;
  wire  T_2632;
  wire [1:0] T_2638_0;
  wire  T_2640;
  wire [3:0] T_2643;
  wire [3:0] GEN_23;
  wire [39:0] GEN_24;
  wire [8:0] GEN_25;
  wire [4:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [4:0] GEN_29;
  wire  GEN_30;
  wire [19:0] GEN_31;
  wire [1:0] GEN_32;
  wire [3:0] GEN_33;
  wire [3:0] GEN_39;
  wire [1:0] GEN_40;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_2671;
  wire  can_finish;
  wire [3:0] GEN_53;
  wire  T_2676;
  wire  T_2677;
  wire  T_2679;
  wire  T_2681;
  wire  T_2682;
  wire [2:0] T_2709_manager_xact_id;
  wire  T_2709_manager_id;
  wire  T_2735;
  wire  T_2736;
  wire  T_2737;
  wire  T_2738;
  wire [8:0] T_2739;
  wire [11:0] GEN_54;
  wire [11:0] T_2740;
  wire [27:0] T_2741;
  wire  T_2743;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_59;
  wire [1:0] GEN_55;
  wire  T_2746;
  wire [1:0] GEN_56;
  wire [2:0] T_2748;
  wire [1:0] T_2749;
  wire [1:0] GEN_42;
  wire  T_2750;
  wire [1:0] GEN_43;
  wire  T_2753;
  wire  T_2762;
  wire  T_2764;
  wire  T_2765;
  wire  T_2766;
  wire  T_2769;
  wire [1:0] T_2776_0;
  wire [1:0] T_2776_1;
  wire [1:0] T_2817_state;
  wire [1:0] T_2842_state;
  wire  T_2867;
  wire [25:0] T_2869;
  wire [1:0] T_2878_0;
  wire  T_2880;
  wire [2:0] T_2883;
  wire [2:0] T_2922_addr_beat;
  wire [25:0] T_2922_addr_block;
  wire [1:0] T_2922_client_xact_id;
  wire  T_2922_voluntary;
  wire [2:0] T_2922_r_type;
  wire [63:0] T_2922_data;
  wire  T_2953;
  wire [25:0] T_2954;
  wire [5:0] T_2970;
  wire [25:0] T_3004_addr_block;
  wire [1:0] T_3004_client_xact_id;
  wire [2:0] T_3004_addr_beat;
  wire  T_3004_is_builtin_type;
  wire [2:0] T_3004_a_type;
  wire [11:0] T_3004_union;
  wire [63:0] T_3004_data;
  wire  T_3037;
  wire [5:0] T_3039;
  wire [31:0] T_3041;
  wire  T_3043;
  wire  GEN_44;
  wire [4:0] GEN_45;
  reg [3:0] GEN_15;
  reg [31:0] GEN_60;
  Queue_73 rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue_74 fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2447;
  assign io_req_sec_rdy = T_2743;
  assign io_idx_match = T_2738;
  assign io_tag = T_2741[19:0];
  assign io_mem_req_valid = T_2953;
  assign io_mem_req_bits_addr_block = T_3004_addr_block;
  assign io_mem_req_bits_client_xact_id = T_3004_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_3004_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_3004_is_builtin_type;
  assign io_mem_req_bits_a_type = T_3004_a_type;
  assign io_mem_req_bits_union = T_3004_union;
  assign io_mem_req_bits_data = T_3004_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2740;
  assign io_meta_read_valid = T_2445;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_15;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2769;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2842_state;
  assign io_replay_valid = T_3037;
  assign io_replay_bits_addr = {{8'd0}, T_3041};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_45;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2735;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2867;
  assign io_wb_req_bits_addr_beat = T_2922_addr_beat;
  assign io_wb_req_bits_addr_block = T_2922_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2922_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2922_voluntary;
  assign io_wb_req_bits_r_type = T_2922_r_type;
  assign io_wb_req_bits_data = T_2922_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2766;
  assign T_1875_state = {{1'd0}, 1'h0};
  assign req_idx = req_addr[11:6];
  assign T_2271 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2271;
  assign T_2272 = io_req_bits_cmd == 5'h1;
  assign T_2273 = io_req_bits_cmd == 5'h7;
  assign T_2274 = T_2272 | T_2273;
  assign T_2275 = io_req_bits_cmd[3];
  assign T_2276 = io_req_bits_cmd == 5'h4;
  assign T_2277 = T_2275 | T_2276;
  assign T_2278 = T_2274 | T_2277;
  assign T_2279 = io_req_bits_cmd == 5'h3;
  assign T_2280 = T_2278 | T_2279;
  assign T_2281 = io_req_bits_cmd == 5'h6;
  assign T_2282 = T_2280 | T_2281;
  assign T_2283 = req_cmd == 5'h1;
  assign T_2284 = req_cmd == 5'h7;
  assign T_2285 = T_2283 | T_2284;
  assign T_2286 = req_cmd[3];
  assign T_2287 = req_cmd == 5'h4;
  assign T_2288 = T_2286 | T_2287;
  assign T_2289 = T_2285 | T_2288;
  assign T_2290 = req_cmd == 5'h3;
  assign T_2291 = T_2289 | T_2290;
  assign T_2292 = req_cmd == 5'h6;
  assign T_2293 = T_2291 | T_2292;
  assign T_2295 = T_2293 == 1'h0;
  assign cmd_requires_second_acquire = T_2282 & T_2295;
  assign states_before_refill_0 = 4'h1;
  assign states_before_refill_1 = 4'h2;
  assign states_before_refill_2 = 4'h3;
  assign T_2302 = states_before_refill_0 == state;
  assign T_2303 = states_before_refill_1 == state;
  assign T_2304 = states_before_refill_2 == state;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2314_0 = 4'h4;
  assign T_2314_1 = 4'h5;
  assign T_2316 = T_2314_0 == state;
  assign T_2317 = T_2314_1 == state;
  assign T_2320 = T_2316 | T_2317;
  assign T_2322 = cmd_requires_second_acquire == 1'h0;
  assign T_2323 = T_2320 & T_2322;
  assign T_2324 = T_2308 | T_2323;
  assign sec_rdy = idx_match & T_2324;
  assign T_2332_0 = 3'h5;
  assign GEN_46 = {{1'd0}, T_2332_0};
  assign T_2334 = GEN_46 == io_mem_grant_bits_g_type;
  assign T_2342_0 = 2'h0;
  assign T_2342_1 = 2'h1;
  assign GEN_47 = {{2'd0}, T_2342_0};
  assign T_2344 = GEN_47 == io_mem_grant_bits_g_type;
  assign GEN_48 = {{2'd0}, T_2342_1};
  assign T_2345 = GEN_48 == io_mem_grant_bits_g_type;
  assign T_2348 = T_2344 | T_2345;
  assign T_2349 = io_mem_grant_bits_is_builtin_type ? T_2334 : T_2348;
  assign T_2350 = io_mem_grant_valid & T_2349;
  assign T_2353 = refill_cnt == 3'h7;
  assign GEN_49 = {{2'd0}, 1'h1};
  assign T_2355 = refill_cnt + GEN_49;
  assign T_2356 = T_2355[2:0];
  assign GEN_0 = T_2350 ? T_2356 : refill_cnt;
  assign refill_count_done = T_2350 & T_2353;
  assign T_2358 = T_2349 == 1'h0;
  assign T_2359 = T_2358 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2359;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2444;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_44;
  assign T_2436 = io_req_pri_val & io_req_pri_rdy;
  assign T_2437 = io_req_sec_val & sec_rdy;
  assign T_2438 = T_2436 | T_2437;
  assign T_2439 = io_req_bits_cmd == 5'h2;
  assign T_2441 = T_2439 | T_2279;
  assign T_2443 = T_2441 == 1'h0;
  assign T_2444 = T_2438 & T_2443;
  assign T_2445 = state == 4'h8;
  assign T_2446 = io_replay_ready & T_2445;
  assign T_2447 = state == 4'h0;
  assign T_2448 = T_2446 | T_2447;
  assign T_2456 = T_2289 ? 2'h3 : 2'h2;
  assign GEN_50 = {{2'd0}, 2'h2};
  assign T_2457 = GEN_50 == io_mem_grant_bits_g_type;
  assign T_2458 = T_2457 ? 2'h3 : 2'h0;
  assign GEN_51 = {{2'd0}, 2'h1};
  assign T_2459 = GEN_51 == io_mem_grant_bits_g_type;
  assign T_2460 = T_2459 ? T_2456 : T_2458;
  assign GEN_52 = {{2'd0}, 2'h0};
  assign T_2461 = GEN_52 == io_mem_grant_bits_g_type;
  assign T_2462 = T_2461 ? 2'h1 : T_2460;
  assign T_2463 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2462;
  assign coh_on_grant_state = T_2463;
  assign T_2520 = T_2278 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2520;
  assign T_2572 = rpq_io_deq_valid == 1'h0;
  assign T_2573 = T_2445 & T_2572;
  assign GEN_1 = T_2573 ? 4'h0 : state;
  assign T_2574 = state == 4'h7;
  assign GEN_2 = T_2574 ? 4'h8 : GEN_1;
  assign T_2575 = state == 4'h6;
  assign T_2576 = T_2575 & io_meta_write_ready;
  assign GEN_3 = T_2576 ? 4'h7 : GEN_2;
  assign T_2577 = state == 4'h5;
  assign T_2578 = T_2577 & refill_done;
  assign GEN_4 = T_2578 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2578 ? coh_on_grant_state : new_coh_state_state;
  assign T_2579 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2579 ? 4'h5 : GEN_4;
  assign T_2580 = state == 4'h3;
  assign T_2581 = T_2580 & io_meta_write_ready;
  assign GEN_7 = T_2581 ? 4'h4 : GEN_6;
  assign T_2582 = state == 4'h2;
  assign T_2583 = T_2582 & io_mem_grant_valid;
  assign GEN_8 = T_2583 ? 4'h3 : GEN_7;
  assign T_2584 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2584 ? 4'h2 : GEN_8;
  assign T_2589 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign GEN_11 = T_2589 ? GEN_10 : req_cmd;
  assign T_2607_0 = 2'h2;
  assign T_2607_1 = 2'h3;
  assign T_2609 = T_2607_0 == io_req_bits_old_meta_coh_state;
  assign T_2610 = T_2607_1 == io_req_bits_old_meta_coh_state;
  assign T_2613 = T_2609 | T_2610;
  assign T_2619_0 = 2'h1;
  assign T_2619_1 = 2'h2;
  assign T_2619_2 = 2'h3;
  assign T_2621 = T_2619_0 == io_req_bits_old_meta_coh_state;
  assign T_2622 = T_2619_1 == io_req_bits_old_meta_coh_state;
  assign T_2623 = T_2619_2 == io_req_bits_old_meta_coh_state;
  assign T_2626 = T_2621 | T_2622;
  assign T_2627 = T_2626 | T_2623;
  assign T_2628 = T_2282 ? T_2613 : T_2627;
  assign GEN_12 = T_2628 ? 4'h6 : GEN_9;
  assign GEN_13 = T_2628 ? coh_on_hit_state : GEN_5;
  assign T_2630 = T_2628 == 1'h0;
  assign GEN_14 = T_2630 ? 4'h4 : GEN_12;
  assign GEN_20 = io_req_bits_tag_match ? GEN_14 : GEN_9;
  assign GEN_21 = io_req_bits_tag_match ? GEN_13 : GEN_5;
  assign T_2632 = io_req_bits_tag_match == 1'h0;
  assign T_2638_0 = 2'h3;
  assign T_2640 = T_2638_0 == io_req_bits_old_meta_coh_state;
  assign T_2643 = T_2640 ? 4'h1 : 4'h3;
  assign GEN_23 = T_2632 ? T_2643 : GEN_20;
  assign GEN_24 = T_2436 ? io_req_bits_addr : req_addr;
  assign GEN_25 = T_2436 ? io_req_bits_tag : req_tag;
  assign GEN_26 = T_2436 ? io_req_bits_cmd : GEN_11;
  assign GEN_27 = T_2436 ? io_req_bits_typ : req_typ;
  assign GEN_28 = T_2436 ? io_req_bits_phys : req_phys;
  assign GEN_29 = T_2436 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_30 = T_2436 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_31 = T_2436 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_32 = T_2436 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_33 = T_2436 ? io_req_bits_way_en : req_way_en;
  assign GEN_39 = T_2436 ? GEN_23 : GEN_9;
  assign GEN_40 = T_2436 ? GEN_21 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2682;
  assign fq_io_enq_bits_manager_xact_id = T_2709_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2709_manager_id;
  assign fq_io_deq_ready = T_2736;
  assign T_2671 = state == 4'h4;
  assign can_finish = T_2447 | T_2671;
  assign GEN_53 = {{1'd0}, 3'h0};
  assign T_2676 = io_mem_grant_bits_g_type == GEN_53;
  assign T_2677 = io_mem_grant_bits_is_builtin_type & T_2676;
  assign T_2679 = T_2677 == 1'h0;
  assign T_2681 = io_mem_grant_valid & T_2679;
  assign T_2682 = T_2681 & refill_done;
  assign T_2709_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2709_manager_id = io_mem_grant_bits_manager_id;
  assign T_2735 = fq_io_deq_valid & can_finish;
  assign T_2736 = io_mem_finish_ready & can_finish;
  assign T_2737 = state != 4'h0;
  assign T_2738 = T_2737 & idx_match;
  assign T_2739 = {req_idx,refill_cnt};
  assign GEN_54 = {{3'd0}, T_2739};
  assign T_2740 = GEN_54 << 3;
  assign T_2741 = req_addr[39:12];
  assign T_2743 = sec_rdy & rpq_io_enq_ready;
  assign GEN_55 = {{1'd0}, 1'h0};
  assign T_2746 = meta_hazard != GEN_55;
  assign GEN_56 = {{1'd0}, 1'h1};
  assign T_2748 = meta_hazard + GEN_56;
  assign T_2749 = T_2748[1:0];
  assign GEN_42 = T_2746 ? T_2749 : meta_hazard;
  assign T_2750 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_43 = T_2750 ? {{1'd0}, 1'h1} : GEN_42;
  assign T_2753 = idx_match == 1'h0;
  assign T_2762 = T_2308 == 1'h0;
  assign T_2764 = meta_hazard == GEN_55;
  assign T_2765 = T_2762 & T_2764;
  assign T_2766 = T_2753 | T_2765;
  assign T_2769 = T_2575 | T_2580;
  assign T_2776_0 = 2'h2;
  assign T_2776_1 = 2'h3;
  assign T_2817_state = 2'h0;
  assign T_2842_state = T_2580 ? T_2817_state : new_coh_state_state;
  assign T_2867 = state == 4'h1;
  assign T_2869 = {req_old_meta_tag,req_idx};
  assign T_2878_0 = 2'h3;
  assign T_2880 = T_2878_0 == req_old_meta_coh_state;
  assign T_2883 = T_2880 ? 3'h0 : 3'h3;
  assign T_2922_addr_beat = {{2'd0}, 1'h0};
  assign T_2922_addr_block = T_2869;
  assign T_2922_client_xact_id = {{1'd0}, 1'h0};
  assign T_2922_voluntary = 1'h1;
  assign T_2922_r_type = T_2883;
  assign T_2922_data = {{63'd0}, 1'h0};
  assign T_2953 = T_2671 & fq_io_enq_ready;
  assign T_2954 = {io_tag,req_idx};
  assign T_2970 = {req_cmd,1'h1};
  assign T_3004_addr_block = T_2954;
  assign T_3004_client_xact_id = {{1'd0}, 1'h0};
  assign T_3004_addr_beat = {{2'd0}, 1'h0};
  assign T_3004_is_builtin_type = 1'h0;
  assign T_3004_a_type = {{2'd0}, T_2293};
  assign T_3004_union = {{6'd0}, T_2970};
  assign T_3004_data = {{63'd0}, 1'h0};
  assign T_3037 = T_2445 & rpq_io_deq_valid;
  assign T_3039 = rpq_io_deq_bits_addr[5:0];
  assign T_3041 = {T_2954,T_3039};
  assign T_3043 = io_meta_read_ready == 1'h0;
  assign GEN_44 = T_3043 ? 1'h0 : T_2448;
  assign GEN_45 = T_3043 ? 5'h5 : rpq_io_deq_bits_cmd;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_16 = {1{$random}};
  state = GEN_16[3:0];
  GEN_17 = {1{$random}};
  new_coh_state_state = GEN_17[1:0];
  GEN_18 = {2{$random}};
  req_addr = GEN_18[39:0];
  GEN_19 = {1{$random}};
  req_tag = GEN_19[8:0];
  GEN_22 = {1{$random}};
  req_cmd = GEN_22[4:0];
  GEN_34 = {1{$random}};
  req_typ = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_phys = GEN_35[0:0];
  GEN_36 = {1{$random}};
  req_sdq_id = GEN_36[4:0];
  GEN_37 = {1{$random}};
  req_tag_match = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_old_meta_tag = GEN_38[19:0];
  GEN_41 = {1{$random}};
  req_old_meta_coh_state = GEN_41[1:0];
  GEN_57 = {1{$random}};
  req_way_en = GEN_57[3:0];
  GEN_58 = {1{$random}};
  refill_cnt = GEN_58[2:0];
  GEN_59 = {1{$random}};
  meta_hazard = GEN_59[1:0];
  GEN_60 = {1{$random}};
  GEN_15 = GEN_60[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      state <= GEN_39;
    end
    if(reset) begin
      new_coh_state_state <= T_1875_state;
    end else begin
      new_coh_state_state <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      req_addr <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      req_tag <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      req_cmd <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      req_typ <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      req_phys <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      req_sdq_id <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      req_tag_match <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      req_old_meta_tag <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      req_old_meta_coh_state <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      req_way_en <= GEN_33;
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      refill_cnt <= GEN_0;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      meta_hazard <= GEN_43;
    end
  end
endmodule
module MSHR_75(
  input   clk,
  input   reset,
  input   io_req_pri_val,
  output  io_req_pri_rdy,
  input   io_req_sec_val,
  output  io_req_sec_rdy,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [4:0] io_req_bits_sdq_id,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  output  io_idx_match,
  output [19:0] io_tag,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [4:0] io_replay_bits_sdq_id,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy
);
  reg [3:0] state;
  reg [31:0] GEN_16;
  wire [1:0] T_1875_state;
  reg [1:0] new_coh_state_state;
  reg [31:0] GEN_17;
  reg [39:0] req_addr;
  reg [63:0] GEN_18;
  reg [8:0] req_tag;
  reg [31:0] GEN_19;
  reg [4:0] req_cmd;
  reg [31:0] GEN_22;
  reg [2:0] req_typ;
  reg [31:0] GEN_34;
  reg  req_phys;
  reg [31:0] GEN_35;
  reg [4:0] req_sdq_id;
  reg [31:0] GEN_36;
  reg  req_tag_match;
  reg [31:0] GEN_37;
  reg [19:0] req_old_meta_tag;
  reg [31:0] GEN_38;
  reg [1:0] req_old_meta_coh_state;
  reg [31:0] GEN_41;
  reg [3:0] req_way_en;
  reg [31:0] GEN_57;
  wire [5:0] req_idx;
  wire [5:0] T_2271;
  wire  idx_match;
  wire  T_2272;
  wire  T_2273;
  wire  T_2274;
  wire  T_2275;
  wire  T_2276;
  wire  T_2277;
  wire  T_2278;
  wire  T_2279;
  wire  T_2280;
  wire  T_2281;
  wire  T_2282;
  wire  T_2283;
  wire  T_2284;
  wire  T_2285;
  wire  T_2286;
  wire  T_2287;
  wire  T_2288;
  wire  T_2289;
  wire  T_2290;
  wire  T_2291;
  wire  T_2292;
  wire  T_2293;
  wire  T_2295;
  wire  cmd_requires_second_acquire;
  wire [3:0] states_before_refill_0;
  wire [3:0] states_before_refill_1;
  wire [3:0] states_before_refill_2;
  wire  T_2302;
  wire  T_2303;
  wire  T_2304;
  wire  T_2307;
  wire  T_2308;
  wire [3:0] T_2314_0;
  wire [3:0] T_2314_1;
  wire  T_2316;
  wire  T_2317;
  wire  T_2320;
  wire  T_2322;
  wire  T_2323;
  wire  T_2324;
  wire  sec_rdy;
  wire [2:0] T_2332_0;
  wire [3:0] GEN_46;
  wire  T_2334;
  wire [1:0] T_2342_0;
  wire [1:0] T_2342_1;
  wire [3:0] GEN_47;
  wire  T_2344;
  wire [3:0] GEN_48;
  wire  T_2345;
  wire  T_2348;
  wire  T_2349;
  wire  T_2350;
  reg [2:0] refill_cnt;
  reg [31:0] GEN_58;
  wire  T_2353;
  wire [2:0] GEN_49;
  wire [3:0] T_2355;
  wire [2:0] T_2356;
  wire [2:0] GEN_0;
  wire  refill_count_done;
  wire  T_2358;
  wire  T_2359;
  wire  refill_done;
  wire  rpq_clk;
  wire  rpq_reset;
  wire  rpq_io_enq_ready;
  wire  rpq_io_enq_valid;
  wire [39:0] rpq_io_enq_bits_addr;
  wire [8:0] rpq_io_enq_bits_tag;
  wire [4:0] rpq_io_enq_bits_cmd;
  wire [2:0] rpq_io_enq_bits_typ;
  wire  rpq_io_enq_bits_phys;
  wire [4:0] rpq_io_enq_bits_sdq_id;
  wire  rpq_io_deq_ready;
  wire  rpq_io_deq_valid;
  wire [39:0] rpq_io_deq_bits_addr;
  wire [8:0] rpq_io_deq_bits_tag;
  wire [4:0] rpq_io_deq_bits_cmd;
  wire [2:0] rpq_io_deq_bits_typ;
  wire  rpq_io_deq_bits_phys;
  wire [4:0] rpq_io_deq_bits_sdq_id;
  wire [4:0] rpq_io_count;
  wire  T_2436;
  wire  T_2437;
  wire  T_2438;
  wire  T_2439;
  wire  T_2441;
  wire  T_2443;
  wire  T_2444;
  wire  T_2445;
  wire  T_2446;
  wire  T_2447;
  wire  T_2448;
  wire [1:0] T_2456;
  wire [3:0] GEN_50;
  wire  T_2457;
  wire [1:0] T_2458;
  wire [3:0] GEN_51;
  wire  T_2459;
  wire [1:0] T_2460;
  wire [3:0] GEN_52;
  wire  T_2461;
  wire [1:0] T_2462;
  wire [1:0] T_2463;
  wire [1:0] coh_on_grant_state;
  wire [1:0] T_2520;
  wire [1:0] coh_on_hit_state;
  wire  T_2572;
  wire  T_2573;
  wire [3:0] GEN_1;
  wire  T_2574;
  wire [3:0] GEN_2;
  wire  T_2575;
  wire  T_2576;
  wire [3:0] GEN_3;
  wire  T_2577;
  wire  T_2578;
  wire [3:0] GEN_4;
  wire [1:0] GEN_5;
  wire  T_2579;
  wire [3:0] GEN_6;
  wire  T_2580;
  wire  T_2581;
  wire [3:0] GEN_7;
  wire  T_2582;
  wire  T_2583;
  wire [3:0] GEN_8;
  wire  T_2584;
  wire [3:0] GEN_9;
  wire  T_2589;
  wire [4:0] GEN_10;
  wire [4:0] GEN_11;
  wire [1:0] T_2607_0;
  wire [1:0] T_2607_1;
  wire  T_2609;
  wire  T_2610;
  wire  T_2613;
  wire [1:0] T_2619_0;
  wire [1:0] T_2619_1;
  wire [1:0] T_2619_2;
  wire  T_2621;
  wire  T_2622;
  wire  T_2623;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire [3:0] GEN_12;
  wire [1:0] GEN_13;
  wire  T_2630;
  wire [3:0] GEN_14;
  wire [3:0] GEN_20;
  wire [1:0] GEN_21;
  wire  T_2632;
  wire [1:0] T_2638_0;
  wire  T_2640;
  wire [3:0] T_2643;
  wire [3:0] GEN_23;
  wire [39:0] GEN_24;
  wire [8:0] GEN_25;
  wire [4:0] GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [4:0] GEN_29;
  wire  GEN_30;
  wire [19:0] GEN_31;
  wire [1:0] GEN_32;
  wire [3:0] GEN_33;
  wire [3:0] GEN_39;
  wire [1:0] GEN_40;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  wire  T_2671;
  wire  can_finish;
  wire [3:0] GEN_53;
  wire  T_2676;
  wire  T_2677;
  wire  T_2679;
  wire  T_2681;
  wire  T_2682;
  wire [2:0] T_2709_manager_xact_id;
  wire  T_2709_manager_id;
  wire  T_2735;
  wire  T_2736;
  wire  T_2737;
  wire  T_2738;
  wire [8:0] T_2739;
  wire [11:0] GEN_54;
  wire [11:0] T_2740;
  wire [27:0] T_2741;
  wire  T_2743;
  reg [1:0] meta_hazard;
  reg [31:0] GEN_59;
  wire [1:0] GEN_55;
  wire  T_2746;
  wire [1:0] GEN_56;
  wire [2:0] T_2748;
  wire [1:0] T_2749;
  wire [1:0] GEN_42;
  wire  T_2750;
  wire [1:0] GEN_43;
  wire  T_2753;
  wire  T_2762;
  wire  T_2764;
  wire  T_2765;
  wire  T_2766;
  wire  T_2769;
  wire [1:0] T_2776_0;
  wire [1:0] T_2776_1;
  wire [1:0] T_2817_state;
  wire [1:0] T_2842_state;
  wire  T_2867;
  wire [25:0] T_2869;
  wire [1:0] T_2878_0;
  wire  T_2880;
  wire [2:0] T_2883;
  wire [2:0] T_2922_addr_beat;
  wire [25:0] T_2922_addr_block;
  wire [1:0] T_2922_client_xact_id;
  wire  T_2922_voluntary;
  wire [2:0] T_2922_r_type;
  wire [63:0] T_2922_data;
  wire  T_2953;
  wire [25:0] T_2954;
  wire [5:0] T_2970;
  wire [25:0] T_3004_addr_block;
  wire [1:0] T_3004_client_xact_id;
  wire [2:0] T_3004_addr_beat;
  wire  T_3004_is_builtin_type;
  wire [2:0] T_3004_a_type;
  wire [11:0] T_3004_union;
  wire [63:0] T_3004_data;
  wire  T_3037;
  wire [5:0] T_3039;
  wire [31:0] T_3041;
  wire  T_3043;
  wire  GEN_44;
  wire [4:0] GEN_45;
  reg [3:0] GEN_15;
  reg [31:0] GEN_60;
  Queue_73 rpq (
    .clk(rpq_clk),
    .reset(rpq_reset),
    .io_enq_ready(rpq_io_enq_ready),
    .io_enq_valid(rpq_io_enq_valid),
    .io_enq_bits_addr(rpq_io_enq_bits_addr),
    .io_enq_bits_tag(rpq_io_enq_bits_tag),
    .io_enq_bits_cmd(rpq_io_enq_bits_cmd),
    .io_enq_bits_typ(rpq_io_enq_bits_typ),
    .io_enq_bits_phys(rpq_io_enq_bits_phys),
    .io_enq_bits_sdq_id(rpq_io_enq_bits_sdq_id),
    .io_deq_ready(rpq_io_deq_ready),
    .io_deq_valid(rpq_io_deq_valid),
    .io_deq_bits_addr(rpq_io_deq_bits_addr),
    .io_deq_bits_tag(rpq_io_deq_bits_tag),
    .io_deq_bits_cmd(rpq_io_deq_bits_cmd),
    .io_deq_bits_typ(rpq_io_deq_bits_typ),
    .io_deq_bits_phys(rpq_io_deq_bits_phys),
    .io_deq_bits_sdq_id(rpq_io_deq_bits_sdq_id),
    .io_count(rpq_io_count)
  );
  FinishQueue_74 fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_pri_rdy = T_2447;
  assign io_req_sec_rdy = T_2743;
  assign io_idx_match = T_2738;
  assign io_tag = T_2741[19:0];
  assign io_mem_req_valid = T_2953;
  assign io_mem_req_bits_addr_block = T_3004_addr_block;
  assign io_mem_req_bits_client_xact_id = T_3004_client_xact_id;
  assign io_mem_req_bits_addr_beat = T_3004_addr_beat;
  assign io_mem_req_bits_is_builtin_type = T_3004_is_builtin_type;
  assign io_mem_req_bits_a_type = T_3004_a_type;
  assign io_mem_req_bits_union = T_3004_union;
  assign io_mem_req_bits_data = T_3004_data;
  assign io_refill_way_en = req_way_en;
  assign io_refill_addr = T_2740;
  assign io_meta_read_valid = T_2445;
  assign io_meta_read_bits_idx = req_idx;
  assign io_meta_read_bits_way_en = GEN_15;
  assign io_meta_read_bits_tag = io_tag;
  assign io_meta_write_valid = T_2769;
  assign io_meta_write_bits_idx = req_idx;
  assign io_meta_write_bits_way_en = req_way_en;
  assign io_meta_write_bits_data_tag = io_tag;
  assign io_meta_write_bits_data_coh_state = T_2842_state;
  assign io_replay_valid = T_3037;
  assign io_replay_bits_addr = {{8'd0}, T_3041};
  assign io_replay_bits_tag = rpq_io_deq_bits_tag;
  assign io_replay_bits_cmd = GEN_45;
  assign io_replay_bits_typ = rpq_io_deq_bits_typ;
  assign io_replay_bits_phys = 1'h1;
  assign io_replay_bits_sdq_id = rpq_io_deq_bits_sdq_id;
  assign io_mem_finish_valid = T_2735;
  assign io_mem_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_wb_req_valid = T_2867;
  assign io_wb_req_bits_addr_beat = T_2922_addr_beat;
  assign io_wb_req_bits_addr_block = T_2922_addr_block;
  assign io_wb_req_bits_client_xact_id = T_2922_client_xact_id;
  assign io_wb_req_bits_voluntary = T_2922_voluntary;
  assign io_wb_req_bits_r_type = T_2922_r_type;
  assign io_wb_req_bits_data = T_2922_data;
  assign io_wb_req_bits_way_en = req_way_en;
  assign io_probe_rdy = T_2766;
  assign T_1875_state = {{1'd0}, 1'h0};
  assign req_idx = req_addr[11:6];
  assign T_2271 = io_req_bits_addr[11:6];
  assign idx_match = req_idx == T_2271;
  assign T_2272 = io_req_bits_cmd == 5'h1;
  assign T_2273 = io_req_bits_cmd == 5'h7;
  assign T_2274 = T_2272 | T_2273;
  assign T_2275 = io_req_bits_cmd[3];
  assign T_2276 = io_req_bits_cmd == 5'h4;
  assign T_2277 = T_2275 | T_2276;
  assign T_2278 = T_2274 | T_2277;
  assign T_2279 = io_req_bits_cmd == 5'h3;
  assign T_2280 = T_2278 | T_2279;
  assign T_2281 = io_req_bits_cmd == 5'h6;
  assign T_2282 = T_2280 | T_2281;
  assign T_2283 = req_cmd == 5'h1;
  assign T_2284 = req_cmd == 5'h7;
  assign T_2285 = T_2283 | T_2284;
  assign T_2286 = req_cmd[3];
  assign T_2287 = req_cmd == 5'h4;
  assign T_2288 = T_2286 | T_2287;
  assign T_2289 = T_2285 | T_2288;
  assign T_2290 = req_cmd == 5'h3;
  assign T_2291 = T_2289 | T_2290;
  assign T_2292 = req_cmd == 5'h6;
  assign T_2293 = T_2291 | T_2292;
  assign T_2295 = T_2293 == 1'h0;
  assign cmd_requires_second_acquire = T_2282 & T_2295;
  assign states_before_refill_0 = 4'h1;
  assign states_before_refill_1 = 4'h2;
  assign states_before_refill_2 = 4'h3;
  assign T_2302 = states_before_refill_0 == state;
  assign T_2303 = states_before_refill_1 == state;
  assign T_2304 = states_before_refill_2 == state;
  assign T_2307 = T_2302 | T_2303;
  assign T_2308 = T_2307 | T_2304;
  assign T_2314_0 = 4'h4;
  assign T_2314_1 = 4'h5;
  assign T_2316 = T_2314_0 == state;
  assign T_2317 = T_2314_1 == state;
  assign T_2320 = T_2316 | T_2317;
  assign T_2322 = cmd_requires_second_acquire == 1'h0;
  assign T_2323 = T_2320 & T_2322;
  assign T_2324 = T_2308 | T_2323;
  assign sec_rdy = idx_match & T_2324;
  assign T_2332_0 = 3'h5;
  assign GEN_46 = {{1'd0}, T_2332_0};
  assign T_2334 = GEN_46 == io_mem_grant_bits_g_type;
  assign T_2342_0 = 2'h0;
  assign T_2342_1 = 2'h1;
  assign GEN_47 = {{2'd0}, T_2342_0};
  assign T_2344 = GEN_47 == io_mem_grant_bits_g_type;
  assign GEN_48 = {{2'd0}, T_2342_1};
  assign T_2345 = GEN_48 == io_mem_grant_bits_g_type;
  assign T_2348 = T_2344 | T_2345;
  assign T_2349 = io_mem_grant_bits_is_builtin_type ? T_2334 : T_2348;
  assign T_2350 = io_mem_grant_valid & T_2349;
  assign T_2353 = refill_cnt == 3'h7;
  assign GEN_49 = {{2'd0}, 1'h1};
  assign T_2355 = refill_cnt + GEN_49;
  assign T_2356 = T_2355[2:0];
  assign GEN_0 = T_2350 ? T_2356 : refill_cnt;
  assign refill_count_done = T_2350 & T_2353;
  assign T_2358 = T_2349 == 1'h0;
  assign T_2359 = T_2358 | refill_count_done;
  assign refill_done = io_mem_grant_valid & T_2359;
  assign rpq_clk = clk;
  assign rpq_reset = reset;
  assign rpq_io_enq_valid = T_2444;
  assign rpq_io_enq_bits_addr = io_req_bits_addr;
  assign rpq_io_enq_bits_tag = io_req_bits_tag;
  assign rpq_io_enq_bits_cmd = io_req_bits_cmd;
  assign rpq_io_enq_bits_typ = io_req_bits_typ;
  assign rpq_io_enq_bits_phys = io_req_bits_phys;
  assign rpq_io_enq_bits_sdq_id = io_req_bits_sdq_id;
  assign rpq_io_deq_ready = GEN_44;
  assign T_2436 = io_req_pri_val & io_req_pri_rdy;
  assign T_2437 = io_req_sec_val & sec_rdy;
  assign T_2438 = T_2436 | T_2437;
  assign T_2439 = io_req_bits_cmd == 5'h2;
  assign T_2441 = T_2439 | T_2279;
  assign T_2443 = T_2441 == 1'h0;
  assign T_2444 = T_2438 & T_2443;
  assign T_2445 = state == 4'h8;
  assign T_2446 = io_replay_ready & T_2445;
  assign T_2447 = state == 4'h0;
  assign T_2448 = T_2446 | T_2447;
  assign T_2456 = T_2289 ? 2'h3 : 2'h2;
  assign GEN_50 = {{2'd0}, 2'h2};
  assign T_2457 = GEN_50 == io_mem_grant_bits_g_type;
  assign T_2458 = T_2457 ? 2'h3 : 2'h0;
  assign GEN_51 = {{2'd0}, 2'h1};
  assign T_2459 = GEN_51 == io_mem_grant_bits_g_type;
  assign T_2460 = T_2459 ? T_2456 : T_2458;
  assign GEN_52 = {{2'd0}, 2'h0};
  assign T_2461 = GEN_52 == io_mem_grant_bits_g_type;
  assign T_2462 = T_2461 ? 2'h1 : T_2460;
  assign T_2463 = io_mem_grant_bits_is_builtin_type ? 2'h0 : T_2462;
  assign coh_on_grant_state = T_2463;
  assign T_2520 = T_2278 ? 2'h3 : io_req_bits_old_meta_coh_state;
  assign coh_on_hit_state = T_2520;
  assign T_2572 = rpq_io_deq_valid == 1'h0;
  assign T_2573 = T_2445 & T_2572;
  assign GEN_1 = T_2573 ? 4'h0 : state;
  assign T_2574 = state == 4'h7;
  assign GEN_2 = T_2574 ? 4'h8 : GEN_1;
  assign T_2575 = state == 4'h6;
  assign T_2576 = T_2575 & io_meta_write_ready;
  assign GEN_3 = T_2576 ? 4'h7 : GEN_2;
  assign T_2577 = state == 4'h5;
  assign T_2578 = T_2577 & refill_done;
  assign GEN_4 = T_2578 ? 4'h6 : GEN_3;
  assign GEN_5 = T_2578 ? coh_on_grant_state : new_coh_state_state;
  assign T_2579 = io_mem_req_ready & io_mem_req_valid;
  assign GEN_6 = T_2579 ? 4'h5 : GEN_4;
  assign T_2580 = state == 4'h3;
  assign T_2581 = T_2580 & io_meta_write_ready;
  assign GEN_7 = T_2581 ? 4'h4 : GEN_6;
  assign T_2582 = state == 4'h2;
  assign T_2583 = T_2582 & io_mem_grant_valid;
  assign GEN_8 = T_2583 ? 4'h3 : GEN_7;
  assign T_2584 = io_wb_req_ready & io_wb_req_valid;
  assign GEN_9 = T_2584 ? 4'h2 : GEN_8;
  assign T_2589 = io_req_sec_val & io_req_sec_rdy;
  assign GEN_10 = cmd_requires_second_acquire ? io_req_bits_cmd : req_cmd;
  assign GEN_11 = T_2589 ? GEN_10 : req_cmd;
  assign T_2607_0 = 2'h2;
  assign T_2607_1 = 2'h3;
  assign T_2609 = T_2607_0 == io_req_bits_old_meta_coh_state;
  assign T_2610 = T_2607_1 == io_req_bits_old_meta_coh_state;
  assign T_2613 = T_2609 | T_2610;
  assign T_2619_0 = 2'h1;
  assign T_2619_1 = 2'h2;
  assign T_2619_2 = 2'h3;
  assign T_2621 = T_2619_0 == io_req_bits_old_meta_coh_state;
  assign T_2622 = T_2619_1 == io_req_bits_old_meta_coh_state;
  assign T_2623 = T_2619_2 == io_req_bits_old_meta_coh_state;
  assign T_2626 = T_2621 | T_2622;
  assign T_2627 = T_2626 | T_2623;
  assign T_2628 = T_2282 ? T_2613 : T_2627;
  assign GEN_12 = T_2628 ? 4'h6 : GEN_9;
  assign GEN_13 = T_2628 ? coh_on_hit_state : GEN_5;
  assign T_2630 = T_2628 == 1'h0;
  assign GEN_14 = T_2630 ? 4'h4 : GEN_12;
  assign GEN_20 = io_req_bits_tag_match ? GEN_14 : GEN_9;
  assign GEN_21 = io_req_bits_tag_match ? GEN_13 : GEN_5;
  assign T_2632 = io_req_bits_tag_match == 1'h0;
  assign T_2638_0 = 2'h3;
  assign T_2640 = T_2638_0 == io_req_bits_old_meta_coh_state;
  assign T_2643 = T_2640 ? 4'h1 : 4'h3;
  assign GEN_23 = T_2632 ? T_2643 : GEN_20;
  assign GEN_24 = T_2436 ? io_req_bits_addr : req_addr;
  assign GEN_25 = T_2436 ? io_req_bits_tag : req_tag;
  assign GEN_26 = T_2436 ? io_req_bits_cmd : GEN_11;
  assign GEN_27 = T_2436 ? io_req_bits_typ : req_typ;
  assign GEN_28 = T_2436 ? io_req_bits_phys : req_phys;
  assign GEN_29 = T_2436 ? io_req_bits_sdq_id : req_sdq_id;
  assign GEN_30 = T_2436 ? io_req_bits_tag_match : req_tag_match;
  assign GEN_31 = T_2436 ? io_req_bits_old_meta_tag : req_old_meta_tag;
  assign GEN_32 = T_2436 ? io_req_bits_old_meta_coh_state : req_old_meta_coh_state;
  assign GEN_33 = T_2436 ? io_req_bits_way_en : req_way_en;
  assign GEN_39 = T_2436 ? GEN_23 : GEN_9;
  assign GEN_40 = T_2436 ? GEN_21 : GEN_5;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_2682;
  assign fq_io_enq_bits_manager_xact_id = T_2709_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_2709_manager_id;
  assign fq_io_deq_ready = T_2736;
  assign T_2671 = state == 4'h4;
  assign can_finish = T_2447 | T_2671;
  assign GEN_53 = {{1'd0}, 3'h0};
  assign T_2676 = io_mem_grant_bits_g_type == GEN_53;
  assign T_2677 = io_mem_grant_bits_is_builtin_type & T_2676;
  assign T_2679 = T_2677 == 1'h0;
  assign T_2681 = io_mem_grant_valid & T_2679;
  assign T_2682 = T_2681 & refill_done;
  assign T_2709_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign T_2709_manager_id = io_mem_grant_bits_manager_id;
  assign T_2735 = fq_io_deq_valid & can_finish;
  assign T_2736 = io_mem_finish_ready & can_finish;
  assign T_2737 = state != 4'h0;
  assign T_2738 = T_2737 & idx_match;
  assign T_2739 = {req_idx,refill_cnt};
  assign GEN_54 = {{3'd0}, T_2739};
  assign T_2740 = GEN_54 << 3;
  assign T_2741 = req_addr[39:12];
  assign T_2743 = sec_rdy & rpq_io_enq_ready;
  assign GEN_55 = {{1'd0}, 1'h0};
  assign T_2746 = meta_hazard != GEN_55;
  assign GEN_56 = {{1'd0}, 1'h1};
  assign T_2748 = meta_hazard + GEN_56;
  assign T_2749 = T_2748[1:0];
  assign GEN_42 = T_2746 ? T_2749 : meta_hazard;
  assign T_2750 = io_meta_write_ready & io_meta_write_valid;
  assign GEN_43 = T_2750 ? {{1'd0}, 1'h1} : GEN_42;
  assign T_2753 = idx_match == 1'h0;
  assign T_2762 = T_2308 == 1'h0;
  assign T_2764 = meta_hazard == GEN_55;
  assign T_2765 = T_2762 & T_2764;
  assign T_2766 = T_2753 | T_2765;
  assign T_2769 = T_2575 | T_2580;
  assign T_2776_0 = 2'h2;
  assign T_2776_1 = 2'h3;
  assign T_2817_state = 2'h0;
  assign T_2842_state = T_2580 ? T_2817_state : new_coh_state_state;
  assign T_2867 = state == 4'h1;
  assign T_2869 = {req_old_meta_tag,req_idx};
  assign T_2878_0 = 2'h3;
  assign T_2880 = T_2878_0 == req_old_meta_coh_state;
  assign T_2883 = T_2880 ? 3'h0 : 3'h3;
  assign T_2922_addr_beat = {{2'd0}, 1'h0};
  assign T_2922_addr_block = T_2869;
  assign T_2922_client_xact_id = {{1'd0}, 1'h1};
  assign T_2922_voluntary = 1'h1;
  assign T_2922_r_type = T_2883;
  assign T_2922_data = {{63'd0}, 1'h0};
  assign T_2953 = T_2671 & fq_io_enq_ready;
  assign T_2954 = {io_tag,req_idx};
  assign T_2970 = {req_cmd,1'h1};
  assign T_3004_addr_block = T_2954;
  assign T_3004_client_xact_id = {{1'd0}, 1'h1};
  assign T_3004_addr_beat = {{2'd0}, 1'h0};
  assign T_3004_is_builtin_type = 1'h0;
  assign T_3004_a_type = {{2'd0}, T_2293};
  assign T_3004_union = {{6'd0}, T_2970};
  assign T_3004_data = {{63'd0}, 1'h0};
  assign T_3037 = T_2445 & rpq_io_deq_valid;
  assign T_3039 = rpq_io_deq_bits_addr[5:0];
  assign T_3041 = {T_2954,T_3039};
  assign T_3043 = io_meta_read_ready == 1'h0;
  assign GEN_44 = T_3043 ? 1'h0 : T_2448;
  assign GEN_45 = T_3043 ? 5'h5 : rpq_io_deq_bits_cmd;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_16 = {1{$random}};
  state = GEN_16[3:0];
  GEN_17 = {1{$random}};
  new_coh_state_state = GEN_17[1:0];
  GEN_18 = {2{$random}};
  req_addr = GEN_18[39:0];
  GEN_19 = {1{$random}};
  req_tag = GEN_19[8:0];
  GEN_22 = {1{$random}};
  req_cmd = GEN_22[4:0];
  GEN_34 = {1{$random}};
  req_typ = GEN_34[2:0];
  GEN_35 = {1{$random}};
  req_phys = GEN_35[0:0];
  GEN_36 = {1{$random}};
  req_sdq_id = GEN_36[4:0];
  GEN_37 = {1{$random}};
  req_tag_match = GEN_37[0:0];
  GEN_38 = {1{$random}};
  req_old_meta_tag = GEN_38[19:0];
  GEN_41 = {1{$random}};
  req_old_meta_coh_state = GEN_41[1:0];
  GEN_57 = {1{$random}};
  req_way_en = GEN_57[3:0];
  GEN_58 = {1{$random}};
  refill_cnt = GEN_58[2:0];
  GEN_59 = {1{$random}};
  meta_hazard = GEN_59[1:0];
  GEN_60 = {1{$random}};
  GEN_15 = GEN_60[3:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 4'h0;
    end else begin
      state <= GEN_39;
    end
    if(reset) begin
      new_coh_state_state <= T_1875_state;
    end else begin
      new_coh_state_state <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      req_addr <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      req_tag <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      req_cmd <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      req_typ <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      req_phys <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      req_sdq_id <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      req_tag_match <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      req_old_meta_tag <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      req_old_meta_coh_state <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      req_way_en <= GEN_33;
    end
    if(reset) begin
      refill_cnt <= 3'h0;
    end else begin
      refill_cnt <= GEN_0;
    end
    if(reset) begin
      meta_hazard <= 2'h0;
    end else begin
      meta_hazard <= GEN_43;
    end
  end
endmodule
module Arbiter_78(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input   io_in_0_bits,
  input   io_out_ready,
  output  io_out_valid,
  output  io_out_bits,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits = io_in_0_bits;
  assign io_chosen = 1'h0;
endmodule
module Arbiter_79(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [39:0] io_in_0_bits_addr,
  input  [8:0] io_in_0_bits_tag,
  input  [4:0] io_in_0_bits_cmd,
  input  [2:0] io_in_0_bits_typ,
  input  [63:0] io_in_0_bits_data,
  input   io_in_0_bits_replay,
  input   io_in_0_bits_has_data,
  input  [63:0] io_in_0_bits_data_word_bypass,
  input  [63:0] io_in_0_bits_store_data,
  input   io_out_ready,
  output  io_out_valid,
  output [39:0] io_out_bits_addr,
  output [8:0] io_out_bits_tag,
  output [4:0] io_out_bits_cmd,
  output [2:0] io_out_bits_typ,
  output [63:0] io_out_bits_data,
  output  io_out_bits_replay,
  output  io_out_bits_has_data,
  output [63:0] io_out_bits_data_word_bypass,
  output [63:0] io_out_bits_store_data,
  output  io_chosen
);
  assign io_in_0_ready = io_out_ready;
  assign io_out_valid = io_in_0_valid;
  assign io_out_bits_addr = io_in_0_bits_addr;
  assign io_out_bits_tag = io_in_0_bits_tag;
  assign io_out_bits_cmd = io_in_0_bits_cmd;
  assign io_out_bits_typ = io_in_0_bits_typ;
  assign io_out_bits_data = io_in_0_bits_data;
  assign io_out_bits_replay = io_in_0_bits_replay;
  assign io_out_bits_has_data = io_in_0_bits_has_data;
  assign io_out_bits_data_word_bypass = io_in_0_bits_data_word_bypass;
  assign io_out_bits_store_data = io_in_0_bits_store_data;
  assign io_chosen = 1'h0;
endmodule
module IOMSHR(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_acquire_ready,
  output  io_acquire_valid,
  output [25:0] io_acquire_bits_addr_block,
  output [1:0] io_acquire_bits_client_xact_id,
  output [2:0] io_acquire_bits_addr_beat,
  output  io_acquire_bits_is_builtin_type,
  output [2:0] io_acquire_bits_a_type,
  output [11:0] io_acquire_bits_union,
  output [63:0] io_acquire_bits_data,
  input   io_grant_valid,
  input  [2:0] io_grant_bits_addr_beat,
  input  [1:0] io_grant_bits_client_xact_id,
  input  [2:0] io_grant_bits_manager_xact_id,
  input   io_grant_bits_is_builtin_type,
  input  [3:0] io_grant_bits_g_type,
  input  [63:0] io_grant_bits_data,
  input   io_grant_bits_manager_id,
  input   io_finish_ready,
  output  io_finish_valid,
  output [2:0] io_finish_bits_manager_xact_id,
  output  io_finish_bits_manager_id,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [8:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_replay_next
);
  reg [39:0] req_addr;
  reg [63:0] GEN_22;
  reg [8:0] req_tag;
  reg [31:0] GEN_24;
  reg [4:0] req_cmd;
  reg [31:0] GEN_27;
  reg [2:0] req_typ;
  reg [31:0] GEN_28;
  reg  req_phys;
  reg [31:0] GEN_29;
  reg [63:0] req_data;
  reg [63:0] GEN_30;
  wire  req_cmd_sc;
  reg [63:0] grant_word;
  reg [63:0] GEN_31;
  wire  fq_clk;
  wire  fq_reset;
  wire  fq_io_enq_ready;
  wire  fq_io_enq_valid;
  wire [2:0] fq_io_enq_bits_manager_xact_id;
  wire  fq_io_enq_bits_manager_id;
  wire  fq_io_deq_ready;
  wire  fq_io_deq_valid;
  wire [2:0] fq_io_deq_bits_manager_xact_id;
  wire  fq_io_deq_bits_manager_id;
  wire  fq_io_count;
  reg [2:0] state;
  reg [31:0] GEN_32;
  wire  T_1211;
  wire [3:0] GEN_13;
  wire  T_1216;
  wire  T_1217;
  wire  T_1219;
  wire  T_1221;
  wire [2:0] T_1248_manager_xact_id;
  wire  T_1248_manager_id;
  wire  T_1274;
  wire  T_1275;
  wire  T_1277;
  wire [1:0] T_1278;
  wire [2:0] T_1280;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  T_1282;
  wire  T_1284;
  wire [1:0] GEN_16;
  wire  T_1288;
  wire  T_1292;
  wire  T_1295;
  wire [1:0] T_1296;
  wire  T_1297;
  wire [1:0] T_1299;
  wire  T_1301;
  wire [1:0] T_1304;
  wire [1:0] T_1305;
  wire [1:0] T_1308;
  wire [3:0] T_1309;
  wire  T_1310;
  wire [3:0] T_1312;
  wire  T_1314;
  wire [3:0] T_1317;
  wire [3:0] T_1318;
  wire [3:0] T_1321;
  wire [7:0] T_1322;
  wire [22:0] GEN_17;
  wire [22:0] beat_mask;
  wire [1:0] GEN_18;
  wire  T_1327;
  wire [7:0] T_1328;
  wire [15:0] T_1329;
  wire [31:0] T_1330;
  wire [63:0] T_1331;
  wire  T_1333;
  wire [15:0] T_1334;
  wire [31:0] T_1335;
  wire [63:0] T_1336;
  wire  T_1338;
  wire [31:0] T_1339;
  wire [63:0] T_1340;
  wire [63:0] T_1341;
  wire [63:0] T_1342;
  wire [63:0] beat_data;
  wire [25:0] addr_block;
  wire [2:0] addr_beat;
  wire [2:0] addr_byte;
  wire [5:0] T_1387;
  wire [11:0] T_1388;
  wire [25:0] get_acquire_addr_block;
  wire [1:0] get_acquire_client_xact_id;
  wire [2:0] get_acquire_addr_beat;
  wire  get_acquire_is_builtin_type;
  wire [2:0] get_acquire_a_type;
  wire [11:0] get_acquire_union;
  wire [63:0] get_acquire_data;
  wire [22:0] GEN_20;
  wire [22:0] T_1518;
  wire [7:0] T_1519;
  wire [8:0] T_1529;
  wire [11:0] T_1549;
  wire [25:0] put_acquire_addr_block;
  wire [1:0] put_acquire_client_xact_id;
  wire [2:0] put_acquire_addr_beat;
  wire  put_acquire_is_builtin_type;
  wire [2:0] put_acquire_a_type;
  wire [11:0] put_acquire_union;
  wire [63:0] put_acquire_data;
  wire [5:0] T_1657;
  wire [11:0] T_1659;
  wire [25:0] putAtomic_acquire_addr_block;
  wire [1:0] putAtomic_acquire_client_xact_id;
  wire [2:0] putAtomic_acquire_addr_beat;
  wire  putAtomic_acquire_is_builtin_type;
  wire [2:0] putAtomic_acquire_a_type;
  wire [11:0] putAtomic_acquire_union;
  wire [63:0] putAtomic_acquire_data;
  wire  T_1750;
  wire  T_1751;
  wire  T_1752;
  wire  T_1753;
  wire  T_1754;
  wire  T_1755;
  wire  T_1756;
  wire  T_1758;
  wire  T_1762;
  wire [25:0] T_1763_addr_block;
  wire [1:0] T_1763_client_xact_id;
  wire [2:0] T_1763_addr_beat;
  wire  T_1763_is_builtin_type;
  wire [2:0] T_1763_a_type;
  wire [11:0] T_1763_union;
  wire [63:0] T_1763_data;
  wire [25:0] T_1794_addr_block;
  wire [1:0] T_1794_client_xact_id;
  wire [2:0] T_1794_addr_beat;
  wire  T_1794_is_builtin_type;
  wire [2:0] T_1794_a_type;
  wire [11:0] T_1794_union;
  wire [63:0] T_1794_data;
  wire  T_1825;
  wire  T_1827;
  wire  T_1828;
  wire  T_1829;
  wire  T_1830;
  wire [31:0] T_1841;
  wire [31:0] T_1842;
  wire [31:0] T_1843;
  wire  T_1851;
  wire  T_1852;
  wire [31:0] GEN_21;
  wire [32:0] T_1854;
  wire [31:0] T_1855;
  wire [31:0] T_1857;
  wire [63:0] T_1858;
  wire [15:0] T_1860;
  wire [15:0] T_1861;
  wire [15:0] T_1862;
  wire  T_1870;
  wire  T_1871;
  wire [47:0] GEN_23;
  wire [48:0] T_1873;
  wire [47:0] T_1874;
  wire [47:0] T_1875;
  wire [47:0] T_1876;
  wire [63:0] T_1877;
  wire [7:0] T_1879;
  wire [7:0] T_1880;
  wire [7:0] T_1881;
  wire [7:0] T_1885;
  wire  T_1888;
  wire  T_1889;
  wire  T_1890;
  wire [55:0] GEN_25;
  wire [56:0] T_1892;
  wire [55:0] T_1893;
  wire [55:0] T_1894;
  wire [55:0] T_1895;
  wire [63:0] T_1896;
  wire [63:0] GEN_26;
  wire [63:0] T_1897;
  wire  T_1899;
  wire [39:0] GEN_0;
  wire [8:0] GEN_1;
  wire [4:0] GEN_2;
  wire [2:0] GEN_3;
  wire  GEN_4;
  wire [63:0] GEN_5;
  wire [2:0] GEN_6;
  wire  T_1900;
  wire [2:0] GEN_7;
  wire  T_1902;
  wire [63:0] T_1915;
  wire [63:0] GEN_8;
  wire [2:0] GEN_9;
  wire [63:0] GEN_10;
  wire  T_1917;
  wire [2:0] GEN_11;
  wire  T_1918;
  wire [2:0] GEN_12;
  reg [63:0] GEN_19;
  reg [63:0] GEN_33;
  FinishQueue_74 fq (
    .clk(fq_clk),
    .reset(fq_reset),
    .io_enq_ready(fq_io_enq_ready),
    .io_enq_valid(fq_io_enq_valid),
    .io_enq_bits_manager_xact_id(fq_io_enq_bits_manager_xact_id),
    .io_enq_bits_manager_id(fq_io_enq_bits_manager_id),
    .io_deq_ready(fq_io_deq_ready),
    .io_deq_valid(fq_io_deq_valid),
    .io_deq_bits_manager_xact_id(fq_io_deq_bits_manager_xact_id),
    .io_deq_bits_manager_id(fq_io_deq_bits_manager_id),
    .io_count(fq_io_count)
  );
  assign io_req_ready = T_1211;
  assign io_acquire_valid = T_1750;
  assign io_acquire_bits_addr_block = T_1794_addr_block;
  assign io_acquire_bits_client_xact_id = T_1794_client_xact_id;
  assign io_acquire_bits_addr_beat = T_1794_addr_beat;
  assign io_acquire_bits_is_builtin_type = T_1794_is_builtin_type;
  assign io_acquire_bits_a_type = T_1794_a_type;
  assign io_acquire_bits_union = T_1794_union;
  assign io_acquire_bits_data = T_1794_data;
  assign io_finish_valid = T_1275;
  assign io_finish_bits_manager_xact_id = fq_io_deq_bits_manager_xact_id;
  assign io_finish_bits_manager_id = fq_io_deq_bits_manager_id;
  assign io_resp_valid = T_1830;
  assign io_resp_bits_addr = req_addr;
  assign io_resp_bits_tag = req_tag;
  assign io_resp_bits_cmd = req_cmd;
  assign io_resp_bits_typ = req_typ;
  assign io_resp_bits_data = T_1897;
  assign io_resp_bits_replay = 1'h1;
  assign io_resp_bits_has_data = T_1762;
  assign io_resp_bits_data_word_bypass = GEN_19;
  assign io_resp_bits_store_data = req_data;
  assign io_replay_next = T_1829;
  assign req_cmd_sc = req_cmd == 5'h7;
  assign fq_clk = clk;
  assign fq_reset = reset;
  assign fq_io_enq_valid = T_1221;
  assign fq_io_enq_bits_manager_xact_id = T_1248_manager_xact_id;
  assign fq_io_enq_bits_manager_id = T_1248_manager_id;
  assign fq_io_deq_ready = T_1277;
  assign T_1211 = state == 3'h0;
  assign GEN_13 = {{1'd0}, 3'h0};
  assign T_1216 = io_grant_bits_g_type == GEN_13;
  assign T_1217 = io_grant_bits_is_builtin_type & T_1216;
  assign T_1219 = T_1217 == 1'h0;
  assign T_1221 = io_grant_valid & T_1219;
  assign T_1248_manager_xact_id = io_grant_bits_manager_xact_id;
  assign T_1248_manager_id = io_grant_bits_manager_id;
  assign T_1274 = state == 3'h4;
  assign T_1275 = fq_io_deq_valid & T_1274;
  assign T_1277 = io_finish_ready & T_1274;
  assign T_1278 = req_typ[1:0];
  assign T_1280 = $signed(req_typ);
  assign GEN_14 = $signed(1'h0);
  assign GEN_15 = {3{GEN_14}};
  assign T_1282 = $signed(T_1280) >= $signed(GEN_15);
  assign T_1284 = req_addr[0];
  assign GEN_16 = {{1'd0}, 1'h1};
  assign T_1288 = T_1278 >= GEN_16;
  assign T_1292 = T_1284 | T_1288;
  assign T_1295 = T_1284 ? 1'h0 : 1'h1;
  assign T_1296 = {T_1292,T_1295};
  assign T_1297 = req_addr[1];
  assign T_1299 = T_1297 ? T_1296 : {{1'd0}, 1'h0};
  assign T_1301 = T_1278 >= 2'h2;
  assign T_1304 = T_1301 ? 2'h3 : {{1'd0}, 1'h0};
  assign T_1305 = T_1299 | T_1304;
  assign T_1308 = T_1297 ? {{1'd0}, 1'h0} : T_1296;
  assign T_1309 = {T_1305,T_1308};
  assign T_1310 = req_addr[2];
  assign T_1312 = T_1310 ? T_1309 : {{3'd0}, 1'h0};
  assign T_1314 = T_1278 >= 2'h3;
  assign T_1317 = T_1314 ? 4'hf : {{3'd0}, 1'h0};
  assign T_1318 = T_1312 | T_1317;
  assign T_1321 = T_1310 ? {{3'd0}, 1'h0} : T_1309;
  assign T_1322 = {T_1318,T_1321};
  assign GEN_17 = {{15'd0}, T_1322};
  assign beat_mask = GEN_17 << 4'h0;
  assign GEN_18 = {{1'd0}, 1'h0};
  assign T_1327 = T_1278 == GEN_18;
  assign T_1328 = req_data[7:0];
  assign T_1329 = {T_1328,T_1328};
  assign T_1330 = {T_1329,T_1329};
  assign T_1331 = {T_1330,T_1330};
  assign T_1333 = T_1278 == GEN_16;
  assign T_1334 = req_data[15:0];
  assign T_1335 = {T_1334,T_1334};
  assign T_1336 = {T_1335,T_1335};
  assign T_1338 = T_1278 == 2'h2;
  assign T_1339 = req_data[31:0];
  assign T_1340 = {T_1339,T_1339};
  assign T_1341 = T_1338 ? T_1340 : req_data;
  assign T_1342 = T_1333 ? T_1336 : T_1341;
  assign beat_data = T_1327 ? T_1331 : T_1342;
  assign addr_block = req_addr[31:6];
  assign addr_beat = req_addr[5:3];
  assign addr_byte = req_addr[2:0];
  assign T_1387 = {addr_byte,req_typ};
  assign T_1388 = {T_1387,6'h0};
  assign get_acquire_addr_block = addr_block;
  assign get_acquire_client_xact_id = 2'h2;
  assign get_acquire_addr_beat = addr_beat;
  assign get_acquire_is_builtin_type = 1'h1;
  assign get_acquire_a_type = 3'h0;
  assign get_acquire_union = T_1388;
  assign get_acquire_data = {{63'd0}, 1'h0};
  assign GEN_20 = {{15'd0}, 8'h0};
  assign T_1518 = GEN_20 | beat_mask;
  assign T_1519 = T_1518[7:0];
  assign T_1529 = {T_1519,1'h0};
  assign T_1549 = 1'h1 ? {{3'd0}, T_1529} : 12'h0;
  assign put_acquire_addr_block = addr_block;
  assign put_acquire_client_xact_id = 2'h2;
  assign put_acquire_addr_beat = addr_beat;
  assign put_acquire_is_builtin_type = 1'h1;
  assign put_acquire_a_type = 3'h2;
  assign put_acquire_union = T_1549;
  assign put_acquire_data = beat_data;
  assign T_1657 = {req_cmd,1'h1};
  assign T_1659 = {T_1387,T_1657};
  assign putAtomic_acquire_addr_block = addr_block;
  assign putAtomic_acquire_client_xact_id = 2'h2;
  assign putAtomic_acquire_addr_beat = addr_beat;
  assign putAtomic_acquire_is_builtin_type = 1'h1;
  assign putAtomic_acquire_a_type = 3'h4;
  assign putAtomic_acquire_union = T_1659;
  assign putAtomic_acquire_data = beat_data;
  assign T_1750 = state == 3'h1;
  assign T_1751 = req_cmd[3];
  assign T_1752 = req_cmd == 5'h4;
  assign T_1753 = T_1751 | T_1752;
  assign T_1754 = req_cmd == 5'h0;
  assign T_1755 = req_cmd == 5'h6;
  assign T_1756 = T_1754 | T_1755;
  assign T_1758 = T_1756 | req_cmd_sc;
  assign T_1762 = T_1758 | T_1753;
  assign T_1763_addr_block = T_1762 ? get_acquire_addr_block : put_acquire_addr_block;
  assign T_1763_client_xact_id = T_1762 ? get_acquire_client_xact_id : put_acquire_client_xact_id;
  assign T_1763_addr_beat = T_1762 ? get_acquire_addr_beat : put_acquire_addr_beat;
  assign T_1763_is_builtin_type = T_1762 ? get_acquire_is_builtin_type : put_acquire_is_builtin_type;
  assign T_1763_a_type = T_1762 ? get_acquire_a_type : put_acquire_a_type;
  assign T_1763_union = T_1762 ? get_acquire_union : put_acquire_union;
  assign T_1763_data = T_1762 ? get_acquire_data : put_acquire_data;
  assign T_1794_addr_block = T_1753 ? putAtomic_acquire_addr_block : T_1763_addr_block;
  assign T_1794_client_xact_id = T_1753 ? putAtomic_acquire_client_xact_id : T_1763_client_xact_id;
  assign T_1794_addr_beat = T_1753 ? putAtomic_acquire_addr_beat : T_1763_addr_beat;
  assign T_1794_is_builtin_type = T_1753 ? putAtomic_acquire_is_builtin_type : T_1763_is_builtin_type;
  assign T_1794_a_type = T_1753 ? putAtomic_acquire_a_type : T_1763_a_type;
  assign T_1794_union = T_1753 ? putAtomic_acquire_union : T_1763_union;
  assign T_1794_data = T_1753 ? putAtomic_acquire_data : T_1763_data;
  assign T_1825 = state == 3'h2;
  assign T_1827 = io_resp_ready == 1'h0;
  assign T_1828 = io_resp_valid & T_1827;
  assign T_1829 = T_1825 | T_1828;
  assign T_1830 = state == 3'h3;
  assign T_1841 = grant_word[63:32];
  assign T_1842 = grant_word[31:0];
  assign T_1843 = T_1310 ? T_1841 : T_1842;
  assign T_1851 = T_1843[31];
  assign T_1852 = T_1282 & T_1851;
  assign GEN_21 = {{31'd0}, T_1852};
  assign T_1854 = 32'h0 - GEN_21;
  assign T_1855 = T_1854[31:0];
  assign T_1857 = T_1338 ? T_1855 : T_1841;
  assign T_1858 = {T_1857,T_1843};
  assign T_1860 = T_1858[31:16];
  assign T_1861 = T_1858[15:0];
  assign T_1862 = T_1297 ? T_1860 : T_1861;
  assign T_1870 = T_1862[15];
  assign T_1871 = T_1282 & T_1870;
  assign GEN_23 = {{47'd0}, T_1871};
  assign T_1873 = 48'h0 - GEN_23;
  assign T_1874 = T_1873[47:0];
  assign T_1875 = T_1858[63:16];
  assign T_1876 = T_1333 ? T_1874 : T_1875;
  assign T_1877 = {T_1876,T_1862};
  assign T_1879 = T_1877[15:8];
  assign T_1880 = T_1877[7:0];
  assign T_1881 = T_1284 ? T_1879 : T_1880;
  assign T_1885 = req_cmd_sc ? {{7'd0}, 1'h0} : T_1881;
  assign T_1888 = T_1327 | req_cmd_sc;
  assign T_1889 = T_1885[7];
  assign T_1890 = T_1282 & T_1889;
  assign GEN_25 = {{55'd0}, T_1890};
  assign T_1892 = 56'h0 - GEN_25;
  assign T_1893 = T_1892[55:0];
  assign T_1894 = T_1877[63:8];
  assign T_1895 = T_1888 ? T_1893 : T_1894;
  assign T_1896 = {T_1895,T_1885};
  assign GEN_26 = {{63'd0}, req_cmd_sc};
  assign T_1897 = T_1896 | GEN_26;
  assign T_1899 = io_req_ready & io_req_valid;
  assign GEN_0 = T_1899 ? io_req_bits_addr : req_addr;
  assign GEN_1 = T_1899 ? io_req_bits_tag : req_tag;
  assign GEN_2 = T_1899 ? io_req_bits_cmd : req_cmd;
  assign GEN_3 = T_1899 ? io_req_bits_typ : req_typ;
  assign GEN_4 = T_1899 ? io_req_bits_phys : req_phys;
  assign GEN_5 = T_1899 ? io_req_bits_data : req_data;
  assign GEN_6 = T_1899 ? 3'h1 : state;
  assign T_1900 = io_acquire_ready & io_acquire_valid;
  assign GEN_7 = T_1900 ? 3'h2 : GEN_6;
  assign T_1902 = T_1825 & io_grant_valid;
  assign T_1915 = io_grant_bits_data >> 7'h0;
  assign GEN_8 = T_1762 ? T_1915 : grant_word;
  assign GEN_9 = T_1902 ? 3'h3 : GEN_7;
  assign GEN_10 = T_1902 ? GEN_8 : grant_word;
  assign T_1917 = io_resp_ready & io_resp_valid;
  assign GEN_11 = T_1917 ? 3'h4 : GEN_9;
  assign T_1918 = io_finish_ready & io_finish_valid;
  assign GEN_12 = T_1918 ? 3'h0 : GEN_11;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_22 = {2{$random}};
  req_addr = GEN_22[39:0];
  GEN_24 = {1{$random}};
  req_tag = GEN_24[8:0];
  GEN_27 = {1{$random}};
  req_cmd = GEN_27[4:0];
  GEN_28 = {1{$random}};
  req_typ = GEN_28[2:0];
  GEN_29 = {1{$random}};
  req_phys = GEN_29[0:0];
  GEN_30 = {2{$random}};
  req_data = GEN_30[63:0];
  GEN_31 = {2{$random}};
  grant_word = GEN_31[63:0];
  GEN_32 = {1{$random}};
  state = GEN_32[2:0];
  GEN_33 = {2{$random}};
  GEN_19 = GEN_33[63:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      req_addr <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      req_tag <= GEN_1;
    end
    if(1'h0) begin
    end else begin
      req_cmd <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      req_typ <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      req_phys <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      req_data <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      grant_word <= GEN_10;
    end
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_12;
    end
  end
endmodule
module MSHRFile(
  input   clk,
  input   reset,
  output  io_req_ready,
  input   io_req_valid,
  input  [39:0] io_req_bits_addr,
  input  [8:0] io_req_bits_tag,
  input  [4:0] io_req_bits_cmd,
  input  [2:0] io_req_bits_typ,
  input   io_req_bits_phys,
  input  [63:0] io_req_bits_data,
  input   io_req_bits_tag_match,
  input  [19:0] io_req_bits_old_meta_tag,
  input  [1:0] io_req_bits_old_meta_coh_state,
  input  [3:0] io_req_bits_way_en,
  input   io_resp_ready,
  output  io_resp_valid,
  output [39:0] io_resp_bits_addr,
  output [8:0] io_resp_bits_tag,
  output [4:0] io_resp_bits_cmd,
  output [2:0] io_resp_bits_typ,
  output [63:0] io_resp_bits_data,
  output  io_resp_bits_replay,
  output  io_resp_bits_has_data,
  output [63:0] io_resp_bits_data_word_bypass,
  output [63:0] io_resp_bits_store_data,
  output  io_secondary_miss,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [25:0] io_mem_req_bits_addr_block,
  output [1:0] io_mem_req_bits_client_xact_id,
  output [2:0] io_mem_req_bits_addr_beat,
  output  io_mem_req_bits_is_builtin_type,
  output [2:0] io_mem_req_bits_a_type,
  output [11:0] io_mem_req_bits_union,
  output [63:0] io_mem_req_bits_data,
  output [3:0] io_refill_way_en,
  output [11:0] io_refill_addr,
  input   io_meta_read_ready,
  output  io_meta_read_valid,
  output [5:0] io_meta_read_bits_idx,
  output [3:0] io_meta_read_bits_way_en,
  output [19:0] io_meta_read_bits_tag,
  input   io_meta_write_ready,
  output  io_meta_write_valid,
  output [5:0] io_meta_write_bits_idx,
  output [3:0] io_meta_write_bits_way_en,
  output [19:0] io_meta_write_bits_data_tag,
  output [1:0] io_meta_write_bits_data_coh_state,
  input   io_replay_ready,
  output  io_replay_valid,
  output [39:0] io_replay_bits_addr,
  output [8:0] io_replay_bits_tag,
  output [4:0] io_replay_bits_cmd,
  output [2:0] io_replay_bits_typ,
  output  io_replay_bits_phys,
  output [63:0] io_replay_bits_data,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id,
  input   io_wb_req_ready,
  output  io_wb_req_valid,
  output [2:0] io_wb_req_bits_addr_beat,
  output [25:0] io_wb_req_bits_addr_block,
  output [1:0] io_wb_req_bits_client_xact_id,
  output  io_wb_req_bits_voluntary,
  output [2:0] io_wb_req_bits_r_type,
  output [63:0] io_wb_req_bits_data,
  output [3:0] io_wb_req_bits_way_en,
  output  io_probe_rdy,
  output  io_fence_rdy,
  output  io_replay_next
);
  wire [39:0] GEN_17;
  wire  T_2615;
  wire [39:0] GEN_18;
  wire  T_2617;
  wire  T_2618;
  reg [16:0] sdq_val;
  reg [31:0] GEN_5;
  wire [16:0] T_2622;
  wire  T_2623;
  wire  T_2624;
  wire  T_2625;
  wire  T_2626;
  wire  T_2627;
  wire  T_2628;
  wire  T_2629;
  wire  T_2630;
  wire  T_2631;
  wire  T_2632;
  wire  T_2633;
  wire  T_2634;
  wire  T_2635;
  wire  T_2636;
  wire  T_2637;
  wire  T_2638;
  wire  T_2639;
  wire [4:0] T_2657;
  wire [4:0] T_2658;
  wire [4:0] T_2659;
  wire [4:0] T_2660;
  wire [4:0] T_2661;
  wire [4:0] T_2662;
  wire [4:0] T_2663;
  wire [4:0] T_2664;
  wire [4:0] T_2665;
  wire [4:0] T_2666;
  wire [4:0] T_2667;
  wire [4:0] T_2668;
  wire [4:0] T_2669;
  wire [4:0] T_2670;
  wire [4:0] T_2671;
  wire [4:0] sdq_alloc_id;
  wire [16:0] GEN_19;
  wire  T_2674;
  wire  sdq_rdy;
  wire  T_2676;
  wire  T_2677;
  wire  T_2678;
  wire  T_2679;
  wire  T_2680;
  wire  T_2681;
  wire  T_2682;
  wire  T_2683;
  wire  T_2684;
  wire  sdq_enq;
  reg [63:0] sdq [0:16];
  reg [63:0] GEN_6;
  wire [63:0] sdq_T_4084_data;
  wire [4:0] sdq_T_4084_addr;
  wire  sdq_T_4084_en;
  wire [63:0] sdq_T_2686_data;
  wire [4:0] sdq_T_2686_addr;
  wire  sdq_T_2686_mask;
  wire  sdq_T_2686_en;
  wire  idxMatch_0;
  wire  idxMatch_1;
  wire [19:0] tagList_0;
  wire [19:0] tagList_1;
  wire [19:0] T_2702;
  wire [19:0] T_2704;
  wire [19:0] T_2706;
  wire [19:0] T_2707;
  wire [27:0] T_2708;
  wire [27:0] GEN_20;
  wire  tag_match;
  wire [19:0] wbTagList_0;
  wire [19:0] wbTagList_1;
  wire [3:0] refillMux_0_way_en;
  wire [11:0] refillMux_0_addr;
  wire [3:0] refillMux_1_way_en;
  wire [11:0] refillMux_1_addr;
  wire  meta_read_arb_clk;
  wire  meta_read_arb_reset;
  wire  meta_read_arb_io_in_0_ready;
  wire  meta_read_arb_io_in_0_valid;
  wire [5:0] meta_read_arb_io_in_0_bits_idx;
  wire [3:0] meta_read_arb_io_in_0_bits_way_en;
  wire [19:0] meta_read_arb_io_in_0_bits_tag;
  wire  meta_read_arb_io_in_1_ready;
  wire  meta_read_arb_io_in_1_valid;
  wire [5:0] meta_read_arb_io_in_1_bits_idx;
  wire [3:0] meta_read_arb_io_in_1_bits_way_en;
  wire [19:0] meta_read_arb_io_in_1_bits_tag;
  wire  meta_read_arb_io_out_ready;
  wire  meta_read_arb_io_out_valid;
  wire [5:0] meta_read_arb_io_out_bits_idx;
  wire [3:0] meta_read_arb_io_out_bits_way_en;
  wire [19:0] meta_read_arb_io_out_bits_tag;
  wire  meta_read_arb_io_chosen;
  wire  meta_write_arb_clk;
  wire  meta_write_arb_reset;
  wire  meta_write_arb_io_in_0_ready;
  wire  meta_write_arb_io_in_0_valid;
  wire [5:0] meta_write_arb_io_in_0_bits_idx;
  wire [3:0] meta_write_arb_io_in_0_bits_way_en;
  wire [19:0] meta_write_arb_io_in_0_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_0_bits_data_coh_state;
  wire  meta_write_arb_io_in_1_ready;
  wire  meta_write_arb_io_in_1_valid;
  wire [5:0] meta_write_arb_io_in_1_bits_idx;
  wire [3:0] meta_write_arb_io_in_1_bits_way_en;
  wire [19:0] meta_write_arb_io_in_1_bits_data_tag;
  wire [1:0] meta_write_arb_io_in_1_bits_data_coh_state;
  wire  meta_write_arb_io_out_ready;
  wire  meta_write_arb_io_out_valid;
  wire [5:0] meta_write_arb_io_out_bits_idx;
  wire [3:0] meta_write_arb_io_out_bits_way_en;
  wire [19:0] meta_write_arb_io_out_bits_data_tag;
  wire [1:0] meta_write_arb_io_out_bits_data_coh_state;
  wire  meta_write_arb_io_chosen;
  wire  mem_req_arb_clk;
  wire  mem_req_arb_reset;
  wire  mem_req_arb_io_in_0_ready;
  wire  mem_req_arb_io_in_0_valid;
  wire [25:0] mem_req_arb_io_in_0_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_0_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_0_bits_addr_beat;
  wire  mem_req_arb_io_in_0_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_0_bits_a_type;
  wire [11:0] mem_req_arb_io_in_0_bits_union;
  wire [63:0] mem_req_arb_io_in_0_bits_data;
  wire  mem_req_arb_io_in_1_ready;
  wire  mem_req_arb_io_in_1_valid;
  wire [25:0] mem_req_arb_io_in_1_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_1_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_1_bits_addr_beat;
  wire  mem_req_arb_io_in_1_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_1_bits_a_type;
  wire [11:0] mem_req_arb_io_in_1_bits_union;
  wire [63:0] mem_req_arb_io_in_1_bits_data;
  wire  mem_req_arb_io_in_2_ready;
  wire  mem_req_arb_io_in_2_valid;
  wire [25:0] mem_req_arb_io_in_2_bits_addr_block;
  wire [1:0] mem_req_arb_io_in_2_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_in_2_bits_addr_beat;
  wire  mem_req_arb_io_in_2_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_in_2_bits_a_type;
  wire [11:0] mem_req_arb_io_in_2_bits_union;
  wire [63:0] mem_req_arb_io_in_2_bits_data;
  wire  mem_req_arb_io_out_ready;
  wire  mem_req_arb_io_out_valid;
  wire [25:0] mem_req_arb_io_out_bits_addr_block;
  wire [1:0] mem_req_arb_io_out_bits_client_xact_id;
  wire [2:0] mem_req_arb_io_out_bits_addr_beat;
  wire  mem_req_arb_io_out_bits_is_builtin_type;
  wire [2:0] mem_req_arb_io_out_bits_a_type;
  wire [11:0] mem_req_arb_io_out_bits_union;
  wire [63:0] mem_req_arb_io_out_bits_data;
  wire [1:0] mem_req_arb_io_chosen;
  wire  mem_finish_arb_clk;
  wire  mem_finish_arb_reset;
  wire  mem_finish_arb_io_in_0_ready;
  wire  mem_finish_arb_io_in_0_valid;
  wire [2:0] mem_finish_arb_io_in_0_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_0_bits_manager_id;
  wire  mem_finish_arb_io_in_1_ready;
  wire  mem_finish_arb_io_in_1_valid;
  wire [2:0] mem_finish_arb_io_in_1_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_1_bits_manager_id;
  wire  mem_finish_arb_io_in_2_ready;
  wire  mem_finish_arb_io_in_2_valid;
  wire [2:0] mem_finish_arb_io_in_2_bits_manager_xact_id;
  wire  mem_finish_arb_io_in_2_bits_manager_id;
  wire  mem_finish_arb_io_out_ready;
  wire  mem_finish_arb_io_out_valid;
  wire [2:0] mem_finish_arb_io_out_bits_manager_xact_id;
  wire  mem_finish_arb_io_out_bits_manager_id;
  wire [1:0] mem_finish_arb_io_chosen;
  wire  wb_req_arb_clk;
  wire  wb_req_arb_reset;
  wire  wb_req_arb_io_in_0_ready;
  wire  wb_req_arb_io_in_0_valid;
  wire [2:0] wb_req_arb_io_in_0_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_0_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_0_bits_client_xact_id;
  wire  wb_req_arb_io_in_0_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_0_bits_r_type;
  wire [63:0] wb_req_arb_io_in_0_bits_data;
  wire [3:0] wb_req_arb_io_in_0_bits_way_en;
  wire  wb_req_arb_io_in_1_ready;
  wire  wb_req_arb_io_in_1_valid;
  wire [2:0] wb_req_arb_io_in_1_bits_addr_beat;
  wire [25:0] wb_req_arb_io_in_1_bits_addr_block;
  wire [1:0] wb_req_arb_io_in_1_bits_client_xact_id;
  wire  wb_req_arb_io_in_1_bits_voluntary;
  wire [2:0] wb_req_arb_io_in_1_bits_r_type;
  wire [63:0] wb_req_arb_io_in_1_bits_data;
  wire [3:0] wb_req_arb_io_in_1_bits_way_en;
  wire  wb_req_arb_io_out_ready;
  wire  wb_req_arb_io_out_valid;
  wire [2:0] wb_req_arb_io_out_bits_addr_beat;
  wire [25:0] wb_req_arb_io_out_bits_addr_block;
  wire [1:0] wb_req_arb_io_out_bits_client_xact_id;
  wire  wb_req_arb_io_out_bits_voluntary;
  wire [2:0] wb_req_arb_io_out_bits_r_type;
  wire [63:0] wb_req_arb_io_out_bits_data;
  wire [3:0] wb_req_arb_io_out_bits_way_en;
  wire  wb_req_arb_io_chosen;
  wire  replay_arb_clk;
  wire  replay_arb_reset;
  wire  replay_arb_io_in_0_ready;
  wire  replay_arb_io_in_0_valid;
  wire [39:0] replay_arb_io_in_0_bits_addr;
  wire [8:0] replay_arb_io_in_0_bits_tag;
  wire [4:0] replay_arb_io_in_0_bits_cmd;
  wire [2:0] replay_arb_io_in_0_bits_typ;
  wire  replay_arb_io_in_0_bits_phys;
  wire [4:0] replay_arb_io_in_0_bits_sdq_id;
  wire  replay_arb_io_in_1_ready;
  wire  replay_arb_io_in_1_valid;
  wire [39:0] replay_arb_io_in_1_bits_addr;
  wire [8:0] replay_arb_io_in_1_bits_tag;
  wire [4:0] replay_arb_io_in_1_bits_cmd;
  wire [2:0] replay_arb_io_in_1_bits_typ;
  wire  replay_arb_io_in_1_bits_phys;
  wire [4:0] replay_arb_io_in_1_bits_sdq_id;
  wire  replay_arb_io_out_ready;
  wire  replay_arb_io_out_valid;
  wire [39:0] replay_arb_io_out_bits_addr;
  wire [8:0] replay_arb_io_out_bits_tag;
  wire [4:0] replay_arb_io_out_bits_cmd;
  wire [2:0] replay_arb_io_out_bits_typ;
  wire  replay_arb_io_out_bits_phys;
  wire [4:0] replay_arb_io_out_bits_sdq_id;
  wire  replay_arb_io_chosen;
  wire  alloc_arb_clk;
  wire  alloc_arb_reset;
  wire  alloc_arb_io_in_0_ready;
  wire  alloc_arb_io_in_0_valid;
  wire  alloc_arb_io_in_0_bits;
  wire  alloc_arb_io_in_1_ready;
  wire  alloc_arb_io_in_1_valid;
  wire  alloc_arb_io_in_1_bits;
  wire  alloc_arb_io_out_ready;
  wire  alloc_arb_io_out_valid;
  wire  alloc_arb_io_out_bits;
  wire  alloc_arb_io_chosen;
  wire  MSHR_3871_clk;
  wire  MSHR_3871_reset;
  wire  MSHR_3871_io_req_pri_val;
  wire  MSHR_3871_io_req_pri_rdy;
  wire  MSHR_3871_io_req_sec_val;
  wire  MSHR_3871_io_req_sec_rdy;
  wire [39:0] MSHR_3871_io_req_bits_addr;
  wire [8:0] MSHR_3871_io_req_bits_tag;
  wire [4:0] MSHR_3871_io_req_bits_cmd;
  wire [2:0] MSHR_3871_io_req_bits_typ;
  wire  MSHR_3871_io_req_bits_phys;
  wire [4:0] MSHR_3871_io_req_bits_sdq_id;
  wire  MSHR_3871_io_req_bits_tag_match;
  wire [19:0] MSHR_3871_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_3871_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_3871_io_req_bits_way_en;
  wire  MSHR_3871_io_idx_match;
  wire [19:0] MSHR_3871_io_tag;
  wire  MSHR_3871_io_mem_req_ready;
  wire  MSHR_3871_io_mem_req_valid;
  wire [25:0] MSHR_3871_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_3871_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_3871_io_mem_req_bits_addr_beat;
  wire  MSHR_3871_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_3871_io_mem_req_bits_a_type;
  wire [11:0] MSHR_3871_io_mem_req_bits_union;
  wire [63:0] MSHR_3871_io_mem_req_bits_data;
  wire [3:0] MSHR_3871_io_refill_way_en;
  wire [11:0] MSHR_3871_io_refill_addr;
  wire  MSHR_3871_io_meta_read_ready;
  wire  MSHR_3871_io_meta_read_valid;
  wire [5:0] MSHR_3871_io_meta_read_bits_idx;
  wire [3:0] MSHR_3871_io_meta_read_bits_way_en;
  wire [19:0] MSHR_3871_io_meta_read_bits_tag;
  wire  MSHR_3871_io_meta_write_ready;
  wire  MSHR_3871_io_meta_write_valid;
  wire [5:0] MSHR_3871_io_meta_write_bits_idx;
  wire [3:0] MSHR_3871_io_meta_write_bits_way_en;
  wire [19:0] MSHR_3871_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_3871_io_meta_write_bits_data_coh_state;
  wire  MSHR_3871_io_replay_ready;
  wire  MSHR_3871_io_replay_valid;
  wire [39:0] MSHR_3871_io_replay_bits_addr;
  wire [8:0] MSHR_3871_io_replay_bits_tag;
  wire [4:0] MSHR_3871_io_replay_bits_cmd;
  wire [2:0] MSHR_3871_io_replay_bits_typ;
  wire  MSHR_3871_io_replay_bits_phys;
  wire [4:0] MSHR_3871_io_replay_bits_sdq_id;
  wire  MSHR_3871_io_mem_grant_valid;
  wire [2:0] MSHR_3871_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_3871_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_3871_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_3871_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_3871_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_3871_io_mem_grant_bits_data;
  wire  MSHR_3871_io_mem_grant_bits_manager_id;
  wire  MSHR_3871_io_mem_finish_ready;
  wire  MSHR_3871_io_mem_finish_valid;
  wire [2:0] MSHR_3871_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_3871_io_mem_finish_bits_manager_id;
  wire  MSHR_3871_io_wb_req_ready;
  wire  MSHR_3871_io_wb_req_valid;
  wire [2:0] MSHR_3871_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_3871_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_3871_io_wb_req_bits_client_xact_id;
  wire  MSHR_3871_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_3871_io_wb_req_bits_r_type;
  wire [63:0] MSHR_3871_io_wb_req_bits_data;
  wire [3:0] MSHR_3871_io_wb_req_bits_way_en;
  wire  MSHR_3871_io_probe_rdy;
  wire [19:0] T_3872;
  wire  T_3873;
  wire  T_3874;
  wire [1:0] GEN_21;
  wire  T_3876;
  wire  T_3877;
  wire  T_3878;
  wire  T_3879;
  wire  T_3880;
  wire  T_3882;
  wire  GEN_7;
  wire  T_3885;
  wire  GEN_8;
  wire  MSHR_75_3887_clk;
  wire  MSHR_75_3887_reset;
  wire  MSHR_75_3887_io_req_pri_val;
  wire  MSHR_75_3887_io_req_pri_rdy;
  wire  MSHR_75_3887_io_req_sec_val;
  wire  MSHR_75_3887_io_req_sec_rdy;
  wire [39:0] MSHR_75_3887_io_req_bits_addr;
  wire [8:0] MSHR_75_3887_io_req_bits_tag;
  wire [4:0] MSHR_75_3887_io_req_bits_cmd;
  wire [2:0] MSHR_75_3887_io_req_bits_typ;
  wire  MSHR_75_3887_io_req_bits_phys;
  wire [4:0] MSHR_75_3887_io_req_bits_sdq_id;
  wire  MSHR_75_3887_io_req_bits_tag_match;
  wire [19:0] MSHR_75_3887_io_req_bits_old_meta_tag;
  wire [1:0] MSHR_75_3887_io_req_bits_old_meta_coh_state;
  wire [3:0] MSHR_75_3887_io_req_bits_way_en;
  wire  MSHR_75_3887_io_idx_match;
  wire [19:0] MSHR_75_3887_io_tag;
  wire  MSHR_75_3887_io_mem_req_ready;
  wire  MSHR_75_3887_io_mem_req_valid;
  wire [25:0] MSHR_75_3887_io_mem_req_bits_addr_block;
  wire [1:0] MSHR_75_3887_io_mem_req_bits_client_xact_id;
  wire [2:0] MSHR_75_3887_io_mem_req_bits_addr_beat;
  wire  MSHR_75_3887_io_mem_req_bits_is_builtin_type;
  wire [2:0] MSHR_75_3887_io_mem_req_bits_a_type;
  wire [11:0] MSHR_75_3887_io_mem_req_bits_union;
  wire [63:0] MSHR_75_3887_io_mem_req_bits_data;
  wire [3:0] MSHR_75_3887_io_refill_way_en;
  wire [11:0] MSHR_75_3887_io_refill_addr;
  wire  MSHR_75_3887_io_meta_read_ready;
  wire  MSHR_75_3887_io_meta_read_valid;
  wire [5:0] MSHR_75_3887_io_meta_read_bits_idx;
  wire [3:0] MSHR_75_3887_io_meta_read_bits_way_en;
  wire [19:0] MSHR_75_3887_io_meta_read_bits_tag;
  wire  MSHR_75_3887_io_meta_write_ready;
  wire  MSHR_75_3887_io_meta_write_valid;
  wire [5:0] MSHR_75_3887_io_meta_write_bits_idx;
  wire [3:0] MSHR_75_3887_io_meta_write_bits_way_en;
  wire [19:0] MSHR_75_3887_io_meta_write_bits_data_tag;
  wire [1:0] MSHR_75_3887_io_meta_write_bits_data_coh_state;
  wire  MSHR_75_3887_io_replay_ready;
  wire  MSHR_75_3887_io_replay_valid;
  wire [39:0] MSHR_75_3887_io_replay_bits_addr;
  wire [8:0] MSHR_75_3887_io_replay_bits_tag;
  wire [4:0] MSHR_75_3887_io_replay_bits_cmd;
  wire [2:0] MSHR_75_3887_io_replay_bits_typ;
  wire  MSHR_75_3887_io_replay_bits_phys;
  wire [4:0] MSHR_75_3887_io_replay_bits_sdq_id;
  wire  MSHR_75_3887_io_mem_grant_valid;
  wire [2:0] MSHR_75_3887_io_mem_grant_bits_addr_beat;
  wire [1:0] MSHR_75_3887_io_mem_grant_bits_client_xact_id;
  wire [2:0] MSHR_75_3887_io_mem_grant_bits_manager_xact_id;
  wire  MSHR_75_3887_io_mem_grant_bits_is_builtin_type;
  wire [3:0] MSHR_75_3887_io_mem_grant_bits_g_type;
  wire [63:0] MSHR_75_3887_io_mem_grant_bits_data;
  wire  MSHR_75_3887_io_mem_grant_bits_manager_id;
  wire  MSHR_75_3887_io_mem_finish_ready;
  wire  MSHR_75_3887_io_mem_finish_valid;
  wire [2:0] MSHR_75_3887_io_mem_finish_bits_manager_xact_id;
  wire  MSHR_75_3887_io_mem_finish_bits_manager_id;
  wire  MSHR_75_3887_io_wb_req_ready;
  wire  MSHR_75_3887_io_wb_req_valid;
  wire [2:0] MSHR_75_3887_io_wb_req_bits_addr_beat;
  wire [25:0] MSHR_75_3887_io_wb_req_bits_addr_block;
  wire [1:0] MSHR_75_3887_io_wb_req_bits_client_xact_id;
  wire  MSHR_75_3887_io_wb_req_bits_voluntary;
  wire [2:0] MSHR_75_3887_io_wb_req_bits_r_type;
  wire [63:0] MSHR_75_3887_io_wb_req_bits_data;
  wire [3:0] MSHR_75_3887_io_wb_req_bits_way_en;
  wire  MSHR_75_3887_io_probe_rdy;
  wire [19:0] T_3888;
  wire [1:0] GEN_22;
  wire  T_3892;
  wire  T_3893;
  wire  pri_rdy;
  wire  sec_rdy;
  wire  idx_match;
  wire  T_3895;
  wire  GEN_9;
  wire  T_3898;
  wire  GEN_10;
  wire  T_3901;
  wire  T_3903;
  wire  T_3904;
  wire  mmio_alloc_arb_clk;
  wire  mmio_alloc_arb_reset;
  wire  mmio_alloc_arb_io_in_0_ready;
  wire  mmio_alloc_arb_io_in_0_valid;
  wire  mmio_alloc_arb_io_in_0_bits;
  wire  mmio_alloc_arb_io_out_ready;
  wire  mmio_alloc_arb_io_out_valid;
  wire  mmio_alloc_arb_io_out_bits;
  wire  mmio_alloc_arb_io_chosen;
  wire  resp_arb_clk;
  wire  resp_arb_reset;
  wire  resp_arb_io_in_0_ready;
  wire  resp_arb_io_in_0_valid;
  wire [39:0] resp_arb_io_in_0_bits_addr;
  wire [8:0] resp_arb_io_in_0_bits_tag;
  wire [4:0] resp_arb_io_in_0_bits_cmd;
  wire [2:0] resp_arb_io_in_0_bits_typ;
  wire [63:0] resp_arb_io_in_0_bits_data;
  wire  resp_arb_io_in_0_bits_replay;
  wire  resp_arb_io_in_0_bits_has_data;
  wire [63:0] resp_arb_io_in_0_bits_data_word_bypass;
  wire [63:0] resp_arb_io_in_0_bits_store_data;
  wire  resp_arb_io_out_ready;
  wire  resp_arb_io_out_valid;
  wire [39:0] resp_arb_io_out_bits_addr;
  wire [8:0] resp_arb_io_out_bits_tag;
  wire [4:0] resp_arb_io_out_bits_cmd;
  wire [2:0] resp_arb_io_out_bits_typ;
  wire [63:0] resp_arb_io_out_bits_data;
  wire  resp_arb_io_out_bits_replay;
  wire  resp_arb_io_out_bits_has_data;
  wire [63:0] resp_arb_io_out_bits_data_word_bypass;
  wire [63:0] resp_arb_io_out_bits_store_data;
  wire  resp_arb_io_chosen;
  wire  IOMSHR_3987_clk;
  wire  IOMSHR_3987_reset;
  wire  IOMSHR_3987_io_req_ready;
  wire  IOMSHR_3987_io_req_valid;
  wire [39:0] IOMSHR_3987_io_req_bits_addr;
  wire [8:0] IOMSHR_3987_io_req_bits_tag;
  wire [4:0] IOMSHR_3987_io_req_bits_cmd;
  wire [2:0] IOMSHR_3987_io_req_bits_typ;
  wire  IOMSHR_3987_io_req_bits_phys;
  wire [63:0] IOMSHR_3987_io_req_bits_data;
  wire  IOMSHR_3987_io_acquire_ready;
  wire  IOMSHR_3987_io_acquire_valid;
  wire [25:0] IOMSHR_3987_io_acquire_bits_addr_block;
  wire [1:0] IOMSHR_3987_io_acquire_bits_client_xact_id;
  wire [2:0] IOMSHR_3987_io_acquire_bits_addr_beat;
  wire  IOMSHR_3987_io_acquire_bits_is_builtin_type;
  wire [2:0] IOMSHR_3987_io_acquire_bits_a_type;
  wire [11:0] IOMSHR_3987_io_acquire_bits_union;
  wire [63:0] IOMSHR_3987_io_acquire_bits_data;
  wire  IOMSHR_3987_io_grant_valid;
  wire [2:0] IOMSHR_3987_io_grant_bits_addr_beat;
  wire [1:0] IOMSHR_3987_io_grant_bits_client_xact_id;
  wire [2:0] IOMSHR_3987_io_grant_bits_manager_xact_id;
  wire  IOMSHR_3987_io_grant_bits_is_builtin_type;
  wire [3:0] IOMSHR_3987_io_grant_bits_g_type;
  wire [63:0] IOMSHR_3987_io_grant_bits_data;
  wire  IOMSHR_3987_io_grant_bits_manager_id;
  wire  IOMSHR_3987_io_finish_ready;
  wire  IOMSHR_3987_io_finish_valid;
  wire [2:0] IOMSHR_3987_io_finish_bits_manager_xact_id;
  wire  IOMSHR_3987_io_finish_bits_manager_id;
  wire  IOMSHR_3987_io_resp_ready;
  wire  IOMSHR_3987_io_resp_valid;
  wire [39:0] IOMSHR_3987_io_resp_bits_addr;
  wire [8:0] IOMSHR_3987_io_resp_bits_tag;
  wire [4:0] IOMSHR_3987_io_resp_bits_cmd;
  wire [2:0] IOMSHR_3987_io_resp_bits_typ;
  wire [63:0] IOMSHR_3987_io_resp_bits_data;
  wire  IOMSHR_3987_io_resp_bits_replay;
  wire  IOMSHR_3987_io_resp_bits_has_data;
  wire [63:0] IOMSHR_3987_io_resp_bits_data_word_bypass;
  wire [63:0] IOMSHR_3987_io_resp_bits_store_data;
  wire  IOMSHR_3987_io_replay_next;
  wire  mmio_rdy;
  wire  T_3989;
  wire  T_3990;
  wire  T_3992;
  wire  GEN_11;
  wire  GEN_12;
  wire  T_3996;
  wire  T_3997;
  wire  T_4000;
  wire  T_4001;
  wire  T_4002;
  wire  T_4003;
  wire [3:0] GEN_0;
  wire [3:0] GEN_13;
  wire [11:0] GEN_1;
  wire [11:0] GEN_14;
  wire  T_4075;
  wire  T_4076;
  wire  T_4077;
  wire  T_4078;
  wire  T_4079;
  wire  T_4080;
  wire  T_4081;
  wire  T_4082;
  wire  free_sdq;
  reg [4:0] T_4083;
  reg [31:0] GEN_23;
  wire [4:0] GEN_15;
  wire  T_4085;
  wire [31:0] GEN_25;
  wire [31:0] T_4087;
  wire [16:0] GEN_26;
  wire [17:0] T_4089;
  wire [16:0] T_4090;
  wire [31:0] GEN_27;
  wire [31:0] T_4091;
  wire [31:0] T_4092;
  wire [31:0] GEN_28;
  wire [31:0] T_4093;
  wire [16:0] T_4132;
  wire [16:0] T_4133;
  wire [16:0] T_4134;
  wire [16:0] T_4135;
  wire [16:0] T_4136;
  wire [16:0] T_4137;
  wire [16:0] T_4138;
  wire [16:0] T_4139;
  wire [16:0] T_4140;
  wire [16:0] T_4141;
  wire [16:0] T_4142;
  wire [16:0] T_4143;
  wire [16:0] T_4144;
  wire [16:0] T_4145;
  wire [16:0] T_4146;
  wire [16:0] T_4147;
  wire [16:0] T_4148;
  wire [16:0] GEN_29;
  wire [17:0] T_4150;
  wire [16:0] T_4151;
  wire [16:0] T_4152;
  wire [31:0] GEN_30;
  wire [31:0] T_4153;
  wire [31:0] GEN_16;
  reg  GEN_2;
  reg [31:0] GEN_24;
  reg  GEN_3;
  reg [31:0] GEN_31;
  reg  GEN_4;
  reg [31:0] GEN_32;
  Arbiter_67 meta_read_arb (
    .clk(meta_read_arb_clk),
    .reset(meta_read_arb_reset),
    .io_in_0_ready(meta_read_arb_io_in_0_ready),
    .io_in_0_valid(meta_read_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_read_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_read_arb_io_in_0_bits_way_en),
    .io_in_0_bits_tag(meta_read_arb_io_in_0_bits_tag),
    .io_in_1_ready(meta_read_arb_io_in_1_ready),
    .io_in_1_valid(meta_read_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_read_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_read_arb_io_in_1_bits_way_en),
    .io_in_1_bits_tag(meta_read_arb_io_in_1_bits_tag),
    .io_out_ready(meta_read_arb_io_out_ready),
    .io_out_valid(meta_read_arb_io_out_valid),
    .io_out_bits_idx(meta_read_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_read_arb_io_out_bits_way_en),
    .io_out_bits_tag(meta_read_arb_io_out_bits_tag),
    .io_chosen(meta_read_arb_io_chosen)
  );
  Arbiter_68 meta_write_arb (
    .clk(meta_write_arb_clk),
    .reset(meta_write_arb_reset),
    .io_in_0_ready(meta_write_arb_io_in_0_ready),
    .io_in_0_valid(meta_write_arb_io_in_0_valid),
    .io_in_0_bits_idx(meta_write_arb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(meta_write_arb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(meta_write_arb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(meta_write_arb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(meta_write_arb_io_in_1_ready),
    .io_in_1_valid(meta_write_arb_io_in_1_valid),
    .io_in_1_bits_idx(meta_write_arb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(meta_write_arb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(meta_write_arb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(meta_write_arb_io_in_1_bits_data_coh_state),
    .io_out_ready(meta_write_arb_io_out_ready),
    .io_out_valid(meta_write_arb_io_out_valid),
    .io_out_bits_idx(meta_write_arb_io_out_bits_idx),
    .io_out_bits_way_en(meta_write_arb_io_out_bits_way_en),
    .io_out_bits_data_tag(meta_write_arb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(meta_write_arb_io_out_bits_data_coh_state),
    .io_chosen(meta_write_arb_io_chosen)
  );
  LockingArbiter mem_req_arb (
    .clk(mem_req_arb_clk),
    .reset(mem_req_arb_reset),
    .io_in_0_ready(mem_req_arb_io_in_0_ready),
    .io_in_0_valid(mem_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_block(mem_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(mem_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_addr_beat(mem_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_is_builtin_type(mem_req_arb_io_in_0_bits_is_builtin_type),
    .io_in_0_bits_a_type(mem_req_arb_io_in_0_bits_a_type),
    .io_in_0_bits_union(mem_req_arb_io_in_0_bits_union),
    .io_in_0_bits_data(mem_req_arb_io_in_0_bits_data),
    .io_in_1_ready(mem_req_arb_io_in_1_ready),
    .io_in_1_valid(mem_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_block(mem_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(mem_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_addr_beat(mem_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_is_builtin_type(mem_req_arb_io_in_1_bits_is_builtin_type),
    .io_in_1_bits_a_type(mem_req_arb_io_in_1_bits_a_type),
    .io_in_1_bits_union(mem_req_arb_io_in_1_bits_union),
    .io_in_1_bits_data(mem_req_arb_io_in_1_bits_data),
    .io_in_2_ready(mem_req_arb_io_in_2_ready),
    .io_in_2_valid(mem_req_arb_io_in_2_valid),
    .io_in_2_bits_addr_block(mem_req_arb_io_in_2_bits_addr_block),
    .io_in_2_bits_client_xact_id(mem_req_arb_io_in_2_bits_client_xact_id),
    .io_in_2_bits_addr_beat(mem_req_arb_io_in_2_bits_addr_beat),
    .io_in_2_bits_is_builtin_type(mem_req_arb_io_in_2_bits_is_builtin_type),
    .io_in_2_bits_a_type(mem_req_arb_io_in_2_bits_a_type),
    .io_in_2_bits_union(mem_req_arb_io_in_2_bits_union),
    .io_in_2_bits_data(mem_req_arb_io_in_2_bits_data),
    .io_out_ready(mem_req_arb_io_out_ready),
    .io_out_valid(mem_req_arb_io_out_valid),
    .io_out_bits_addr_block(mem_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(mem_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_addr_beat(mem_req_arb_io_out_bits_addr_beat),
    .io_out_bits_is_builtin_type(mem_req_arb_io_out_bits_is_builtin_type),
    .io_out_bits_a_type(mem_req_arb_io_out_bits_a_type),
    .io_out_bits_union(mem_req_arb_io_out_bits_union),
    .io_out_bits_data(mem_req_arb_io_out_bits_data),
    .io_chosen(mem_req_arb_io_chosen)
  );
  Arbiter_69 mem_finish_arb (
    .clk(mem_finish_arb_clk),
    .reset(mem_finish_arb_reset),
    .io_in_0_ready(mem_finish_arb_io_in_0_ready),
    .io_in_0_valid(mem_finish_arb_io_in_0_valid),
    .io_in_0_bits_manager_xact_id(mem_finish_arb_io_in_0_bits_manager_xact_id),
    .io_in_0_bits_manager_id(mem_finish_arb_io_in_0_bits_manager_id),
    .io_in_1_ready(mem_finish_arb_io_in_1_ready),
    .io_in_1_valid(mem_finish_arb_io_in_1_valid),
    .io_in_1_bits_manager_xact_id(mem_finish_arb_io_in_1_bits_manager_xact_id),
    .io_in_1_bits_manager_id(mem_finish_arb_io_in_1_bits_manager_id),
    .io_in_2_ready(mem_finish_arb_io_in_2_ready),
    .io_in_2_valid(mem_finish_arb_io_in_2_valid),
    .io_in_2_bits_manager_xact_id(mem_finish_arb_io_in_2_bits_manager_xact_id),
    .io_in_2_bits_manager_id(mem_finish_arb_io_in_2_bits_manager_id),
    .io_out_ready(mem_finish_arb_io_out_ready),
    .io_out_valid(mem_finish_arb_io_out_valid),
    .io_out_bits_manager_xact_id(mem_finish_arb_io_out_bits_manager_xact_id),
    .io_out_bits_manager_id(mem_finish_arb_io_out_bits_manager_id),
    .io_chosen(mem_finish_arb_io_chosen)
  );
  Arbiter_70 wb_req_arb (
    .clk(wb_req_arb_clk),
    .reset(wb_req_arb_reset),
    .io_in_0_ready(wb_req_arb_io_in_0_ready),
    .io_in_0_valid(wb_req_arb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wb_req_arb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wb_req_arb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wb_req_arb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wb_req_arb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wb_req_arb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wb_req_arb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wb_req_arb_io_in_0_bits_way_en),
    .io_in_1_ready(wb_req_arb_io_in_1_ready),
    .io_in_1_valid(wb_req_arb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wb_req_arb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wb_req_arb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wb_req_arb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wb_req_arb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wb_req_arb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wb_req_arb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wb_req_arb_io_in_1_bits_way_en),
    .io_out_ready(wb_req_arb_io_out_ready),
    .io_out_valid(wb_req_arb_io_out_valid),
    .io_out_bits_addr_beat(wb_req_arb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wb_req_arb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wb_req_arb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wb_req_arb_io_out_bits_voluntary),
    .io_out_bits_r_type(wb_req_arb_io_out_bits_r_type),
    .io_out_bits_data(wb_req_arb_io_out_bits_data),
    .io_out_bits_way_en(wb_req_arb_io_out_bits_way_en),
    .io_chosen(wb_req_arb_io_chosen)
  );
  Arbiter_71 replay_arb (
    .clk(replay_arb_clk),
    .reset(replay_arb_reset),
    .io_in_0_ready(replay_arb_io_in_0_ready),
    .io_in_0_valid(replay_arb_io_in_0_valid),
    .io_in_0_bits_addr(replay_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(replay_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(replay_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(replay_arb_io_in_0_bits_typ),
    .io_in_0_bits_phys(replay_arb_io_in_0_bits_phys),
    .io_in_0_bits_sdq_id(replay_arb_io_in_0_bits_sdq_id),
    .io_in_1_ready(replay_arb_io_in_1_ready),
    .io_in_1_valid(replay_arb_io_in_1_valid),
    .io_in_1_bits_addr(replay_arb_io_in_1_bits_addr),
    .io_in_1_bits_tag(replay_arb_io_in_1_bits_tag),
    .io_in_1_bits_cmd(replay_arb_io_in_1_bits_cmd),
    .io_in_1_bits_typ(replay_arb_io_in_1_bits_typ),
    .io_in_1_bits_phys(replay_arb_io_in_1_bits_phys),
    .io_in_1_bits_sdq_id(replay_arb_io_in_1_bits_sdq_id),
    .io_out_ready(replay_arb_io_out_ready),
    .io_out_valid(replay_arb_io_out_valid),
    .io_out_bits_addr(replay_arb_io_out_bits_addr),
    .io_out_bits_tag(replay_arb_io_out_bits_tag),
    .io_out_bits_cmd(replay_arb_io_out_bits_cmd),
    .io_out_bits_typ(replay_arb_io_out_bits_typ),
    .io_out_bits_phys(replay_arb_io_out_bits_phys),
    .io_out_bits_sdq_id(replay_arb_io_out_bits_sdq_id),
    .io_chosen(replay_arb_io_chosen)
  );
  Arbiter_72 alloc_arb (
    .clk(alloc_arb_clk),
    .reset(alloc_arb_reset),
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_0_bits(alloc_arb_io_in_0_bits),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_in_1_bits(alloc_arb_io_in_1_bits),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid),
    .io_out_bits(alloc_arb_io_out_bits),
    .io_chosen(alloc_arb_io_chosen)
  );
  MSHR MSHR_3871 (
    .clk(MSHR_3871_clk),
    .reset(MSHR_3871_reset),
    .io_req_pri_val(MSHR_3871_io_req_pri_val),
    .io_req_pri_rdy(MSHR_3871_io_req_pri_rdy),
    .io_req_sec_val(MSHR_3871_io_req_sec_val),
    .io_req_sec_rdy(MSHR_3871_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_3871_io_req_bits_addr),
    .io_req_bits_tag(MSHR_3871_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_3871_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_3871_io_req_bits_typ),
    .io_req_bits_phys(MSHR_3871_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_3871_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_3871_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_3871_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_3871_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_3871_io_req_bits_way_en),
    .io_idx_match(MSHR_3871_io_idx_match),
    .io_tag(MSHR_3871_io_tag),
    .io_mem_req_ready(MSHR_3871_io_mem_req_ready),
    .io_mem_req_valid(MSHR_3871_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_3871_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_3871_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_3871_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_3871_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_3871_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_3871_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_3871_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_3871_io_refill_way_en),
    .io_refill_addr(MSHR_3871_io_refill_addr),
    .io_meta_read_ready(MSHR_3871_io_meta_read_ready),
    .io_meta_read_valid(MSHR_3871_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_3871_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_3871_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_3871_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_3871_io_meta_write_ready),
    .io_meta_write_valid(MSHR_3871_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_3871_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_3871_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_3871_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_3871_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_3871_io_replay_ready),
    .io_replay_valid(MSHR_3871_io_replay_valid),
    .io_replay_bits_addr(MSHR_3871_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_3871_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_3871_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_3871_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_3871_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_3871_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_3871_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_3871_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_3871_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_3871_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_3871_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_3871_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_3871_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_3871_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_3871_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_3871_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_3871_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_3871_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_3871_io_wb_req_ready),
    .io_wb_req_valid(MSHR_3871_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_3871_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_3871_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_3871_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_3871_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_3871_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_3871_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_3871_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_3871_io_probe_rdy)
  );
  MSHR_75 MSHR_75_3887 (
    .clk(MSHR_75_3887_clk),
    .reset(MSHR_75_3887_reset),
    .io_req_pri_val(MSHR_75_3887_io_req_pri_val),
    .io_req_pri_rdy(MSHR_75_3887_io_req_pri_rdy),
    .io_req_sec_val(MSHR_75_3887_io_req_sec_val),
    .io_req_sec_rdy(MSHR_75_3887_io_req_sec_rdy),
    .io_req_bits_addr(MSHR_75_3887_io_req_bits_addr),
    .io_req_bits_tag(MSHR_75_3887_io_req_bits_tag),
    .io_req_bits_cmd(MSHR_75_3887_io_req_bits_cmd),
    .io_req_bits_typ(MSHR_75_3887_io_req_bits_typ),
    .io_req_bits_phys(MSHR_75_3887_io_req_bits_phys),
    .io_req_bits_sdq_id(MSHR_75_3887_io_req_bits_sdq_id),
    .io_req_bits_tag_match(MSHR_75_3887_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(MSHR_75_3887_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(MSHR_75_3887_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(MSHR_75_3887_io_req_bits_way_en),
    .io_idx_match(MSHR_75_3887_io_idx_match),
    .io_tag(MSHR_75_3887_io_tag),
    .io_mem_req_ready(MSHR_75_3887_io_mem_req_ready),
    .io_mem_req_valid(MSHR_75_3887_io_mem_req_valid),
    .io_mem_req_bits_addr_block(MSHR_75_3887_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(MSHR_75_3887_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(MSHR_75_3887_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(MSHR_75_3887_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(MSHR_75_3887_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(MSHR_75_3887_io_mem_req_bits_union),
    .io_mem_req_bits_data(MSHR_75_3887_io_mem_req_bits_data),
    .io_refill_way_en(MSHR_75_3887_io_refill_way_en),
    .io_refill_addr(MSHR_75_3887_io_refill_addr),
    .io_meta_read_ready(MSHR_75_3887_io_meta_read_ready),
    .io_meta_read_valid(MSHR_75_3887_io_meta_read_valid),
    .io_meta_read_bits_idx(MSHR_75_3887_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(MSHR_75_3887_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(MSHR_75_3887_io_meta_read_bits_tag),
    .io_meta_write_ready(MSHR_75_3887_io_meta_write_ready),
    .io_meta_write_valid(MSHR_75_3887_io_meta_write_valid),
    .io_meta_write_bits_idx(MSHR_75_3887_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(MSHR_75_3887_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(MSHR_75_3887_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(MSHR_75_3887_io_meta_write_bits_data_coh_state),
    .io_replay_ready(MSHR_75_3887_io_replay_ready),
    .io_replay_valid(MSHR_75_3887_io_replay_valid),
    .io_replay_bits_addr(MSHR_75_3887_io_replay_bits_addr),
    .io_replay_bits_tag(MSHR_75_3887_io_replay_bits_tag),
    .io_replay_bits_cmd(MSHR_75_3887_io_replay_bits_cmd),
    .io_replay_bits_typ(MSHR_75_3887_io_replay_bits_typ),
    .io_replay_bits_phys(MSHR_75_3887_io_replay_bits_phys),
    .io_replay_bits_sdq_id(MSHR_75_3887_io_replay_bits_sdq_id),
    .io_mem_grant_valid(MSHR_75_3887_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(MSHR_75_3887_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(MSHR_75_3887_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(MSHR_75_3887_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(MSHR_75_3887_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(MSHR_75_3887_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(MSHR_75_3887_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(MSHR_75_3887_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(MSHR_75_3887_io_mem_finish_ready),
    .io_mem_finish_valid(MSHR_75_3887_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(MSHR_75_3887_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(MSHR_75_3887_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(MSHR_75_3887_io_wb_req_ready),
    .io_wb_req_valid(MSHR_75_3887_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(MSHR_75_3887_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(MSHR_75_3887_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(MSHR_75_3887_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(MSHR_75_3887_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(MSHR_75_3887_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(MSHR_75_3887_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(MSHR_75_3887_io_wb_req_bits_way_en),
    .io_probe_rdy(MSHR_75_3887_io_probe_rdy)
  );
  Arbiter_78 mmio_alloc_arb (
    .clk(mmio_alloc_arb_clk),
    .reset(mmio_alloc_arb_reset),
    .io_in_0_ready(mmio_alloc_arb_io_in_0_ready),
    .io_in_0_valid(mmio_alloc_arb_io_in_0_valid),
    .io_in_0_bits(mmio_alloc_arb_io_in_0_bits),
    .io_out_ready(mmio_alloc_arb_io_out_ready),
    .io_out_valid(mmio_alloc_arb_io_out_valid),
    .io_out_bits(mmio_alloc_arb_io_out_bits),
    .io_chosen(mmio_alloc_arb_io_chosen)
  );
  Arbiter_79 resp_arb (
    .clk(resp_arb_clk),
    .reset(resp_arb_reset),
    .io_in_0_ready(resp_arb_io_in_0_ready),
    .io_in_0_valid(resp_arb_io_in_0_valid),
    .io_in_0_bits_addr(resp_arb_io_in_0_bits_addr),
    .io_in_0_bits_tag(resp_arb_io_in_0_bits_tag),
    .io_in_0_bits_cmd(resp_arb_io_in_0_bits_cmd),
    .io_in_0_bits_typ(resp_arb_io_in_0_bits_typ),
    .io_in_0_bits_data(resp_arb_io_in_0_bits_data),
    .io_in_0_bits_replay(resp_arb_io_in_0_bits_replay),
    .io_in_0_bits_has_data(resp_arb_io_in_0_bits_has_data),
    .io_in_0_bits_data_word_bypass(resp_arb_io_in_0_bits_data_word_bypass),
    .io_in_0_bits_store_data(resp_arb_io_in_0_bits_store_data),
    .io_out_ready(resp_arb_io_out_ready),
    .io_out_valid(resp_arb_io_out_valid),
    .io_out_bits_addr(resp_arb_io_out_bits_addr),
    .io_out_bits_tag(resp_arb_io_out_bits_tag),
    .io_out_bits_cmd(resp_arb_io_out_bits_cmd),
    .io_out_bits_typ(resp_arb_io_out_bits_typ),
    .io_out_bits_data(resp_arb_io_out_bits_data),
    .io_out_bits_replay(resp_arb_io_out_bits_replay),
    .io_out_bits_has_data(resp_arb_io_out_bits_has_data),
    .io_out_bits_data_word_bypass(resp_arb_io_out_bits_data_word_bypass),
    .io_out_bits_store_data(resp_arb_io_out_bits_store_data),
    .io_chosen(resp_arb_io_chosen)
  );
  IOMSHR IOMSHR_3987 (
    .clk(IOMSHR_3987_clk),
    .reset(IOMSHR_3987_reset),
    .io_req_ready(IOMSHR_3987_io_req_ready),
    .io_req_valid(IOMSHR_3987_io_req_valid),
    .io_req_bits_addr(IOMSHR_3987_io_req_bits_addr),
    .io_req_bits_tag(IOMSHR_3987_io_req_bits_tag),
    .io_req_bits_cmd(IOMSHR_3987_io_req_bits_cmd),
    .io_req_bits_typ(IOMSHR_3987_io_req_bits_typ),
    .io_req_bits_phys(IOMSHR_3987_io_req_bits_phys),
    .io_req_bits_data(IOMSHR_3987_io_req_bits_data),
    .io_acquire_ready(IOMSHR_3987_io_acquire_ready),
    .io_acquire_valid(IOMSHR_3987_io_acquire_valid),
    .io_acquire_bits_addr_block(IOMSHR_3987_io_acquire_bits_addr_block),
    .io_acquire_bits_client_xact_id(IOMSHR_3987_io_acquire_bits_client_xact_id),
    .io_acquire_bits_addr_beat(IOMSHR_3987_io_acquire_bits_addr_beat),
    .io_acquire_bits_is_builtin_type(IOMSHR_3987_io_acquire_bits_is_builtin_type),
    .io_acquire_bits_a_type(IOMSHR_3987_io_acquire_bits_a_type),
    .io_acquire_bits_union(IOMSHR_3987_io_acquire_bits_union),
    .io_acquire_bits_data(IOMSHR_3987_io_acquire_bits_data),
    .io_grant_valid(IOMSHR_3987_io_grant_valid),
    .io_grant_bits_addr_beat(IOMSHR_3987_io_grant_bits_addr_beat),
    .io_grant_bits_client_xact_id(IOMSHR_3987_io_grant_bits_client_xact_id),
    .io_grant_bits_manager_xact_id(IOMSHR_3987_io_grant_bits_manager_xact_id),
    .io_grant_bits_is_builtin_type(IOMSHR_3987_io_grant_bits_is_builtin_type),
    .io_grant_bits_g_type(IOMSHR_3987_io_grant_bits_g_type),
    .io_grant_bits_data(IOMSHR_3987_io_grant_bits_data),
    .io_grant_bits_manager_id(IOMSHR_3987_io_grant_bits_manager_id),
    .io_finish_ready(IOMSHR_3987_io_finish_ready),
    .io_finish_valid(IOMSHR_3987_io_finish_valid),
    .io_finish_bits_manager_xact_id(IOMSHR_3987_io_finish_bits_manager_xact_id),
    .io_finish_bits_manager_id(IOMSHR_3987_io_finish_bits_manager_id),
    .io_resp_ready(IOMSHR_3987_io_resp_ready),
    .io_resp_valid(IOMSHR_3987_io_resp_valid),
    .io_resp_bits_addr(IOMSHR_3987_io_resp_bits_addr),
    .io_resp_bits_tag(IOMSHR_3987_io_resp_bits_tag),
    .io_resp_bits_cmd(IOMSHR_3987_io_resp_bits_cmd),
    .io_resp_bits_typ(IOMSHR_3987_io_resp_bits_typ),
    .io_resp_bits_data(IOMSHR_3987_io_resp_bits_data),
    .io_resp_bits_replay(IOMSHR_3987_io_resp_bits_replay),
    .io_resp_bits_has_data(IOMSHR_3987_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(IOMSHR_3987_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(IOMSHR_3987_io_resp_bits_store_data),
    .io_replay_next(IOMSHR_3987_io_replay_next)
  );
  assign io_req_ready = T_4003;
  assign io_resp_valid = resp_arb_io_out_valid;
  assign io_resp_bits_addr = resp_arb_io_out_bits_addr;
  assign io_resp_bits_tag = resp_arb_io_out_bits_tag;
  assign io_resp_bits_cmd = resp_arb_io_out_bits_cmd;
  assign io_resp_bits_typ = resp_arb_io_out_bits_typ;
  assign io_resp_bits_data = resp_arb_io_out_bits_data;
  assign io_resp_bits_replay = resp_arb_io_out_bits_replay;
  assign io_resp_bits_has_data = resp_arb_io_out_bits_has_data;
  assign io_resp_bits_data_word_bypass = resp_arb_io_out_bits_data_word_bypass;
  assign io_resp_bits_store_data = resp_arb_io_out_bits_store_data;
  assign io_secondary_miss = idx_match;
  assign io_mem_req_valid = mem_req_arb_io_out_valid;
  assign io_mem_req_bits_addr_block = mem_req_arb_io_out_bits_addr_block;
  assign io_mem_req_bits_client_xact_id = mem_req_arb_io_out_bits_client_xact_id;
  assign io_mem_req_bits_addr_beat = mem_req_arb_io_out_bits_addr_beat;
  assign io_mem_req_bits_is_builtin_type = mem_req_arb_io_out_bits_is_builtin_type;
  assign io_mem_req_bits_a_type = mem_req_arb_io_out_bits_a_type;
  assign io_mem_req_bits_union = mem_req_arb_io_out_bits_union;
  assign io_mem_req_bits_data = mem_req_arb_io_out_bits_data;
  assign io_refill_way_en = GEN_0;
  assign io_refill_addr = GEN_1;
  assign io_meta_read_valid = meta_read_arb_io_out_valid;
  assign io_meta_read_bits_idx = meta_read_arb_io_out_bits_idx;
  assign io_meta_read_bits_way_en = meta_read_arb_io_out_bits_way_en;
  assign io_meta_read_bits_tag = meta_read_arb_io_out_bits_tag;
  assign io_meta_write_valid = meta_write_arb_io_out_valid;
  assign io_meta_write_bits_idx = meta_write_arb_io_out_bits_idx;
  assign io_meta_write_bits_way_en = meta_write_arb_io_out_bits_way_en;
  assign io_meta_write_bits_data_tag = meta_write_arb_io_out_bits_data_tag;
  assign io_meta_write_bits_data_coh_state = meta_write_arb_io_out_bits_data_coh_state;
  assign io_replay_valid = replay_arb_io_out_valid;
  assign io_replay_bits_addr = replay_arb_io_out_bits_addr;
  assign io_replay_bits_tag = replay_arb_io_out_bits_tag;
  assign io_replay_bits_cmd = replay_arb_io_out_bits_cmd;
  assign io_replay_bits_typ = replay_arb_io_out_bits_typ;
  assign io_replay_bits_phys = replay_arb_io_out_bits_phys;
  assign io_replay_bits_data = sdq_T_4084_data;
  assign io_mem_finish_valid = mem_finish_arb_io_out_valid;
  assign io_mem_finish_bits_manager_xact_id = mem_finish_arb_io_out_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mem_finish_arb_io_out_bits_manager_id;
  assign io_wb_req_valid = wb_req_arb_io_out_valid;
  assign io_wb_req_bits_addr_beat = wb_req_arb_io_out_bits_addr_beat;
  assign io_wb_req_bits_addr_block = wb_req_arb_io_out_bits_addr_block;
  assign io_wb_req_bits_client_xact_id = wb_req_arb_io_out_bits_client_xact_id;
  assign io_wb_req_bits_voluntary = wb_req_arb_io_out_bits_voluntary;
  assign io_wb_req_bits_r_type = wb_req_arb_io_out_bits_r_type;
  assign io_wb_req_bits_data = wb_req_arb_io_out_bits_data;
  assign io_wb_req_bits_way_en = wb_req_arb_io_out_bits_way_en;
  assign io_probe_rdy = GEN_10;
  assign io_fence_rdy = GEN_11;
  assign io_replay_next = GEN_12;
  assign GEN_17 = {{8'd0}, 32'h80000000};
  assign T_2615 = GEN_17 <= io_req_bits_addr;
  assign GEN_18 = {{7'd0}, 33'h100000000};
  assign T_2617 = io_req_bits_addr < GEN_18;
  assign T_2618 = T_2615 & T_2617;
  assign T_2622 = ~ sdq_val;
  assign T_2623 = T_2622[0];
  assign T_2624 = T_2622[1];
  assign T_2625 = T_2622[2];
  assign T_2626 = T_2622[3];
  assign T_2627 = T_2622[4];
  assign T_2628 = T_2622[5];
  assign T_2629 = T_2622[6];
  assign T_2630 = T_2622[7];
  assign T_2631 = T_2622[8];
  assign T_2632 = T_2622[9];
  assign T_2633 = T_2622[10];
  assign T_2634 = T_2622[11];
  assign T_2635 = T_2622[12];
  assign T_2636 = T_2622[13];
  assign T_2637 = T_2622[14];
  assign T_2638 = T_2622[15];
  assign T_2639 = T_2622[16];
  assign T_2657 = T_2638 ? {{1'd0}, 4'hf} : 5'h10;
  assign T_2658 = T_2637 ? {{1'd0}, 4'he} : T_2657;
  assign T_2659 = T_2636 ? {{1'd0}, 4'hd} : T_2658;
  assign T_2660 = T_2635 ? {{1'd0}, 4'hc} : T_2659;
  assign T_2661 = T_2634 ? {{1'd0}, 4'hb} : T_2660;
  assign T_2662 = T_2633 ? {{1'd0}, 4'ha} : T_2661;
  assign T_2663 = T_2632 ? {{1'd0}, 4'h9} : T_2662;
  assign T_2664 = T_2631 ? {{1'd0}, 4'h8} : T_2663;
  assign T_2665 = T_2630 ? {{2'd0}, 3'h7} : T_2664;
  assign T_2666 = T_2629 ? {{2'd0}, 3'h6} : T_2665;
  assign T_2667 = T_2628 ? {{2'd0}, 3'h5} : T_2666;
  assign T_2668 = T_2627 ? {{2'd0}, 3'h4} : T_2667;
  assign T_2669 = T_2626 ? {{3'd0}, 2'h3} : T_2668;
  assign T_2670 = T_2625 ? {{3'd0}, 2'h2} : T_2669;
  assign T_2671 = T_2624 ? {{4'd0}, 1'h1} : T_2670;
  assign sdq_alloc_id = T_2623 ? {{4'd0}, 1'h0} : T_2671;
  assign GEN_19 = {{16'd0}, 1'h0};
  assign T_2674 = T_2622 == GEN_19;
  assign sdq_rdy = T_2674 == 1'h0;
  assign T_2676 = io_req_valid & io_req_ready;
  assign T_2677 = T_2676 & T_2618;
  assign T_2678 = io_req_bits_cmd == 5'h1;
  assign T_2679 = io_req_bits_cmd == 5'h7;
  assign T_2680 = T_2678 | T_2679;
  assign T_2681 = io_req_bits_cmd[3];
  assign T_2682 = io_req_bits_cmd == 5'h4;
  assign T_2683 = T_2681 | T_2682;
  assign T_2684 = T_2680 | T_2683;
  assign sdq_enq = T_2677 & T_2684;
  assign sdq_T_4084_addr = T_4083;
  assign sdq_T_4084_en = 1'h1;
  `ifdef SYNTHESIS
  assign sdq_T_4084_data = sdq[sdq_T_4084_addr];
  `else
  assign sdq_T_4084_data = sdq_T_4084_addr >= 5'h11 ? $random : sdq[sdq_T_4084_addr];
  `endif
  assign sdq_T_2686_data = io_req_bits_data;
  assign sdq_T_2686_addr = sdq_alloc_id;
  assign sdq_T_2686_mask = sdq_enq;
  assign sdq_T_2686_en = sdq_enq;
  assign idxMatch_0 = MSHR_3871_io_idx_match;
  assign idxMatch_1 = MSHR_75_3887_io_idx_match;
  assign tagList_0 = MSHR_3871_io_tag;
  assign tagList_1 = MSHR_75_3887_io_tag;
  assign T_2702 = idxMatch_0 ? tagList_0 : {{19'd0}, 1'h0};
  assign T_2704 = idxMatch_1 ? tagList_1 : {{19'd0}, 1'h0};
  assign T_2706 = T_2702 | T_2704;
  assign T_2707 = T_2706;
  assign T_2708 = io_req_bits_addr[39:12];
  assign GEN_20 = {{8'd0}, T_2707};
  assign tag_match = GEN_20 == T_2708;
  assign wbTagList_0 = T_3872;
  assign wbTagList_1 = T_3888;
  assign refillMux_0_way_en = MSHR_3871_io_refill_way_en;
  assign refillMux_0_addr = MSHR_3871_io_refill_addr;
  assign refillMux_1_way_en = MSHR_75_3887_io_refill_way_en;
  assign refillMux_1_addr = MSHR_75_3887_io_refill_addr;
  assign meta_read_arb_clk = clk;
  assign meta_read_arb_reset = reset;
  assign meta_read_arb_io_in_0_valid = MSHR_3871_io_meta_read_valid;
  assign meta_read_arb_io_in_0_bits_idx = MSHR_3871_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_0_bits_way_en = MSHR_3871_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_0_bits_tag = MSHR_3871_io_meta_read_bits_tag;
  assign meta_read_arb_io_in_1_valid = MSHR_75_3887_io_meta_read_valid;
  assign meta_read_arb_io_in_1_bits_idx = MSHR_75_3887_io_meta_read_bits_idx;
  assign meta_read_arb_io_in_1_bits_way_en = MSHR_75_3887_io_meta_read_bits_way_en;
  assign meta_read_arb_io_in_1_bits_tag = MSHR_75_3887_io_meta_read_bits_tag;
  assign meta_read_arb_io_out_ready = io_meta_read_ready;
  assign meta_write_arb_clk = clk;
  assign meta_write_arb_reset = reset;
  assign meta_write_arb_io_in_0_valid = MSHR_3871_io_meta_write_valid;
  assign meta_write_arb_io_in_0_bits_idx = MSHR_3871_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_0_bits_way_en = MSHR_3871_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_0_bits_data_tag = MSHR_3871_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_0_bits_data_coh_state = MSHR_3871_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_in_1_valid = MSHR_75_3887_io_meta_write_valid;
  assign meta_write_arb_io_in_1_bits_idx = MSHR_75_3887_io_meta_write_bits_idx;
  assign meta_write_arb_io_in_1_bits_way_en = MSHR_75_3887_io_meta_write_bits_way_en;
  assign meta_write_arb_io_in_1_bits_data_tag = MSHR_75_3887_io_meta_write_bits_data_tag;
  assign meta_write_arb_io_in_1_bits_data_coh_state = MSHR_75_3887_io_meta_write_bits_data_coh_state;
  assign meta_write_arb_io_out_ready = io_meta_write_ready;
  assign mem_req_arb_clk = clk;
  assign mem_req_arb_reset = reset;
  assign mem_req_arb_io_in_0_valid = MSHR_3871_io_mem_req_valid;
  assign mem_req_arb_io_in_0_bits_addr_block = MSHR_3871_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_0_bits_client_xact_id = MSHR_3871_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_0_bits_addr_beat = MSHR_3871_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_0_bits_is_builtin_type = MSHR_3871_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_0_bits_a_type = MSHR_3871_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_0_bits_union = MSHR_3871_io_mem_req_bits_union;
  assign mem_req_arb_io_in_0_bits_data = MSHR_3871_io_mem_req_bits_data;
  assign mem_req_arb_io_in_1_valid = MSHR_75_3887_io_mem_req_valid;
  assign mem_req_arb_io_in_1_bits_addr_block = MSHR_75_3887_io_mem_req_bits_addr_block;
  assign mem_req_arb_io_in_1_bits_client_xact_id = MSHR_75_3887_io_mem_req_bits_client_xact_id;
  assign mem_req_arb_io_in_1_bits_addr_beat = MSHR_75_3887_io_mem_req_bits_addr_beat;
  assign mem_req_arb_io_in_1_bits_is_builtin_type = MSHR_75_3887_io_mem_req_bits_is_builtin_type;
  assign mem_req_arb_io_in_1_bits_a_type = MSHR_75_3887_io_mem_req_bits_a_type;
  assign mem_req_arb_io_in_1_bits_union = MSHR_75_3887_io_mem_req_bits_union;
  assign mem_req_arb_io_in_1_bits_data = MSHR_75_3887_io_mem_req_bits_data;
  assign mem_req_arb_io_in_2_valid = IOMSHR_3987_io_acquire_valid;
  assign mem_req_arb_io_in_2_bits_addr_block = IOMSHR_3987_io_acquire_bits_addr_block;
  assign mem_req_arb_io_in_2_bits_client_xact_id = IOMSHR_3987_io_acquire_bits_client_xact_id;
  assign mem_req_arb_io_in_2_bits_addr_beat = IOMSHR_3987_io_acquire_bits_addr_beat;
  assign mem_req_arb_io_in_2_bits_is_builtin_type = IOMSHR_3987_io_acquire_bits_is_builtin_type;
  assign mem_req_arb_io_in_2_bits_a_type = IOMSHR_3987_io_acquire_bits_a_type;
  assign mem_req_arb_io_in_2_bits_union = IOMSHR_3987_io_acquire_bits_union;
  assign mem_req_arb_io_in_2_bits_data = IOMSHR_3987_io_acquire_bits_data;
  assign mem_req_arb_io_out_ready = io_mem_req_ready;
  assign mem_finish_arb_clk = clk;
  assign mem_finish_arb_reset = reset;
  assign mem_finish_arb_io_in_0_valid = MSHR_3871_io_mem_finish_valid;
  assign mem_finish_arb_io_in_0_bits_manager_xact_id = MSHR_3871_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_0_bits_manager_id = MSHR_3871_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_1_valid = MSHR_75_3887_io_mem_finish_valid;
  assign mem_finish_arb_io_in_1_bits_manager_xact_id = MSHR_75_3887_io_mem_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_1_bits_manager_id = MSHR_75_3887_io_mem_finish_bits_manager_id;
  assign mem_finish_arb_io_in_2_valid = IOMSHR_3987_io_finish_valid;
  assign mem_finish_arb_io_in_2_bits_manager_xact_id = IOMSHR_3987_io_finish_bits_manager_xact_id;
  assign mem_finish_arb_io_in_2_bits_manager_id = IOMSHR_3987_io_finish_bits_manager_id;
  assign mem_finish_arb_io_out_ready = io_mem_finish_ready;
  assign wb_req_arb_clk = clk;
  assign wb_req_arb_reset = reset;
  assign wb_req_arb_io_in_0_valid = MSHR_3871_io_wb_req_valid;
  assign wb_req_arb_io_in_0_bits_addr_beat = MSHR_3871_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_0_bits_addr_block = MSHR_3871_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_0_bits_client_xact_id = MSHR_3871_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_0_bits_voluntary = MSHR_3871_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_0_bits_r_type = MSHR_3871_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_0_bits_data = MSHR_3871_io_wb_req_bits_data;
  assign wb_req_arb_io_in_0_bits_way_en = MSHR_3871_io_wb_req_bits_way_en;
  assign wb_req_arb_io_in_1_valid = MSHR_75_3887_io_wb_req_valid;
  assign wb_req_arb_io_in_1_bits_addr_beat = MSHR_75_3887_io_wb_req_bits_addr_beat;
  assign wb_req_arb_io_in_1_bits_addr_block = MSHR_75_3887_io_wb_req_bits_addr_block;
  assign wb_req_arb_io_in_1_bits_client_xact_id = MSHR_75_3887_io_wb_req_bits_client_xact_id;
  assign wb_req_arb_io_in_1_bits_voluntary = MSHR_75_3887_io_wb_req_bits_voluntary;
  assign wb_req_arb_io_in_1_bits_r_type = MSHR_75_3887_io_wb_req_bits_r_type;
  assign wb_req_arb_io_in_1_bits_data = MSHR_75_3887_io_wb_req_bits_data;
  assign wb_req_arb_io_in_1_bits_way_en = MSHR_75_3887_io_wb_req_bits_way_en;
  assign wb_req_arb_io_out_ready = io_wb_req_ready;
  assign replay_arb_clk = clk;
  assign replay_arb_reset = reset;
  assign replay_arb_io_in_0_valid = MSHR_3871_io_replay_valid;
  assign replay_arb_io_in_0_bits_addr = MSHR_3871_io_replay_bits_addr;
  assign replay_arb_io_in_0_bits_tag = MSHR_3871_io_replay_bits_tag;
  assign replay_arb_io_in_0_bits_cmd = MSHR_3871_io_replay_bits_cmd;
  assign replay_arb_io_in_0_bits_typ = MSHR_3871_io_replay_bits_typ;
  assign replay_arb_io_in_0_bits_phys = MSHR_3871_io_replay_bits_phys;
  assign replay_arb_io_in_0_bits_sdq_id = MSHR_3871_io_replay_bits_sdq_id;
  assign replay_arb_io_in_1_valid = MSHR_75_3887_io_replay_valid;
  assign replay_arb_io_in_1_bits_addr = MSHR_75_3887_io_replay_bits_addr;
  assign replay_arb_io_in_1_bits_tag = MSHR_75_3887_io_replay_bits_tag;
  assign replay_arb_io_in_1_bits_cmd = MSHR_75_3887_io_replay_bits_cmd;
  assign replay_arb_io_in_1_bits_typ = MSHR_75_3887_io_replay_bits_typ;
  assign replay_arb_io_in_1_bits_phys = MSHR_75_3887_io_replay_bits_phys;
  assign replay_arb_io_in_1_bits_sdq_id = MSHR_75_3887_io_replay_bits_sdq_id;
  assign replay_arb_io_out_ready = io_replay_ready;
  assign alloc_arb_clk = clk;
  assign alloc_arb_reset = reset;
  assign alloc_arb_io_in_0_valid = MSHR_3871_io_req_pri_rdy;
  assign alloc_arb_io_in_0_bits = GEN_2;
  assign alloc_arb_io_in_1_valid = MSHR_75_3887_io_req_pri_rdy;
  assign alloc_arb_io_in_1_bits = GEN_3;
  assign alloc_arb_io_out_ready = T_3904;
  assign MSHR_3871_clk = clk;
  assign MSHR_3871_reset = reset;
  assign MSHR_3871_io_req_pri_val = alloc_arb_io_in_0_ready;
  assign MSHR_3871_io_req_sec_val = T_3874;
  assign MSHR_3871_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_3871_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_3871_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_3871_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_3871_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_3871_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_3871_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_3871_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_3871_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_3871_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_3871_io_mem_req_ready = mem_req_arb_io_in_0_ready;
  assign MSHR_3871_io_meta_read_ready = meta_read_arb_io_in_0_ready;
  assign MSHR_3871_io_meta_write_ready = meta_write_arb_io_in_0_ready;
  assign MSHR_3871_io_replay_ready = replay_arb_io_in_0_ready;
  assign MSHR_3871_io_mem_grant_valid = T_3877;
  assign MSHR_3871_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_3871_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_3871_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_3871_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_3871_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_3871_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_3871_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_3871_io_mem_finish_ready = mem_finish_arb_io_in_0_ready;
  assign MSHR_3871_io_wb_req_ready = wb_req_arb_io_in_0_ready;
  assign T_3872 = MSHR_3871_io_wb_req_bits_addr_block[25:6];
  assign T_3873 = io_req_valid & sdq_rdy;
  assign T_3874 = T_3873 & tag_match;
  assign GEN_21 = {{1'd0}, 1'h0};
  assign T_3876 = io_mem_grant_bits_client_xact_id == GEN_21;
  assign T_3877 = io_mem_grant_valid & T_3876;
  assign T_3878 = MSHR_3871_io_req_pri_rdy;
  assign T_3879 = MSHR_3871_io_req_sec_rdy;
  assign T_3880 = MSHR_3871_io_idx_match;
  assign T_3882 = MSHR_3871_io_req_pri_rdy == 1'h0;
  assign GEN_7 = T_3882 ? 1'h0 : 1'h1;
  assign T_3885 = MSHR_3871_io_probe_rdy == 1'h0;
  assign GEN_8 = T_3885 ? 1'h0 : 1'h1;
  assign MSHR_75_3887_clk = clk;
  assign MSHR_75_3887_reset = reset;
  assign MSHR_75_3887_io_req_pri_val = alloc_arb_io_in_1_ready;
  assign MSHR_75_3887_io_req_sec_val = T_3874;
  assign MSHR_75_3887_io_req_bits_addr = io_req_bits_addr;
  assign MSHR_75_3887_io_req_bits_tag = io_req_bits_tag;
  assign MSHR_75_3887_io_req_bits_cmd = io_req_bits_cmd;
  assign MSHR_75_3887_io_req_bits_typ = io_req_bits_typ;
  assign MSHR_75_3887_io_req_bits_phys = io_req_bits_phys;
  assign MSHR_75_3887_io_req_bits_sdq_id = sdq_alloc_id;
  assign MSHR_75_3887_io_req_bits_tag_match = io_req_bits_tag_match;
  assign MSHR_75_3887_io_req_bits_old_meta_tag = io_req_bits_old_meta_tag;
  assign MSHR_75_3887_io_req_bits_old_meta_coh_state = io_req_bits_old_meta_coh_state;
  assign MSHR_75_3887_io_req_bits_way_en = io_req_bits_way_en;
  assign MSHR_75_3887_io_mem_req_ready = mem_req_arb_io_in_1_ready;
  assign MSHR_75_3887_io_meta_read_ready = meta_read_arb_io_in_1_ready;
  assign MSHR_75_3887_io_meta_write_ready = meta_write_arb_io_in_1_ready;
  assign MSHR_75_3887_io_replay_ready = replay_arb_io_in_1_ready;
  assign MSHR_75_3887_io_mem_grant_valid = T_3893;
  assign MSHR_75_3887_io_mem_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign MSHR_75_3887_io_mem_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign MSHR_75_3887_io_mem_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign MSHR_75_3887_io_mem_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign MSHR_75_3887_io_mem_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign MSHR_75_3887_io_mem_grant_bits_data = io_mem_grant_bits_data;
  assign MSHR_75_3887_io_mem_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign MSHR_75_3887_io_mem_finish_ready = mem_finish_arb_io_in_1_ready;
  assign MSHR_75_3887_io_wb_req_ready = wb_req_arb_io_in_1_ready;
  assign T_3888 = MSHR_75_3887_io_wb_req_bits_addr_block[25:6];
  assign GEN_22 = {{1'd0}, 1'h1};
  assign T_3892 = io_mem_grant_bits_client_xact_id == GEN_22;
  assign T_3893 = io_mem_grant_valid & T_3892;
  assign pri_rdy = T_3878 | MSHR_75_3887_io_req_pri_rdy;
  assign sec_rdy = T_3879 | MSHR_75_3887_io_req_sec_rdy;
  assign idx_match = T_3880 | MSHR_75_3887_io_idx_match;
  assign T_3895 = MSHR_75_3887_io_req_pri_rdy == 1'h0;
  assign GEN_9 = T_3895 ? 1'h0 : GEN_7;
  assign T_3898 = MSHR_75_3887_io_probe_rdy == 1'h0;
  assign GEN_10 = T_3898 ? 1'h0 : GEN_8;
  assign T_3901 = T_3873 & T_2618;
  assign T_3903 = idx_match == 1'h0;
  assign T_3904 = T_3901 & T_3903;
  assign mmio_alloc_arb_clk = clk;
  assign mmio_alloc_arb_reset = reset;
  assign mmio_alloc_arb_io_in_0_valid = IOMSHR_3987_io_req_ready;
  assign mmio_alloc_arb_io_in_0_bits = GEN_4;
  assign mmio_alloc_arb_io_out_ready = T_3997;
  assign resp_arb_clk = clk;
  assign resp_arb_reset = reset;
  assign resp_arb_io_in_0_valid = IOMSHR_3987_io_resp_valid;
  assign resp_arb_io_in_0_bits_addr = IOMSHR_3987_io_resp_bits_addr;
  assign resp_arb_io_in_0_bits_tag = IOMSHR_3987_io_resp_bits_tag;
  assign resp_arb_io_in_0_bits_cmd = IOMSHR_3987_io_resp_bits_cmd;
  assign resp_arb_io_in_0_bits_typ = IOMSHR_3987_io_resp_bits_typ;
  assign resp_arb_io_in_0_bits_data = IOMSHR_3987_io_resp_bits_data;
  assign resp_arb_io_in_0_bits_replay = IOMSHR_3987_io_resp_bits_replay;
  assign resp_arb_io_in_0_bits_has_data = IOMSHR_3987_io_resp_bits_has_data;
  assign resp_arb_io_in_0_bits_data_word_bypass = IOMSHR_3987_io_resp_bits_data_word_bypass;
  assign resp_arb_io_in_0_bits_store_data = IOMSHR_3987_io_resp_bits_store_data;
  assign resp_arb_io_out_ready = io_resp_ready;
  assign IOMSHR_3987_clk = clk;
  assign IOMSHR_3987_reset = reset;
  assign IOMSHR_3987_io_req_valid = mmio_alloc_arb_io_in_0_ready;
  assign IOMSHR_3987_io_req_bits_addr = io_req_bits_addr;
  assign IOMSHR_3987_io_req_bits_tag = io_req_bits_tag;
  assign IOMSHR_3987_io_req_bits_cmd = io_req_bits_cmd;
  assign IOMSHR_3987_io_req_bits_typ = io_req_bits_typ;
  assign IOMSHR_3987_io_req_bits_phys = io_req_bits_phys;
  assign IOMSHR_3987_io_req_bits_data = io_req_bits_data;
  assign IOMSHR_3987_io_acquire_ready = mem_req_arb_io_in_2_ready;
  assign IOMSHR_3987_io_grant_valid = T_3990;
  assign IOMSHR_3987_io_grant_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign IOMSHR_3987_io_grant_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign IOMSHR_3987_io_grant_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign IOMSHR_3987_io_grant_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign IOMSHR_3987_io_grant_bits_g_type = io_mem_grant_bits_g_type;
  assign IOMSHR_3987_io_grant_bits_data = io_mem_grant_bits_data;
  assign IOMSHR_3987_io_grant_bits_manager_id = io_mem_grant_bits_manager_id;
  assign IOMSHR_3987_io_finish_ready = mem_finish_arb_io_in_2_ready;
  assign IOMSHR_3987_io_resp_ready = resp_arb_io_in_0_ready;
  assign mmio_rdy = IOMSHR_3987_io_req_ready;
  assign T_3989 = io_mem_grant_bits_client_xact_id == 2'h2;
  assign T_3990 = io_mem_grant_valid & T_3989;
  assign T_3992 = IOMSHR_3987_io_req_ready == 1'h0;
  assign GEN_11 = T_3992 ? 1'h0 : GEN_9;
  assign GEN_12 = IOMSHR_3987_io_replay_next;
  assign T_3996 = T_2618 == 1'h0;
  assign T_3997 = io_req_valid & T_3996;
  assign T_4000 = tag_match & sec_rdy;
  assign T_4001 = idx_match ? T_4000 : pri_rdy;
  assign T_4002 = T_4001 & sdq_rdy;
  assign T_4003 = T_3996 ? mmio_rdy : T_4002;
  assign GEN_0 = GEN_13;
  assign GEN_13 = GEN_22 == io_mem_grant_bits_client_xact_id ? refillMux_1_way_en : refillMux_0_way_en;
  assign GEN_1 = GEN_14;
  assign GEN_14 = GEN_22 == io_mem_grant_bits_client_xact_id ? refillMux_1_addr : refillMux_0_addr;
  assign T_4075 = io_replay_ready & io_replay_valid;
  assign T_4076 = io_replay_bits_cmd == 5'h1;
  assign T_4077 = io_replay_bits_cmd == 5'h7;
  assign T_4078 = T_4076 | T_4077;
  assign T_4079 = io_replay_bits_cmd[3];
  assign T_4080 = io_replay_bits_cmd == 5'h4;
  assign T_4081 = T_4079 | T_4080;
  assign T_4082 = T_4078 | T_4081;
  assign free_sdq = T_4075 & T_4082;
  assign GEN_15 = free_sdq ? replay_arb_io_out_bits_sdq_id : T_4083;
  assign T_4085 = io_replay_valid | sdq_enq;
  assign GEN_25 = {{31'd0}, 1'h1};
  assign T_4087 = GEN_25 << replay_arb_io_out_bits_sdq_id;
  assign GEN_26 = {{16'd0}, free_sdq};
  assign T_4089 = 17'h0 - GEN_26;
  assign T_4090 = T_4089[16:0];
  assign GEN_27 = {{15'd0}, T_4090};
  assign T_4091 = T_4087 & GEN_27;
  assign T_4092 = ~ T_4091;
  assign GEN_28 = {{15'd0}, sdq_val};
  assign T_4093 = GEN_28 & T_4092;
  assign T_4132 = T_2639 ? 17'h10000 : 17'h0;
  assign T_4133 = T_2638 ? 17'h8000 : T_4132;
  assign T_4134 = T_2637 ? 17'h4000 : T_4133;
  assign T_4135 = T_2636 ? 17'h2000 : T_4134;
  assign T_4136 = T_2635 ? 17'h1000 : T_4135;
  assign T_4137 = T_2634 ? 17'h800 : T_4136;
  assign T_4138 = T_2633 ? 17'h400 : T_4137;
  assign T_4139 = T_2632 ? 17'h200 : T_4138;
  assign T_4140 = T_2631 ? 17'h100 : T_4139;
  assign T_4141 = T_2630 ? 17'h80 : T_4140;
  assign T_4142 = T_2629 ? 17'h40 : T_4141;
  assign T_4143 = T_2628 ? 17'h20 : T_4142;
  assign T_4144 = T_2627 ? 17'h10 : T_4143;
  assign T_4145 = T_2626 ? 17'h8 : T_4144;
  assign T_4146 = T_2625 ? 17'h4 : T_4145;
  assign T_4147 = T_2624 ? 17'h2 : T_4146;
  assign T_4148 = T_2623 ? 17'h1 : T_4147;
  assign GEN_29 = {{16'd0}, sdq_enq};
  assign T_4150 = 17'h0 - GEN_29;
  assign T_4151 = T_4150[16:0];
  assign T_4152 = T_4148 & T_4151;
  assign GEN_30 = {{15'd0}, T_4152};
  assign T_4153 = T_4093 | GEN_30;
  assign GEN_16 = T_4085 ? T_4153 : {{15'd0}, sdq_val};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_5 = {1{$random}};
  sdq_val = GEN_5[16:0];
  GEN_6 = {2{$random}};
  for (initvar = 0; initvar < 17; initvar = initvar+1)
    sdq[initvar] = GEN_6[63:0];
  GEN_23 = {1{$random}};
  T_4083 = GEN_23[4:0];
  GEN_24 = {1{$random}};
  GEN_2 = GEN_24[0:0];
  GEN_31 = {1{$random}};
  GEN_3 = GEN_31[0:0];
  GEN_32 = {1{$random}};
  GEN_4 = GEN_32[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      sdq_val <= 17'h0;
    end else begin
      sdq_val <= GEN_16[16:0];
    end
    if(sdq_T_2686_en & sdq_T_2686_mask) begin
      sdq[sdq_T_2686_addr] <= sdq_T_2686_data;
    end
    if(1'h0) begin
    end else begin
      T_4083 <= GEN_15;
    end
  end
endmodule
module MetadataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [5:0] io_read_bits_idx,
  input  [3:0] io_read_bits_way_en,
  output  io_write_ready,
  input   io_write_valid,
  input  [5:0] io_write_bits_idx,
  input  [3:0] io_write_bits_way_en,
  input  [19:0] io_write_bits_data_tag,
  input  [1:0] io_write_bits_data_coh_state,
  output [19:0] io_resp_0_tag,
  output [1:0] io_resp_0_coh_state,
  output [19:0] io_resp_1_tag,
  output [1:0] io_resp_1_coh_state,
  output [19:0] io_resp_2_tag,
  output [1:0] io_resp_2_coh_state,
  output [19:0] io_resp_3_tag,
  output [1:0] io_resp_3_coh_state
);
  wire [1:0] T_50_state;
  wire [19:0] rstVal_tag;
  wire [1:0] rstVal_coh_state;
  reg [6:0] rst_cnt;
  reg [31:0] GEN_1;
  wire  rst;
  wire [6:0] waddr;
  wire [19:0] T_2358_tag;
  wire [1:0] T_2358_coh_state;
  wire [21:0] wdata;
  wire [3:0] T_2457;
  wire  GEN_25;
  wire [3:0] T_2458;
  wire  T_2459;
  wire  T_2460;
  wire  T_2461;
  wire  T_2462;
  wire [6:0] GEN_27;
  wire [7:0] T_2473;
  wire [6:0] T_2474;
  wire [6:0] GEN_0;
  reg [21:0] T_2483_0 [0:63];
  reg [31:0] GEN_2;
  wire [21:0] T_2483_0_T_2500_data;
  wire [5:0] T_2483_0_T_2500_addr;
  wire  T_2483_0_T_2500_en;
  reg [5:0] GEN_3;
  reg  GEN_4;
  wire [21:0] T_2483_0_T_2494_data;
  wire [5:0] T_2483_0_T_2494_addr;
  wire  T_2483_0_T_2494_mask;
  wire  T_2483_0_T_2494_en;
  reg [21:0] T_2483_1 [0:63];
  reg [31:0] GEN_5;
  wire [21:0] T_2483_1_T_2500_data;
  wire [5:0] T_2483_1_T_2500_addr;
  wire  T_2483_1_T_2500_en;
  reg [5:0] GEN_6;
  reg  GEN_7;
  wire [21:0] T_2483_1_T_2494_data;
  wire [5:0] T_2483_1_T_2494_addr;
  wire  T_2483_1_T_2494_mask;
  wire  T_2483_1_T_2494_en;
  reg [21:0] T_2483_2 [0:63];
  reg [31:0] GEN_8;
  wire [21:0] T_2483_2_T_2500_data;
  wire [5:0] T_2483_2_T_2500_addr;
  wire  T_2483_2_T_2500_en;
  reg [5:0] GEN_9;
  reg  GEN_10;
  wire [21:0] T_2483_2_T_2494_data;
  wire [5:0] T_2483_2_T_2494_addr;
  wire  T_2483_2_T_2494_mask;
  wire  T_2483_2_T_2494_en;
  reg [21:0] T_2483_3 [0:63];
  reg [31:0] GEN_11;
  wire [21:0] T_2483_3_T_2500_data;
  wire [5:0] T_2483_3_T_2500_addr;
  wire  T_2483_3_T_2500_en;
  reg [5:0] GEN_12;
  reg  GEN_13;
  wire [21:0] T_2483_3_T_2494_data;
  wire [5:0] T_2483_3_T_2494_addr;
  wire  T_2483_3_T_2494_mask;
  wire  T_2483_3_T_2494_en;
  wire  T_2484;
  wire [21:0] T_2490_0;
  wire [21:0] T_2490_1;
  wire [21:0] T_2490_2;
  wire [21:0] T_2490_3;
  wire  GEN_17;
  wire  GEN_19;
  wire  GEN_21;
  wire  GEN_23;
  wire [5:0] T_2497;
  wire [43:0] T_2502;
  wire [43:0] T_2503;
  wire [87:0] T_2504;
  wire [19:0] T_3366_0_tag;
  wire [1:0] T_3366_0_coh_state;
  wire [19:0] T_3366_1_tag;
  wire [1:0] T_3366_1_coh_state;
  wire [19:0] T_3366_2_tag;
  wire [1:0] T_3366_2_coh_state;
  wire [19:0] T_3366_3_tag;
  wire [1:0] T_3366_3_coh_state;
  wire [1:0] T_3843;
  wire [19:0] T_3844;
  wire [1:0] T_3845;
  wire [19:0] T_3846;
  wire [1:0] T_3847;
  wire [19:0] T_3848;
  wire [1:0] T_3849;
  wire [19:0] T_3850;
  wire  T_3852;
  wire  T_3854;
  wire  T_3855;
  assign io_read_ready = T_3855;
  assign io_write_ready = T_3852;
  assign io_resp_0_tag = T_3366_0_tag;
  assign io_resp_0_coh_state = T_3366_0_coh_state;
  assign io_resp_1_tag = T_3366_1_tag;
  assign io_resp_1_coh_state = T_3366_1_coh_state;
  assign io_resp_2_tag = T_3366_2_tag;
  assign io_resp_2_coh_state = T_3366_2_coh_state;
  assign io_resp_3_tag = T_3366_3_tag;
  assign io_resp_3_coh_state = T_3366_3_coh_state;
  assign T_50_state = {{1'd0}, 1'h0};
  assign rstVal_tag = {{19'd0}, 1'h0};
  assign rstVal_coh_state = T_50_state;
  assign rst = rst_cnt < 7'h40;
  assign waddr = rst ? rst_cnt : {{1'd0}, io_write_bits_idx};
  assign T_2358_tag = rst ? rstVal_tag : io_write_bits_data_tag;
  assign T_2358_coh_state = rst ? rstVal_coh_state : io_write_bits_data_coh_state;
  assign wdata = {T_2358_tag,T_2358_coh_state};
  assign T_2457 = $signed(io_write_bits_way_en);
  assign GEN_25 = $signed(1'h1);
  assign T_2458 = rst ? $signed({4{GEN_25}}) : $signed(T_2457);
  assign T_2459 = T_2458[0];
  assign T_2460 = T_2458[1];
  assign T_2461 = T_2458[2];
  assign T_2462 = T_2458[3];
  assign GEN_27 = {{6'd0}, 1'h1};
  assign T_2473 = rst_cnt + GEN_27;
  assign T_2474 = T_2473[6:0];
  assign GEN_0 = rst ? T_2474 : rst_cnt;
  assign T_2483_0_T_2500_addr = T_2497;
  assign T_2483_0_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_0_T_2500_data = T_2483_0[GEN_3];
  `else
  assign T_2483_0_T_2500_data = GEN_3 >= 7'h40 ? $random : T_2483_0[GEN_3];
  `endif
  assign T_2483_0_T_2494_data = T_2490_0;
  assign T_2483_0_T_2494_addr = waddr[5:0];
  assign T_2483_0_T_2494_mask = GEN_17;
  assign T_2483_0_T_2494_en = T_2484;
  assign T_2483_1_T_2500_addr = T_2497;
  assign T_2483_1_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_1_T_2500_data = T_2483_1[GEN_6];
  `else
  assign T_2483_1_T_2500_data = GEN_6 >= 7'h40 ? $random : T_2483_1[GEN_6];
  `endif
  assign T_2483_1_T_2494_data = T_2490_1;
  assign T_2483_1_T_2494_addr = waddr[5:0];
  assign T_2483_1_T_2494_mask = GEN_19;
  assign T_2483_1_T_2494_en = T_2484;
  assign T_2483_2_T_2500_addr = T_2497;
  assign T_2483_2_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_2_T_2500_data = T_2483_2[GEN_9];
  `else
  assign T_2483_2_T_2500_data = GEN_9 >= 7'h40 ? $random : T_2483_2[GEN_9];
  `endif
  assign T_2483_2_T_2494_data = T_2490_2;
  assign T_2483_2_T_2494_addr = waddr[5:0];
  assign T_2483_2_T_2494_mask = GEN_21;
  assign T_2483_2_T_2494_en = T_2484;
  assign T_2483_3_T_2500_addr = T_2497;
  assign T_2483_3_T_2500_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_2483_3_T_2500_data = T_2483_3[GEN_12];
  `else
  assign T_2483_3_T_2500_data = GEN_12 >= 7'h40 ? $random : T_2483_3[GEN_12];
  `endif
  assign T_2483_3_T_2494_data = T_2490_3;
  assign T_2483_3_T_2494_addr = waddr[5:0];
  assign T_2483_3_T_2494_mask = GEN_23;
  assign T_2483_3_T_2494_en = T_2484;
  assign T_2484 = rst | io_write_valid;
  assign T_2490_0 = wdata;
  assign T_2490_1 = wdata;
  assign T_2490_2 = wdata;
  assign T_2490_3 = wdata;
  assign GEN_17 = T_2484 ? T_2459 : 1'h0;
  assign GEN_19 = T_2484 ? T_2460 : 1'h0;
  assign GEN_21 = T_2484 ? T_2461 : 1'h0;
  assign GEN_23 = T_2484 ? T_2462 : 1'h0;
  assign T_2497 = io_read_bits_idx;
  assign T_2502 = {T_2483_1_T_2500_data,T_2483_0_T_2500_data};
  assign T_2503 = {T_2483_3_T_2500_data,T_2483_2_T_2500_data};
  assign T_2504 = {T_2503,T_2502};
  assign T_3366_0_tag = T_3844;
  assign T_3366_0_coh_state = T_3843;
  assign T_3366_1_tag = T_3846;
  assign T_3366_1_coh_state = T_3845;
  assign T_3366_2_tag = T_3848;
  assign T_3366_2_coh_state = T_3847;
  assign T_3366_3_tag = T_3850;
  assign T_3366_3_coh_state = T_3849;
  assign T_3843 = T_2504[1:0];
  assign T_3844 = T_2504[21:2];
  assign T_3845 = T_2504[23:22];
  assign T_3846 = T_2504[43:24];
  assign T_3847 = T_2504[45:44];
  assign T_3848 = T_2504[65:46];
  assign T_3849 = T_2504[67:66];
  assign T_3850 = T_2504[87:68];
  assign T_3852 = rst == 1'h0;
  assign T_3854 = io_write_valid == 1'h0;
  assign T_3855 = T_3852 & T_3854;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  rst_cnt = GEN_1[6:0];
  GEN_2 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_0[initvar] = GEN_2[21:0];
  GEN_5 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_1[initvar] = GEN_5[21:0];
  GEN_8 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_2[initvar] = GEN_8[21:0];
  GEN_11 = {1{$random}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    T_2483_3[initvar] = GEN_11[21:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      rst_cnt <= 7'h0;
    end else begin
      rst_cnt <= GEN_0;
    end
    GEN_3 <= T_2483_0_T_2500_addr;
    GEN_4 <= T_2483_0_T_2500_en;
    if(T_2483_0_T_2494_en & T_2483_0_T_2494_mask) begin
      T_2483_0[T_2483_0_T_2494_addr] <= T_2483_0_T_2494_data;
    end
    GEN_6 <= T_2483_1_T_2500_addr;
    GEN_7 <= T_2483_1_T_2500_en;
    if(T_2483_1_T_2494_en & T_2483_1_T_2494_mask) begin
      T_2483_1[T_2483_1_T_2494_addr] <= T_2483_1_T_2494_data;
    end
    GEN_9 <= T_2483_2_T_2500_addr;
    GEN_10 <= T_2483_2_T_2500_en;
    if(T_2483_2_T_2494_en & T_2483_2_T_2494_mask) begin
      T_2483_2[T_2483_2_T_2494_addr] <= T_2483_2_T_2494_data;
    end
    GEN_12 <= T_2483_3_T_2500_addr;
    GEN_13 <= T_2483_3_T_2500_en;
    if(T_2483_3_T_2494_en & T_2483_3_T_2494_mask) begin
      T_2483_3[T_2483_3_T_2494_addr] <= T_2483_3_T_2494_data;
    end
  end
endmodule
module Arbiter_83(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [5:0] io_in_0_bits_idx,
  input  [3:0] io_in_0_bits_way_en,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [5:0] io_in_1_bits_idx,
  input  [3:0] io_in_1_bits_way_en,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [5:0] io_in_2_bits_idx,
  input  [3:0] io_in_2_bits_way_en,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [5:0] io_in_3_bits_idx,
  input  [3:0] io_in_3_bits_way_en,
  output  io_in_4_ready,
  input   io_in_4_valid,
  input  [5:0] io_in_4_bits_idx,
  input  [3:0] io_in_4_bits_way_en,
  input   io_out_ready,
  output  io_out_valid,
  output [5:0] io_out_bits_idx,
  output [3:0] io_out_bits_way_en,
  output [2:0] io_chosen
);
  wire [2:0] GEN_0;
  wire [5:0] GEN_1;
  wire [3:0] GEN_2;
  wire [2:0] GEN_3;
  wire [5:0] GEN_4;
  wire [3:0] GEN_5;
  wire [2:0] GEN_6;
  wire [5:0] GEN_7;
  wire [3:0] GEN_8;
  wire [2:0] GEN_9;
  wire [5:0] GEN_10;
  wire [3:0] GEN_11;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_938;
  wire  T_940;
  wire  T_942;
  wire  T_944;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire  T_949;
  wire  T_951;
  wire  T_952;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_946;
  assign io_in_2_ready = T_947;
  assign io_in_3_ready = T_948;
  assign io_in_4_ready = T_949;
  assign io_out_valid = T_952;
  assign io_out_bits_idx = GEN_10;
  assign io_out_bits_way_en = GEN_11;
  assign io_chosen = GEN_9;
  assign GEN_0 = io_in_3_valid ? {{1'd0}, 2'h3} : 3'h4;
  assign GEN_1 = io_in_3_valid ? io_in_3_bits_idx : io_in_4_bits_idx;
  assign GEN_2 = io_in_3_valid ? io_in_3_bits_way_en : io_in_4_bits_way_en;
  assign GEN_3 = io_in_2_valid ? {{1'd0}, 2'h2} : GEN_0;
  assign GEN_4 = io_in_2_valid ? io_in_2_bits_idx : GEN_1;
  assign GEN_5 = io_in_2_valid ? io_in_2_bits_way_en : GEN_2;
  assign GEN_6 = io_in_1_valid ? {{2'd0}, 1'h1} : GEN_3;
  assign GEN_7 = io_in_1_valid ? io_in_1_bits_idx : GEN_4;
  assign GEN_8 = io_in_1_valid ? io_in_1_bits_way_en : GEN_5;
  assign GEN_9 = io_in_0_valid ? {{2'd0}, 1'h0} : GEN_6;
  assign GEN_10 = io_in_0_valid ? io_in_0_bits_idx : GEN_7;
  assign GEN_11 = io_in_0_valid ? io_in_0_bits_way_en : GEN_8;
  assign T_934 = io_in_0_valid | io_in_1_valid;
  assign T_935 = T_934 | io_in_2_valid;
  assign T_936 = T_935 | io_in_3_valid;
  assign T_938 = io_in_0_valid == 1'h0;
  assign T_940 = T_934 == 1'h0;
  assign T_942 = T_935 == 1'h0;
  assign T_944 = T_936 == 1'h0;
  assign T_946 = T_938 & io_out_ready;
  assign T_947 = T_940 & io_out_ready;
  assign T_948 = T_942 & io_out_ready;
  assign T_949 = T_944 & io_out_ready;
  assign T_951 = T_944 == 1'h0;
  assign T_952 = T_951 | io_in_4_valid;
endmodule
module DataArray(
  input   clk,
  input   reset,
  output  io_read_ready,
  input   io_read_valid,
  input  [3:0] io_read_bits_way_en,
  input  [11:0] io_read_bits_addr,
  output  io_write_ready,
  input   io_write_valid,
  input  [3:0] io_write_bits_way_en,
  input  [11:0] io_write_bits_addr,
  input   io_write_bits_wmask,
  input  [63:0] io_write_bits_data,
  output [63:0] io_resp_0,
  output [63:0] io_resp_1,
  output [63:0] io_resp_2,
  output [63:0] io_resp_3
);
  wire [8:0] waddr;
  wire [8:0] raddr;
  wire  T_815;
  wire [63:0] T_823_0;
  reg [11:0] T_825;
  reg [31:0] GEN_1;
  wire [11:0] GEN_0;
  reg [63:0] T_834_0 [0:511];
  reg [63:0] GEN_2;
  wire [63:0] T_834_0_T_860_data;
  wire [8:0] T_834_0_T_860_addr;
  wire  T_834_0_T_860_en;
  reg [8:0] GEN_3;
  reg  GEN_4;
  wire [63:0] T_834_0_T_851_data;
  wire [8:0] T_834_0_T_851_addr;
  wire  T_834_0_T_851_mask;
  wire  T_834_0_T_851_en;
  wire  T_837;
  wire  T_839;
  wire [63:0] T_846_0;
  wire  GEN_8;
  wire [8:0] T_857;
  wire [63:0] T_868_0;
  wire  T_870;
  wire [63:0] T_878_0;
  reg [11:0] T_880;
  reg [31:0] GEN_5;
  wire [11:0] GEN_10;
  reg [63:0] T_889_0 [0:511];
  reg [63:0] GEN_6;
  wire [63:0] T_889_0_T_915_data;
  wire [8:0] T_889_0_T_915_addr;
  wire  T_889_0_T_915_en;
  reg [8:0] GEN_7;
  reg  GEN_9;
  wire [63:0] T_889_0_T_906_data;
  wire [8:0] T_889_0_T_906_addr;
  wire  T_889_0_T_906_mask;
  wire  T_889_0_T_906_en;
  wire  T_892;
  wire  T_894;
  wire [63:0] T_901_0;
  wire  GEN_18;
  wire [8:0] T_912;
  wire [63:0] T_923_0;
  wire  T_925;
  wire [63:0] T_933_0;
  reg [11:0] T_935;
  reg [31:0] GEN_11;
  wire [11:0] GEN_20;
  reg [63:0] T_944_0 [0:511];
  reg [63:0] GEN_12;
  wire [63:0] T_944_0_T_970_data;
  wire [8:0] T_944_0_T_970_addr;
  wire  T_944_0_T_970_en;
  reg [8:0] GEN_13;
  reg  GEN_14;
  wire [63:0] T_944_0_T_961_data;
  wire [8:0] T_944_0_T_961_addr;
  wire  T_944_0_T_961_mask;
  wire  T_944_0_T_961_en;
  wire  T_947;
  wire  T_949;
  wire [63:0] T_956_0;
  wire  GEN_28;
  wire [8:0] T_967;
  wire [63:0] T_978_0;
  wire  T_980;
  wire [63:0] T_988_0;
  reg [11:0] T_990;
  reg [31:0] GEN_15;
  wire [11:0] GEN_30;
  reg [63:0] T_999_0 [0:511];
  reg [63:0] GEN_16;
  wire [63:0] T_999_0_T_1025_data;
  wire [8:0] T_999_0_T_1025_addr;
  wire  T_999_0_T_1025_en;
  reg [8:0] GEN_17;
  reg  GEN_19;
  wire [63:0] T_999_0_T_1016_data;
  wire [8:0] T_999_0_T_1016_addr;
  wire  T_999_0_T_1016_mask;
  wire  T_999_0_T_1016_en;
  wire  T_1002;
  wire  T_1004;
  wire [63:0] T_1011_0;
  wire  GEN_38;
  wire [8:0] T_1022;
  wire [63:0] T_1033_0;
  assign io_read_ready = 1'h1;
  assign io_write_ready = 1'h1;
  assign io_resp_0 = T_868_0;
  assign io_resp_1 = T_923_0;
  assign io_resp_2 = T_978_0;
  assign io_resp_3 = T_1033_0;
  assign waddr = io_write_bits_addr[11:3];
  assign raddr = io_read_bits_addr[11:3];
  assign T_815 = io_write_bits_way_en[0];
  assign T_823_0 = T_834_0_T_860_data;
  assign GEN_0 = io_read_valid ? io_read_bits_addr : T_825;
  assign T_834_0_T_860_addr = T_857;
  assign T_834_0_T_860_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_834_0_T_860_data = T_834_0[GEN_3];
  `else
  assign T_834_0_T_860_data = GEN_3 >= 10'h200 ? $random : T_834_0[GEN_3];
  `endif
  assign T_834_0_T_851_data = T_846_0;
  assign T_834_0_T_851_addr = waddr;
  assign T_834_0_T_851_mask = GEN_8;
  assign T_834_0_T_851_en = T_839;
  assign T_837 = T_815 & io_write_valid;
  assign T_839 = T_837 & io_write_bits_wmask;
  assign T_846_0 = io_write_bits_data;
  assign GEN_8 = T_839 ? T_815 : 1'h0;
  assign T_857 = raddr;
  assign T_868_0 = T_823_0;
  assign T_870 = io_write_bits_way_en[1];
  assign T_878_0 = T_889_0_T_915_data;
  assign GEN_10 = io_read_valid ? io_read_bits_addr : T_880;
  assign T_889_0_T_915_addr = T_912;
  assign T_889_0_T_915_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_889_0_T_915_data = T_889_0[GEN_7];
  `else
  assign T_889_0_T_915_data = GEN_7 >= 10'h200 ? $random : T_889_0[GEN_7];
  `endif
  assign T_889_0_T_906_data = T_901_0;
  assign T_889_0_T_906_addr = waddr;
  assign T_889_0_T_906_mask = GEN_18;
  assign T_889_0_T_906_en = T_894;
  assign T_892 = T_870 & io_write_valid;
  assign T_894 = T_892 & io_write_bits_wmask;
  assign T_901_0 = io_write_bits_data;
  assign GEN_18 = T_894 ? T_870 : 1'h0;
  assign T_912 = raddr;
  assign T_923_0 = T_878_0;
  assign T_925 = io_write_bits_way_en[2];
  assign T_933_0 = T_944_0_T_970_data;
  assign GEN_20 = io_read_valid ? io_read_bits_addr : T_935;
  assign T_944_0_T_970_addr = T_967;
  assign T_944_0_T_970_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_944_0_T_970_data = T_944_0[GEN_13];
  `else
  assign T_944_0_T_970_data = GEN_13 >= 10'h200 ? $random : T_944_0[GEN_13];
  `endif
  assign T_944_0_T_961_data = T_956_0;
  assign T_944_0_T_961_addr = waddr;
  assign T_944_0_T_961_mask = GEN_28;
  assign T_944_0_T_961_en = T_949;
  assign T_947 = T_925 & io_write_valid;
  assign T_949 = T_947 & io_write_bits_wmask;
  assign T_956_0 = io_write_bits_data;
  assign GEN_28 = T_949 ? T_925 : 1'h0;
  assign T_967 = raddr;
  assign T_978_0 = T_933_0;
  assign T_980 = io_write_bits_way_en[3];
  assign T_988_0 = T_999_0_T_1025_data;
  assign GEN_30 = io_read_valid ? io_read_bits_addr : T_990;
  assign T_999_0_T_1025_addr = T_1022;
  assign T_999_0_T_1025_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_999_0_T_1025_data = T_999_0[GEN_17];
  `else
  assign T_999_0_T_1025_data = GEN_17 >= 10'h200 ? $random : T_999_0[GEN_17];
  `endif
  assign T_999_0_T_1016_data = T_1011_0;
  assign T_999_0_T_1016_addr = waddr;
  assign T_999_0_T_1016_mask = GEN_38;
  assign T_999_0_T_1016_en = T_1004;
  assign T_1002 = T_980 & io_write_valid;
  assign T_1004 = T_1002 & io_write_bits_wmask;
  assign T_1011_0 = io_write_bits_data;
  assign GEN_38 = T_1004 ? T_980 : 1'h0;
  assign T_1022 = raddr;
  assign T_1033_0 = T_988_0;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_1 = {1{$random}};
  T_825 = GEN_1[11:0];
  GEN_2 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_834_0[initvar] = GEN_2[63:0];
  GEN_5 = {1{$random}};
  T_880 = GEN_5[11:0];
  GEN_6 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_889_0[initvar] = GEN_6[63:0];
  GEN_11 = {1{$random}};
  T_935 = GEN_11[11:0];
  GEN_12 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_944_0[initvar] = GEN_12[63:0];
  GEN_15 = {1{$random}};
  T_990 = GEN_15[11:0];
  GEN_16 = {2{$random}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    T_999_0[initvar] = GEN_16[63:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      T_825 <= GEN_0;
    end
    GEN_3 <= T_834_0_T_860_addr;
    GEN_4 <= T_834_0_T_860_en;
    if(T_834_0_T_851_en & T_834_0_T_851_mask) begin
      T_834_0[T_834_0_T_851_addr] <= T_834_0_T_851_data;
    end
    if(1'h0) begin
    end else begin
      T_880 <= GEN_10;
    end
    GEN_7 <= T_889_0_T_915_addr;
    GEN_9 <= T_889_0_T_915_en;
    if(T_889_0_T_906_en & T_889_0_T_906_mask) begin
      T_889_0[T_889_0_T_906_addr] <= T_889_0_T_906_data;
    end
    if(1'h0) begin
    end else begin
      T_935 <= GEN_20;
    end
    GEN_13 <= T_944_0_T_970_addr;
    GEN_14 <= T_944_0_T_970_en;
    if(T_944_0_T_961_en & T_944_0_T_961_mask) begin
      T_944_0[T_944_0_T_961_addr] <= T_944_0_T_961_data;
    end
    if(1'h0) begin
    end else begin
      T_990 <= GEN_30;
    end
    GEN_17 <= T_999_0_T_1025_addr;
    GEN_19 <= T_999_0_T_1025_en;
    if(T_999_0_T_1016_en & T_999_0_T_1016_mask) begin
      T_999_0[T_999_0_T_1016_addr] <= T_999_0_T_1016_data;
    end
  end
endmodule
module Arbiter_85(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  output  io_in_2_ready,
  input   io_in_2_valid,
  input  [3:0] io_in_2_bits_way_en,
  input  [11:0] io_in_2_bits_addr,
  output  io_in_3_ready,
  input   io_in_3_valid,
  input  [3:0] io_in_3_bits_way_en,
  input  [11:0] io_in_3_bits_addr,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output [1:0] io_chosen
);
  wire [1:0] GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire [1:0] GEN_3;
  wire [3:0] GEN_4;
  wire [11:0] GEN_5;
  wire [1:0] GEN_6;
  wire [3:0] GEN_7;
  wire [11:0] GEN_8;
  wire  T_2205;
  wire  T_2206;
  wire  T_2208;
  wire  T_2210;
  wire  T_2212;
  wire  T_2214;
  wire  T_2215;
  wire  T_2216;
  wire  T_2218;
  wire  T_2219;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_2214;
  assign io_in_2_ready = T_2215;
  assign io_in_3_ready = T_2216;
  assign io_out_valid = T_2219;
  assign io_out_bits_way_en = GEN_7;
  assign io_out_bits_addr = GEN_8;
  assign io_chosen = GEN_6;
  assign GEN_0 = io_in_2_valid ? 2'h2 : 2'h3;
  assign GEN_1 = io_in_2_valid ? io_in_2_bits_way_en : io_in_3_bits_way_en;
  assign GEN_2 = io_in_2_valid ? io_in_2_bits_addr : io_in_3_bits_addr;
  assign GEN_3 = io_in_1_valid ? {{1'd0}, 1'h1} : GEN_0;
  assign GEN_4 = io_in_1_valid ? io_in_1_bits_way_en : GEN_1;
  assign GEN_5 = io_in_1_valid ? io_in_1_bits_addr : GEN_2;
  assign GEN_6 = io_in_0_valid ? {{1'd0}, 1'h0} : GEN_3;
  assign GEN_7 = io_in_0_valid ? io_in_0_bits_way_en : GEN_4;
  assign GEN_8 = io_in_0_valid ? io_in_0_bits_addr : GEN_5;
  assign T_2205 = io_in_0_valid | io_in_1_valid;
  assign T_2206 = T_2205 | io_in_2_valid;
  assign T_2208 = io_in_0_valid == 1'h0;
  assign T_2210 = T_2205 == 1'h0;
  assign T_2212 = T_2206 == 1'h0;
  assign T_2214 = T_2208 & io_out_ready;
  assign T_2215 = T_2210 & io_out_ready;
  assign T_2216 = T_2212 & io_out_ready;
  assign T_2218 = T_2212 == 1'h0;
  assign T_2219 = T_2218 | io_in_3_valid;
endmodule
module Arbiter_86(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [3:0] io_in_0_bits_way_en,
  input  [11:0] io_in_0_bits_addr,
  input   io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [3:0] io_in_1_bits_way_en,
  input  [11:0] io_in_1_bits_addr,
  input   io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [3:0] io_out_bits_way_en,
  output [11:0] io_out_bits_addr,
  output  io_out_bits_wmask,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  GEN_0;
  wire [3:0] GEN_1;
  wire [11:0] GEN_2;
  wire  GEN_3;
  wire [63:0] GEN_4;
  wire  T_1664;
  wire  T_1666;
  wire  T_1668;
  wire  T_1669;
  assign io_in_0_ready = io_out_ready;
  assign io_in_1_ready = T_1666;
  assign io_out_valid = T_1669;
  assign io_out_bits_way_en = GEN_1;
  assign io_out_bits_addr = GEN_2;
  assign io_out_bits_wmask = GEN_3;
  assign io_out_bits_data = GEN_4;
  assign io_chosen = GEN_0;
  assign GEN_0 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_1 = io_in_0_valid ? io_in_0_bits_way_en : io_in_1_bits_way_en;
  assign GEN_2 = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr;
  assign GEN_3 = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask;
  assign GEN_4 = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data;
  assign T_1664 = io_in_0_valid == 1'h0;
  assign T_1666 = T_1664 & io_out_ready;
  assign T_1668 = T_1664 == 1'h0;
  assign T_1669 = T_1668 | io_in_1_valid;
endmodule
module AMOALU(
  input   clk,
  input   reset,
  input  [5:0] io_addr,
  input  [4:0] io_cmd,
  input  [2:0] io_typ,
  input  [63:0] io_lhs,
  input  [63:0] io_rhs,
  output [63:0] io_out
);
  wire [1:0] T_6;
  wire  T_8;
  wire [31:0] T_9;
  wire [63:0] T_10;
  wire [63:0] rhs;
  wire  T_11;
  wire  T_12;
  wire  sgned;
  wire  T_14;
  wire  max;
  wire  T_16;
  wire  min;
  wire  T_17;
  wire  T_18;
  wire  T_19;
  wire  T_20;
  wire  T_21;
  wire  T_22;
  wire  word;
  wire  T_25;
  wire [31:0] GEN_0;
  wire [31:0] T_26;
  wire [63:0] GEN_1;
  wire [63:0] T_27;
  wire [63:0] T_28;
  wire [63:0] T_29;
  wire [64:0] T_30;
  wire [63:0] adder_out;
  wire  T_33;
  wire  T_34;
  wire  T_35;
  wire  T_36;
  wire  T_37;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire [31:0] T_45;
  wire [31:0] T_46;
  wire  T_47;
  wire [31:0] T_48;
  wire [31:0] T_49;
  wire  T_50;
  wire  T_53;
  wire  T_55;
  wire  T_56;
  wire  T_57;
  wire  T_58;
  wire  T_59;
  wire  T_60;
  wire  less;
  wire  T_61;
  wire  T_62;
  wire [63:0] T_63;
  wire  T_64;
  wire [63:0] T_65;
  wire  T_66;
  wire [63:0] T_67;
  wire  T_68;
  wire [1:0] GEN_2;
  wire  T_70;
  wire [7:0] T_71;
  wire [15:0] T_72;
  wire [31:0] T_73;
  wire [63:0] T_74;
  wire [1:0] GEN_3;
  wire  T_76;
  wire [15:0] T_77;
  wire [31:0] T_78;
  wire [63:0] T_79;
  wire [63:0] T_85;
  wire [63:0] T_86;
  wire [63:0] T_87;
  wire [63:0] T_88;
  wire [63:0] T_89;
  wire [63:0] T_90;
  wire [63:0] out;
  wire  T_92;
  wire  T_96;
  wire  T_100;
  wire  T_103;
  wire [1:0] T_104;
  wire  T_105;
  wire [1:0] T_107;
  wire  T_109;
  wire [1:0] T_112;
  wire [1:0] T_113;
  wire [1:0] T_116;
  wire [3:0] T_117;
  wire [3:0] T_120;
  wire  T_122;
  wire [3:0] T_125;
  wire [3:0] T_126;
  wire [3:0] T_129;
  wire [7:0] T_130;
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire  T_134;
  wire  T_135;
  wire  T_136;
  wire  T_137;
  wire  T_138;
  wire [7:0] GEN_5;
  wire [8:0] T_140;
  wire [7:0] T_141;
  wire [7:0] GEN_6;
  wire [8:0] T_143;
  wire [7:0] T_144;
  wire [7:0] GEN_7;
  wire [8:0] T_146;
  wire [7:0] T_147;
  wire [7:0] GEN_8;
  wire [8:0] T_149;
  wire [7:0] T_150;
  wire [7:0] GEN_9;
  wire [8:0] T_152;
  wire [7:0] T_153;
  wire [7:0] GEN_10;
  wire [8:0] T_155;
  wire [7:0] T_156;
  wire [7:0] GEN_11;
  wire [8:0] T_158;
  wire [7:0] T_159;
  wire [7:0] GEN_12;
  wire [8:0] T_161;
  wire [7:0] T_162;
  wire [7:0] T_168_0;
  wire [7:0] T_168_1;
  wire [7:0] T_168_2;
  wire [7:0] T_168_3;
  wire [7:0] T_168_4;
  wire [7:0] T_168_5;
  wire [7:0] T_168_6;
  wire [7:0] T_168_7;
  wire [15:0] T_170;
  wire [15:0] T_171;
  wire [31:0] T_172;
  wire [15:0] T_173;
  wire [15:0] T_174;
  wire [31:0] T_175;
  wire [63:0] wmask;
  wire [63:0] T_176;
  wire [63:0] T_177;
  wire [63:0] T_178;
  wire [63:0] T_179;
  assign io_out = T_179;
  assign T_6 = io_typ[1:0];
  assign T_8 = T_6 == 2'h2;
  assign T_9 = io_rhs[31:0];
  assign T_10 = {T_9,T_9};
  assign rhs = T_8 ? T_10 : io_rhs;
  assign T_11 = io_cmd == 5'hc;
  assign T_12 = io_cmd == 5'hd;
  assign sgned = T_11 | T_12;
  assign T_14 = io_cmd == 5'hf;
  assign max = T_12 | T_14;
  assign T_16 = io_cmd == 5'he;
  assign min = T_11 | T_16;
  assign T_17 = io_typ == 3'h2;
  assign T_18 = io_typ == 3'h6;
  assign T_19 = T_17 | T_18;
  assign T_20 = io_typ == 3'h0;
  assign T_21 = T_19 | T_20;
  assign T_22 = io_typ == 3'h4;
  assign word = T_21 | T_22;
  assign T_25 = io_addr[2];
  assign GEN_0 = {{31'd0}, T_25};
  assign T_26 = GEN_0 << 31;
  assign GEN_1 = {{32'd0}, T_26};
  assign T_27 = 64'hffffffffffffffff ^ GEN_1;
  assign T_28 = io_lhs & T_27;
  assign T_29 = rhs & T_27;
  assign T_30 = T_28 + T_29;
  assign adder_out = T_30[63:0];
  assign T_33 = T_25 == 1'h0;
  assign T_34 = word & T_33;
  assign T_35 = io_lhs[31];
  assign T_36 = io_lhs[63];
  assign T_37 = T_34 ? T_35 : T_36;
  assign T_42 = rhs[31];
  assign T_43 = rhs[63];
  assign T_44 = T_34 ? T_42 : T_43;
  assign T_45 = io_lhs[31:0];
  assign T_46 = rhs[31:0];
  assign T_47 = T_45 < T_46;
  assign T_48 = io_lhs[63:32];
  assign T_49 = rhs[63:32];
  assign T_50 = T_48 < T_49;
  assign T_53 = T_48 == T_49;
  assign T_55 = T_25 ? T_50 : T_47;
  assign T_56 = T_53 & T_47;
  assign T_57 = T_50 | T_56;
  assign T_58 = word ? T_55 : T_57;
  assign T_59 = T_37 == T_44;
  assign T_60 = sgned ? T_37 : T_44;
  assign less = T_59 ? T_58 : T_60;
  assign T_61 = io_cmd == 5'h8;
  assign T_62 = io_cmd == 5'hb;
  assign T_63 = io_lhs & rhs;
  assign T_64 = io_cmd == 5'ha;
  assign T_65 = io_lhs | rhs;
  assign T_66 = io_cmd == 5'h9;
  assign T_67 = io_lhs ^ rhs;
  assign T_68 = less ? min : max;
  assign GEN_2 = {{1'd0}, 1'h0};
  assign T_70 = T_6 == GEN_2;
  assign T_71 = io_rhs[7:0];
  assign T_72 = {T_71,T_71};
  assign T_73 = {T_72,T_72};
  assign T_74 = {T_73,T_73};
  assign GEN_3 = {{1'd0}, 1'h1};
  assign T_76 = T_6 == GEN_3;
  assign T_77 = io_rhs[15:0];
  assign T_78 = {T_77,T_77};
  assign T_79 = {T_78,T_78};
  assign T_85 = T_76 ? T_79 : rhs;
  assign T_86 = T_70 ? T_74 : T_85;
  assign T_87 = T_68 ? io_lhs : T_86;
  assign T_88 = T_66 ? T_67 : T_87;
  assign T_89 = T_64 ? T_65 : T_88;
  assign T_90 = T_62 ? T_63 : T_89;
  assign out = T_61 ? adder_out : T_90;
  assign T_92 = io_addr[0];
  assign T_96 = T_6 >= GEN_3;
  assign T_100 = T_92 | T_96;
  assign T_103 = T_92 ? 1'h0 : 1'h1;
  assign T_104 = {T_100,T_103};
  assign T_105 = io_addr[1];
  assign T_107 = T_105 ? T_104 : {{1'd0}, 1'h0};
  assign T_109 = T_6 >= 2'h2;
  assign T_112 = T_109 ? 2'h3 : {{1'd0}, 1'h0};
  assign T_113 = T_107 | T_112;
  assign T_116 = T_105 ? {{1'd0}, 1'h0} : T_104;
  assign T_117 = {T_113,T_116};
  assign T_120 = T_25 ? T_117 : {{3'd0}, 1'h0};
  assign T_122 = T_6 >= 2'h3;
  assign T_125 = T_122 ? 4'hf : {{3'd0}, 1'h0};
  assign T_126 = T_120 | T_125;
  assign T_129 = T_25 ? {{3'd0}, 1'h0} : T_117;
  assign T_130 = {T_126,T_129};
  assign T_131 = T_130[0];
  assign T_132 = T_130[1];
  assign T_133 = T_130[2];
  assign T_134 = T_130[3];
  assign T_135 = T_130[4];
  assign T_136 = T_130[5];
  assign T_137 = T_130[6];
  assign T_138 = T_130[7];
  assign GEN_5 = {{7'd0}, T_131};
  assign T_140 = 8'h0 - GEN_5;
  assign T_141 = T_140[7:0];
  assign GEN_6 = {{7'd0}, T_132};
  assign T_143 = 8'h0 - GEN_6;
  assign T_144 = T_143[7:0];
  assign GEN_7 = {{7'd0}, T_133};
  assign T_146 = 8'h0 - GEN_7;
  assign T_147 = T_146[7:0];
  assign GEN_8 = {{7'd0}, T_134};
  assign T_149 = 8'h0 - GEN_8;
  assign T_150 = T_149[7:0];
  assign GEN_9 = {{7'd0}, T_135};
  assign T_152 = 8'h0 - GEN_9;
  assign T_153 = T_152[7:0];
  assign GEN_10 = {{7'd0}, T_136};
  assign T_155 = 8'h0 - GEN_10;
  assign T_156 = T_155[7:0];
  assign GEN_11 = {{7'd0}, T_137};
  assign T_158 = 8'h0 - GEN_11;
  assign T_159 = T_158[7:0];
  assign GEN_12 = {{7'd0}, T_138};
  assign T_161 = 8'h0 - GEN_12;
  assign T_162 = T_161[7:0];
  assign T_168_0 = T_141;
  assign T_168_1 = T_144;
  assign T_168_2 = T_147;
  assign T_168_3 = T_150;
  assign T_168_4 = T_153;
  assign T_168_5 = T_156;
  assign T_168_6 = T_159;
  assign T_168_7 = T_162;
  assign T_170 = {T_168_1,T_168_0};
  assign T_171 = {T_168_3,T_168_2};
  assign T_172 = {T_171,T_170};
  assign T_173 = {T_168_5,T_168_4};
  assign T_174 = {T_168_7,T_168_6};
  assign T_175 = {T_174,T_173};
  assign wmask = {T_175,T_172};
  assign T_176 = wmask & out;
  assign T_177 = ~ wmask;
  assign T_178 = T_177 & io_lhs;
  assign T_179 = T_176 | T_178;
endmodule
module LockingArbiter_87(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [2:0] io_in_0_bits_addr_beat,
  input  [25:0] io_in_0_bits_addr_block,
  input  [1:0] io_in_0_bits_client_xact_id,
  input   io_in_0_bits_voluntary,
  input  [2:0] io_in_0_bits_r_type,
  input  [63:0] io_in_0_bits_data,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [2:0] io_in_1_bits_addr_beat,
  input  [25:0] io_in_1_bits_addr_block,
  input  [1:0] io_in_1_bits_client_xact_id,
  input   io_in_1_bits_voluntary,
  input  [2:0] io_in_1_bits_r_type,
  input  [63:0] io_in_1_bits_data,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [25:0] io_out_bits_addr_block,
  output [1:0] io_out_bits_client_xact_id,
  output  io_out_bits_voluntary,
  output [2:0] io_out_bits_r_type,
  output [63:0] io_out_bits_data,
  output  io_chosen
);
  wire  choice;
  wire  GEN_0;
  wire  GEN_7;
  wire [2:0] GEN_1;
  wire [2:0] GEN_8;
  wire [25:0] GEN_2;
  wire [25:0] GEN_9;
  wire [1:0] GEN_3;
  wire [1:0] GEN_10;
  wire  GEN_4;
  wire  GEN_11;
  wire [2:0] GEN_5;
  wire [2:0] GEN_12;
  wire [63:0] GEN_6;
  wire [63:0] GEN_13;
  reg [2:0] T_818;
  reg [31:0] GEN_20;
  reg  T_820;
  reg [31:0] GEN_21;
  wire [2:0] GEN_18;
  wire  T_822;
  wire [2:0] T_829_0;
  wire [2:0] T_829_1;
  wire [2:0] T_829_2;
  wire  T_831;
  wire  T_832;
  wire  T_833;
  wire  T_836;
  wire  T_837;
  wire  T_839;
  wire  T_840;
  wire [2:0] GEN_19;
  wire [3:0] T_844;
  wire [2:0] T_845;
  wire  GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire  T_848;
  wire  T_850;
  wire  T_851;
  wire  T_852;
  wire  T_855;
  wire  T_856;
  wire  GEN_17;
  assign io_in_0_ready = T_852;
  assign io_in_1_ready = T_856;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr_beat = GEN_1;
  assign io_out_bits_addr_block = GEN_2;
  assign io_out_bits_client_xact_id = GEN_3;
  assign io_out_bits_voluntary = GEN_4;
  assign io_out_bits_r_type = GEN_5;
  assign io_out_bits_data = GEN_6;
  assign io_chosen = GEN_16;
  assign choice = GEN_17;
  assign GEN_0 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_addr_beat : io_in_0_bits_addr_beat;
  assign GEN_2 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_addr_block : io_in_0_bits_addr_block;
  assign GEN_3 = GEN_10;
  assign GEN_10 = io_chosen ? io_in_1_bits_client_xact_id : io_in_0_bits_client_xact_id;
  assign GEN_4 = GEN_11;
  assign GEN_11 = io_chosen ? io_in_1_bits_voluntary : io_in_0_bits_voluntary;
  assign GEN_5 = GEN_12;
  assign GEN_12 = io_chosen ? io_in_1_bits_r_type : io_in_0_bits_r_type;
  assign GEN_6 = GEN_13;
  assign GEN_13 = io_chosen ? io_in_1_bits_data : io_in_0_bits_data;
  assign GEN_18 = {{2'd0}, 1'h0};
  assign T_822 = T_818 != GEN_18;
  assign T_829_0 = 3'h0;
  assign T_829_1 = 3'h1;
  assign T_829_2 = 3'h2;
  assign T_831 = T_829_0 == io_out_bits_r_type;
  assign T_832 = T_829_1 == io_out_bits_r_type;
  assign T_833 = T_829_2 == io_out_bits_r_type;
  assign T_836 = T_831 | T_832;
  assign T_837 = T_836 | T_833;
  assign T_839 = io_out_ready & io_out_valid;
  assign T_840 = T_839 & T_837;
  assign GEN_19 = {{2'd0}, 1'h1};
  assign T_844 = T_818 + GEN_19;
  assign T_845 = T_844[2:0];
  assign GEN_14 = T_840 ? io_chosen : T_820;
  assign GEN_15 = T_840 ? T_845 : T_818;
  assign GEN_16 = T_822 ? T_820 : choice;
  assign T_848 = io_in_0_valid == 1'h0;
  assign T_850 = T_820 == 1'h0;
  assign T_851 = T_822 ? T_850 : 1'h1;
  assign T_852 = T_851 & io_out_ready;
  assign T_855 = T_822 ? T_820 : T_848;
  assign T_856 = T_855 & io_out_ready;
  assign GEN_17 = io_in_0_valid ? 1'h0 : 1'h1;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  T_818 = GEN_20[2:0];
  GEN_21 = {1{$random}};
  T_820 = GEN_21[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_818 <= 3'h0;
    end else begin
      T_818 <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_820 <= GEN_14;
    end
  end
endmodule
module FlowThroughSerializer_88(
  input   clk,
  input   reset,
  output  io_in_ready,
  input   io_in_valid,
  input  [2:0] io_in_bits_addr_beat,
  input  [1:0] io_in_bits_client_xact_id,
  input  [2:0] io_in_bits_manager_xact_id,
  input   io_in_bits_is_builtin_type,
  input  [3:0] io_in_bits_g_type,
  input  [63:0] io_in_bits_data,
  input   io_in_bits_manager_id,
  input   io_out_ready,
  output  io_out_valid,
  output [2:0] io_out_bits_addr_beat,
  output [1:0] io_out_bits_client_xact_id,
  output [2:0] io_out_bits_manager_xact_id,
  output  io_out_bits_is_builtin_type,
  output [3:0] io_out_bits_g_type,
  output [63:0] io_out_bits_data,
  output  io_out_bits_manager_id,
  output  io_cnt,
  output  io_done
);
  assign io_in_ready = io_out_ready;
  assign io_out_valid = io_in_valid;
  assign io_out_bits_addr_beat = io_in_bits_addr_beat;
  assign io_out_bits_client_xact_id = io_in_bits_client_xact_id;
  assign io_out_bits_manager_xact_id = io_in_bits_manager_xact_id;
  assign io_out_bits_is_builtin_type = io_in_bits_is_builtin_type;
  assign io_out_bits_g_type = io_in_bits_g_type;
  assign io_out_bits_data = io_in_bits_data;
  assign io_out_bits_manager_id = io_in_bits_manager_id;
  assign io_cnt = 1'h0;
  assign io_done = 1'h1;
endmodule
module HellaCache(
  input   clk,
  input   reset,
  output  io_cpu_req_ready,
  input   io_cpu_req_valid,
  input  [39:0] io_cpu_req_bits_addr,
  input  [8:0] io_cpu_req_bits_tag,
  input  [4:0] io_cpu_req_bits_cmd,
  input  [2:0] io_cpu_req_bits_typ,
  input   io_cpu_req_bits_phys,
  input  [63:0] io_cpu_req_bits_data,
  input   io_cpu_s1_kill,
  input  [63:0] io_cpu_s1_data,
  output  io_cpu_s2_nack,
  output  io_cpu_resp_valid,
  output [39:0] io_cpu_resp_bits_addr,
  output [8:0] io_cpu_resp_bits_tag,
  output [4:0] io_cpu_resp_bits_cmd,
  output [2:0] io_cpu_resp_bits_typ,
  output [63:0] io_cpu_resp_bits_data,
  output  io_cpu_resp_bits_replay,
  output  io_cpu_resp_bits_has_data,
  output [63:0] io_cpu_resp_bits_data_word_bypass,
  output [63:0] io_cpu_resp_bits_store_data,
  output  io_cpu_replay_next,
  output  io_cpu_xcpt_ma_ld,
  output  io_cpu_xcpt_ma_st,
  output  io_cpu_xcpt_pf_ld,
  output  io_cpu_xcpt_pf_st,
  input   io_cpu_invalidate_lr,
  output  io_cpu_ordered,
  input   io_ptw_req_ready,
  output  io_ptw_req_valid,
  output [26:0] io_ptw_req_bits_addr,
  output [1:0] io_ptw_req_bits_prv,
  output  io_ptw_req_bits_store,
  output  io_ptw_req_bits_fetch,
  input   io_ptw_resp_valid,
  input  [19:0] io_ptw_resp_bits_pte_ppn,
  input  [2:0] io_ptw_resp_bits_pte_reserved_for_software,
  input   io_ptw_resp_bits_pte_d,
  input   io_ptw_resp_bits_pte_r,
  input  [3:0] io_ptw_resp_bits_pte_typ,
  input   io_ptw_resp_bits_pte_v,
  input   io_ptw_status_debug,
  input  [1:0] io_ptw_status_prv,
  input   io_ptw_status_sd,
  input  [30:0] io_ptw_status_zero3,
  input   io_ptw_status_sd_rv32,
  input  [1:0] io_ptw_status_zero2,
  input  [4:0] io_ptw_status_vm,
  input  [4:0] io_ptw_status_zero1,
  input   io_ptw_status_pum,
  input   io_ptw_status_mprv,
  input  [1:0] io_ptw_status_xs,
  input  [1:0] io_ptw_status_fs,
  input  [1:0] io_ptw_status_mpp,
  input  [1:0] io_ptw_status_hpp,
  input   io_ptw_status_spp,
  input   io_ptw_status_mpie,
  input   io_ptw_status_hpie,
  input   io_ptw_status_spie,
  input   io_ptw_status_upie,
  input   io_ptw_status_mie,
  input   io_ptw_status_hie,
  input   io_ptw_status_sie,
  input   io_ptw_status_uie,
  input   io_ptw_invalidate,
  input   io_mem_acquire_ready,
  output  io_mem_acquire_valid,
  output [25:0] io_mem_acquire_bits_addr_block,
  output [1:0] io_mem_acquire_bits_client_xact_id,
  output [2:0] io_mem_acquire_bits_addr_beat,
  output  io_mem_acquire_bits_is_builtin_type,
  output [2:0] io_mem_acquire_bits_a_type,
  output [11:0] io_mem_acquire_bits_union,
  output [63:0] io_mem_acquire_bits_data,
  output  io_mem_probe_ready,
  input   io_mem_probe_valid,
  input  [25:0] io_mem_probe_bits_addr_block,
  input  [1:0] io_mem_probe_bits_p_type,
  input   io_mem_release_ready,
  output  io_mem_release_valid,
  output [2:0] io_mem_release_bits_addr_beat,
  output [25:0] io_mem_release_bits_addr_block,
  output [1:0] io_mem_release_bits_client_xact_id,
  output  io_mem_release_bits_voluntary,
  output [2:0] io_mem_release_bits_r_type,
  output [63:0] io_mem_release_bits_data,
  output  io_mem_grant_ready,
  input   io_mem_grant_valid,
  input  [2:0] io_mem_grant_bits_addr_beat,
  input  [1:0] io_mem_grant_bits_client_xact_id,
  input  [2:0] io_mem_grant_bits_manager_xact_id,
  input   io_mem_grant_bits_is_builtin_type,
  input  [3:0] io_mem_grant_bits_g_type,
  input  [63:0] io_mem_grant_bits_data,
  input   io_mem_grant_bits_manager_id,
  input   io_mem_finish_ready,
  output  io_mem_finish_valid,
  output [2:0] io_mem_finish_bits_manager_xact_id,
  output  io_mem_finish_bits_manager_id
);
  wire  wb_clk;
  wire  wb_reset;
  wire  wb_io_req_ready;
  wire  wb_io_req_valid;
  wire [2:0] wb_io_req_bits_addr_beat;
  wire [25:0] wb_io_req_bits_addr_block;
  wire [1:0] wb_io_req_bits_client_xact_id;
  wire  wb_io_req_bits_voluntary;
  wire [2:0] wb_io_req_bits_r_type;
  wire [63:0] wb_io_req_bits_data;
  wire [3:0] wb_io_req_bits_way_en;
  wire  wb_io_meta_read_ready;
  wire  wb_io_meta_read_valid;
  wire [5:0] wb_io_meta_read_bits_idx;
  wire [3:0] wb_io_meta_read_bits_way_en;
  wire [19:0] wb_io_meta_read_bits_tag;
  wire  wb_io_data_req_ready;
  wire  wb_io_data_req_valid;
  wire [3:0] wb_io_data_req_bits_way_en;
  wire [11:0] wb_io_data_req_bits_addr;
  wire [63:0] wb_io_data_resp;
  wire  wb_io_release_ready;
  wire  wb_io_release_valid;
  wire [2:0] wb_io_release_bits_addr_beat;
  wire [25:0] wb_io_release_bits_addr_block;
  wire [1:0] wb_io_release_bits_client_xact_id;
  wire  wb_io_release_bits_voluntary;
  wire [2:0] wb_io_release_bits_r_type;
  wire [63:0] wb_io_release_bits_data;
  wire  prober_clk;
  wire  prober_reset;
  wire  prober_io_req_ready;
  wire  prober_io_req_valid;
  wire [25:0] prober_io_req_bits_addr_block;
  wire [1:0] prober_io_req_bits_p_type;
  wire [1:0] prober_io_req_bits_client_xact_id;
  wire  prober_io_rep_ready;
  wire  prober_io_rep_valid;
  wire [2:0] prober_io_rep_bits_addr_beat;
  wire [25:0] prober_io_rep_bits_addr_block;
  wire [1:0] prober_io_rep_bits_client_xact_id;
  wire  prober_io_rep_bits_voluntary;
  wire [2:0] prober_io_rep_bits_r_type;
  wire [63:0] prober_io_rep_bits_data;
  wire  prober_io_meta_read_ready;
  wire  prober_io_meta_read_valid;
  wire [5:0] prober_io_meta_read_bits_idx;
  wire [3:0] prober_io_meta_read_bits_way_en;
  wire [19:0] prober_io_meta_read_bits_tag;
  wire  prober_io_meta_write_ready;
  wire  prober_io_meta_write_valid;
  wire [5:0] prober_io_meta_write_bits_idx;
  wire [3:0] prober_io_meta_write_bits_way_en;
  wire [19:0] prober_io_meta_write_bits_data_tag;
  wire [1:0] prober_io_meta_write_bits_data_coh_state;
  wire  prober_io_wb_req_ready;
  wire  prober_io_wb_req_valid;
  wire [2:0] prober_io_wb_req_bits_addr_beat;
  wire [25:0] prober_io_wb_req_bits_addr_block;
  wire [1:0] prober_io_wb_req_bits_client_xact_id;
  wire  prober_io_wb_req_bits_voluntary;
  wire [2:0] prober_io_wb_req_bits_r_type;
  wire [63:0] prober_io_wb_req_bits_data;
  wire [3:0] prober_io_wb_req_bits_way_en;
  wire [3:0] prober_io_way_en;
  wire  prober_io_mshr_rdy;
  wire [1:0] prober_io_block_state_state;
  wire  mshrs_clk;
  wire  mshrs_reset;
  wire  mshrs_io_req_ready;
  wire  mshrs_io_req_valid;
  wire [39:0] mshrs_io_req_bits_addr;
  wire [8:0] mshrs_io_req_bits_tag;
  wire [4:0] mshrs_io_req_bits_cmd;
  wire [2:0] mshrs_io_req_bits_typ;
  wire  mshrs_io_req_bits_phys;
  wire [63:0] mshrs_io_req_bits_data;
  wire  mshrs_io_req_bits_tag_match;
  wire [19:0] mshrs_io_req_bits_old_meta_tag;
  wire [1:0] mshrs_io_req_bits_old_meta_coh_state;
  wire [3:0] mshrs_io_req_bits_way_en;
  wire  mshrs_io_resp_ready;
  wire  mshrs_io_resp_valid;
  wire [39:0] mshrs_io_resp_bits_addr;
  wire [8:0] mshrs_io_resp_bits_tag;
  wire [4:0] mshrs_io_resp_bits_cmd;
  wire [2:0] mshrs_io_resp_bits_typ;
  wire [63:0] mshrs_io_resp_bits_data;
  wire  mshrs_io_resp_bits_replay;
  wire  mshrs_io_resp_bits_has_data;
  wire [63:0] mshrs_io_resp_bits_data_word_bypass;
  wire [63:0] mshrs_io_resp_bits_store_data;
  wire  mshrs_io_secondary_miss;
  wire  mshrs_io_mem_req_ready;
  wire  mshrs_io_mem_req_valid;
  wire [25:0] mshrs_io_mem_req_bits_addr_block;
  wire [1:0] mshrs_io_mem_req_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_req_bits_addr_beat;
  wire  mshrs_io_mem_req_bits_is_builtin_type;
  wire [2:0] mshrs_io_mem_req_bits_a_type;
  wire [11:0] mshrs_io_mem_req_bits_union;
  wire [63:0] mshrs_io_mem_req_bits_data;
  wire [3:0] mshrs_io_refill_way_en;
  wire [11:0] mshrs_io_refill_addr;
  wire  mshrs_io_meta_read_ready;
  wire  mshrs_io_meta_read_valid;
  wire [5:0] mshrs_io_meta_read_bits_idx;
  wire [3:0] mshrs_io_meta_read_bits_way_en;
  wire [19:0] mshrs_io_meta_read_bits_tag;
  wire  mshrs_io_meta_write_ready;
  wire  mshrs_io_meta_write_valid;
  wire [5:0] mshrs_io_meta_write_bits_idx;
  wire [3:0] mshrs_io_meta_write_bits_way_en;
  wire [19:0] mshrs_io_meta_write_bits_data_tag;
  wire [1:0] mshrs_io_meta_write_bits_data_coh_state;
  wire  mshrs_io_replay_ready;
  wire  mshrs_io_replay_valid;
  wire [39:0] mshrs_io_replay_bits_addr;
  wire [8:0] mshrs_io_replay_bits_tag;
  wire [4:0] mshrs_io_replay_bits_cmd;
  wire [2:0] mshrs_io_replay_bits_typ;
  wire  mshrs_io_replay_bits_phys;
  wire [63:0] mshrs_io_replay_bits_data;
  wire  mshrs_io_mem_grant_valid;
  wire [2:0] mshrs_io_mem_grant_bits_addr_beat;
  wire [1:0] mshrs_io_mem_grant_bits_client_xact_id;
  wire [2:0] mshrs_io_mem_grant_bits_manager_xact_id;
  wire  mshrs_io_mem_grant_bits_is_builtin_type;
  wire [3:0] mshrs_io_mem_grant_bits_g_type;
  wire [63:0] mshrs_io_mem_grant_bits_data;
  wire  mshrs_io_mem_grant_bits_manager_id;
  wire  mshrs_io_mem_finish_ready;
  wire  mshrs_io_mem_finish_valid;
  wire [2:0] mshrs_io_mem_finish_bits_manager_xact_id;
  wire  mshrs_io_mem_finish_bits_manager_id;
  wire  mshrs_io_wb_req_ready;
  wire  mshrs_io_wb_req_valid;
  wire [2:0] mshrs_io_wb_req_bits_addr_beat;
  wire [25:0] mshrs_io_wb_req_bits_addr_block;
  wire [1:0] mshrs_io_wb_req_bits_client_xact_id;
  wire  mshrs_io_wb_req_bits_voluntary;
  wire [2:0] mshrs_io_wb_req_bits_r_type;
  wire [63:0] mshrs_io_wb_req_bits_data;
  wire [3:0] mshrs_io_wb_req_bits_way_en;
  wire  mshrs_io_probe_rdy;
  wire  mshrs_io_fence_rdy;
  wire  mshrs_io_replay_next;
  wire  T_2075;
  reg  s1_valid;
  reg [31:0] GEN_94;
  reg [39:0] s1_req_addr;
  reg [63:0] GEN_104;
  reg [8:0] s1_req_tag;
  reg [31:0] GEN_105;
  reg [4:0] s1_req_cmd;
  reg [31:0] GEN_109;
  reg [2:0] s1_req_typ;
  reg [31:0] GEN_114;
  reg  s1_req_phys;
  reg [31:0] GEN_115;
  reg [63:0] s1_req_data;
  reg [63:0] GEN_116;
  wire  T_2153;
  wire  s1_valid_masked;
  reg  s1_replay;
  reg [31:0] GEN_117;
  reg  s1_clk_en;
  reg [31:0] GEN_118;
  reg  s2_valid;
  reg [31:0] GEN_119;
  reg [39:0] s2_req_addr;
  reg [63:0] GEN_120;
  reg [8:0] s2_req_tag;
  reg [31:0] GEN_121;
  reg [4:0] s2_req_cmd;
  reg [31:0] GEN_122;
  reg [2:0] s2_req_typ;
  reg [31:0] GEN_123;
  reg  s2_req_phys;
  reg [31:0] GEN_124;
  reg [63:0] s2_req_data;
  reg [63:0] GEN_125;
  reg  T_2233;
  reg [31:0] GEN_126;
  wire  T_2234;
  wire  s2_replay;
  wire  s2_recycle;
  wire  s2_valid_masked;
  reg  s3_valid;
  reg [31:0] GEN_127;
  reg [39:0] s3_req_addr;
  reg [63:0] GEN_128;
  reg [8:0] s3_req_tag;
  reg [31:0] GEN_129;
  reg [4:0] s3_req_cmd;
  reg [31:0] GEN_130;
  reg [2:0] s3_req_typ;
  reg [31:0] GEN_131;
  reg  s3_req_phys;
  reg [31:0] GEN_132;
  reg [63:0] s3_req_data;
  reg [63:0] GEN_133;
  reg [3:0] s3_way;
  reg [31:0] GEN_134;
  reg  s1_recycled;
  reg [31:0] GEN_135;
  wire  GEN_0;
  wire  T_2315;
  wire  T_2316;
  wire  T_2317;
  wire  T_2318;
  wire  T_2319;
  wire  T_2320;
  wire  T_2321;
  wire  T_2322;
  wire  s1_read;
  wire  T_2323;
  wire  T_2325;
  wire  s1_write;
  wire  T_2329;
  wire  T_2330;
  wire  T_2331;
  wire  T_2332;
  wire  s1_readwrite;
  wire  dtlb_clk;
  wire  dtlb_reset;
  wire  dtlb_io_req_ready;
  wire  dtlb_io_req_valid;
  wire [6:0] dtlb_io_req_bits_asid;
  wire [27:0] dtlb_io_req_bits_vpn;
  wire  dtlb_io_req_bits_passthrough;
  wire  dtlb_io_req_bits_instruction;
  wire  dtlb_io_req_bits_store;
  wire  dtlb_io_resp_miss;
  wire [19:0] dtlb_io_resp_ppn;
  wire  dtlb_io_resp_xcpt_ld;
  wire  dtlb_io_resp_xcpt_st;
  wire  dtlb_io_resp_xcpt_if;
  wire [7:0] dtlb_io_resp_hit_idx;
  wire  dtlb_io_ptw_req_ready;
  wire  dtlb_io_ptw_req_valid;
  wire [26:0] dtlb_io_ptw_req_bits_addr;
  wire [1:0] dtlb_io_ptw_req_bits_prv;
  wire  dtlb_io_ptw_req_bits_store;
  wire  dtlb_io_ptw_req_bits_fetch;
  wire  dtlb_io_ptw_resp_valid;
  wire [19:0] dtlb_io_ptw_resp_bits_pte_ppn;
  wire [2:0] dtlb_io_ptw_resp_bits_pte_reserved_for_software;
  wire  dtlb_io_ptw_resp_bits_pte_d;
  wire  dtlb_io_ptw_resp_bits_pte_r;
  wire [3:0] dtlb_io_ptw_resp_bits_pte_typ;
  wire  dtlb_io_ptw_resp_bits_pte_v;
  wire  dtlb_io_ptw_status_debug;
  wire [1:0] dtlb_io_ptw_status_prv;
  wire  dtlb_io_ptw_status_sd;
  wire [30:0] dtlb_io_ptw_status_zero3;
  wire  dtlb_io_ptw_status_sd_rv32;
  wire [1:0] dtlb_io_ptw_status_zero2;
  wire [4:0] dtlb_io_ptw_status_vm;
  wire [4:0] dtlb_io_ptw_status_zero1;
  wire  dtlb_io_ptw_status_pum;
  wire  dtlb_io_ptw_status_mprv;
  wire [1:0] dtlb_io_ptw_status_xs;
  wire [1:0] dtlb_io_ptw_status_fs;
  wire [1:0] dtlb_io_ptw_status_mpp;
  wire [1:0] dtlb_io_ptw_status_hpp;
  wire  dtlb_io_ptw_status_spp;
  wire  dtlb_io_ptw_status_mpie;
  wire  dtlb_io_ptw_status_hpie;
  wire  dtlb_io_ptw_status_spie;
  wire  dtlb_io_ptw_status_upie;
  wire  dtlb_io_ptw_status_mie;
  wire  dtlb_io_ptw_status_hie;
  wire  dtlb_io_ptw_status_sie;
  wire  dtlb_io_ptw_status_uie;
  wire  dtlb_io_ptw_invalidate;
  wire  T_2333;
  wire [27:0] T_2335;
  wire  T_2338;
  wire  T_2340;
  wire  T_2341;
  wire  GEN_1;
  wire [39:0] GEN_2;
  wire [8:0] GEN_3;
  wire [4:0] GEN_4;
  wire [2:0] GEN_5;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire [25:0] T_2343;
  wire [31:0] GEN_83;
  wire [31:0] T_2344;
  wire [39:0] GEN_8;
  wire  GEN_9;
  wire [25:0] T_2346;
  wire [31:0] GEN_84;
  wire [31:0] T_2347;
  wire [39:0] GEN_10;
  wire  GEN_11;
  wire [39:0] GEN_12;
  wire [8:0] GEN_13;
  wire [4:0] GEN_14;
  wire [2:0] GEN_15;
  wire  GEN_16;
  wire [63:0] GEN_17;
  wire [39:0] GEN_18;
  wire [8:0] GEN_19;
  wire [4:0] GEN_20;
  wire [2:0] GEN_21;
  wire  GEN_22;
  wire [63:0] GEN_23;
  wire [11:0] T_2349;
  wire [31:0] s1_addr;
  wire [63:0] T_2350;
  wire [63:0] GEN_24;
  wire [63:0] GEN_25;
  wire [2:0] GEN_26;
  wire  GEN_27;
  wire [39:0] GEN_28;
  wire [63:0] GEN_29;
  wire [8:0] GEN_30;
  wire [4:0] GEN_31;
  wire [1:0] T_2352;
  wire [3:0] GEN_85;
  wire [3:0] T_2354;
  wire [4:0] T_2356;
  wire [3:0] T_2357;
  wire [2:0] T_2358;
  wire [39:0] GEN_87;
  wire [39:0] T_2359;
  wire [39:0] GEN_88;
  wire  misaligned;
  wire  T_2361;
  wire  T_2362;
  wire  T_2363;
  wire  T_2364;
  wire  T_2365;
  wire  T_2366;
  wire  T_2367;
  reg  T_2368;
  reg [31:0] GEN_136;
  wire  T_2369;
  wire  T_2371;
  wire  T_2372;
  wire  T_2374;
  wire  meta_clk;
  wire  meta_reset;
  wire  meta_io_read_ready;
  wire  meta_io_read_valid;
  wire [5:0] meta_io_read_bits_idx;
  wire [3:0] meta_io_read_bits_way_en;
  wire  meta_io_write_ready;
  wire  meta_io_write_valid;
  wire [5:0] meta_io_write_bits_idx;
  wire [3:0] meta_io_write_bits_way_en;
  wire [19:0] meta_io_write_bits_data_tag;
  wire [1:0] meta_io_write_bits_data_coh_state;
  wire [19:0] meta_io_resp_0_tag;
  wire [1:0] meta_io_resp_0_coh_state;
  wire [19:0] meta_io_resp_1_tag;
  wire [1:0] meta_io_resp_1_coh_state;
  wire [19:0] meta_io_resp_2_tag;
  wire [1:0] meta_io_resp_2_coh_state;
  wire [19:0] meta_io_resp_3_tag;
  wire [1:0] meta_io_resp_3_coh_state;
  wire  metaReadArb_clk;
  wire  metaReadArb_reset;
  wire  metaReadArb_io_in_0_ready;
  wire  metaReadArb_io_in_0_valid;
  wire [5:0] metaReadArb_io_in_0_bits_idx;
  wire [3:0] metaReadArb_io_in_0_bits_way_en;
  wire  metaReadArb_io_in_1_ready;
  wire  metaReadArb_io_in_1_valid;
  wire [5:0] metaReadArb_io_in_1_bits_idx;
  wire [3:0] metaReadArb_io_in_1_bits_way_en;
  wire  metaReadArb_io_in_2_ready;
  wire  metaReadArb_io_in_2_valid;
  wire [5:0] metaReadArb_io_in_2_bits_idx;
  wire [3:0] metaReadArb_io_in_2_bits_way_en;
  wire  metaReadArb_io_in_3_ready;
  wire  metaReadArb_io_in_3_valid;
  wire [5:0] metaReadArb_io_in_3_bits_idx;
  wire [3:0] metaReadArb_io_in_3_bits_way_en;
  wire  metaReadArb_io_in_4_ready;
  wire  metaReadArb_io_in_4_valid;
  wire [5:0] metaReadArb_io_in_4_bits_idx;
  wire [3:0] metaReadArb_io_in_4_bits_way_en;
  wire  metaReadArb_io_out_ready;
  wire  metaReadArb_io_out_valid;
  wire [5:0] metaReadArb_io_out_bits_idx;
  wire [3:0] metaReadArb_io_out_bits_way_en;
  wire [2:0] metaReadArb_io_chosen;
  wire  metaWriteArb_clk;
  wire  metaWriteArb_reset;
  wire  metaWriteArb_io_in_0_ready;
  wire  metaWriteArb_io_in_0_valid;
  wire [5:0] metaWriteArb_io_in_0_bits_idx;
  wire [3:0] metaWriteArb_io_in_0_bits_way_en;
  wire [19:0] metaWriteArb_io_in_0_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_0_bits_data_coh_state;
  wire  metaWriteArb_io_in_1_ready;
  wire  metaWriteArb_io_in_1_valid;
  wire [5:0] metaWriteArb_io_in_1_bits_idx;
  wire [3:0] metaWriteArb_io_in_1_bits_way_en;
  wire [19:0] metaWriteArb_io_in_1_bits_data_tag;
  wire [1:0] metaWriteArb_io_in_1_bits_data_coh_state;
  wire  metaWriteArb_io_out_ready;
  wire  metaWriteArb_io_out_valid;
  wire [5:0] metaWriteArb_io_out_bits_idx;
  wire [3:0] metaWriteArb_io_out_bits_way_en;
  wire [19:0] metaWriteArb_io_out_bits_data_tag;
  wire [1:0] metaWriteArb_io_out_bits_data_coh_state;
  wire  metaWriteArb_io_chosen;
  wire  data_clk;
  wire  data_reset;
  wire  data_io_read_ready;
  wire  data_io_read_valid;
  wire [3:0] data_io_read_bits_way_en;
  wire [11:0] data_io_read_bits_addr;
  wire  data_io_write_ready;
  wire  data_io_write_valid;
  wire [3:0] data_io_write_bits_way_en;
  wire [11:0] data_io_write_bits_addr;
  wire  data_io_write_bits_wmask;
  wire [63:0] data_io_write_bits_data;
  wire [63:0] data_io_resp_0;
  wire [63:0] data_io_resp_1;
  wire [63:0] data_io_resp_2;
  wire [63:0] data_io_resp_3;
  wire  readArb_clk;
  wire  readArb_reset;
  wire  readArb_io_in_0_ready;
  wire  readArb_io_in_0_valid;
  wire [3:0] readArb_io_in_0_bits_way_en;
  wire [11:0] readArb_io_in_0_bits_addr;
  wire  readArb_io_in_1_ready;
  wire  readArb_io_in_1_valid;
  wire [3:0] readArb_io_in_1_bits_way_en;
  wire [11:0] readArb_io_in_1_bits_addr;
  wire  readArb_io_in_2_ready;
  wire  readArb_io_in_2_valid;
  wire [3:0] readArb_io_in_2_bits_way_en;
  wire [11:0] readArb_io_in_2_bits_addr;
  wire  readArb_io_in_3_ready;
  wire  readArb_io_in_3_valid;
  wire [3:0] readArb_io_in_3_bits_way_en;
  wire [11:0] readArb_io_in_3_bits_addr;
  wire  readArb_io_out_ready;
  wire  readArb_io_out_valid;
  wire [3:0] readArb_io_out_bits_way_en;
  wire [11:0] readArb_io_out_bits_addr;
  wire [1:0] readArb_io_chosen;
  wire  writeArb_clk;
  wire  writeArb_reset;
  wire  writeArb_io_in_0_ready;
  wire  writeArb_io_in_0_valid;
  wire [3:0] writeArb_io_in_0_bits_way_en;
  wire [11:0] writeArb_io_in_0_bits_addr;
  wire  writeArb_io_in_0_bits_wmask;
  wire [63:0] writeArb_io_in_0_bits_data;
  wire  writeArb_io_in_1_ready;
  wire  writeArb_io_in_1_valid;
  wire [3:0] writeArb_io_in_1_bits_way_en;
  wire [11:0] writeArb_io_in_1_bits_addr;
  wire  writeArb_io_in_1_bits_wmask;
  wire [63:0] writeArb_io_in_1_bits_data;
  wire  writeArb_io_out_ready;
  wire  writeArb_io_out_valid;
  wire [3:0] writeArb_io_out_bits_way_en;
  wire [11:0] writeArb_io_out_bits_addr;
  wire  writeArb_io_out_bits_wmask;
  wire [63:0] writeArb_io_out_bits_data;
  wire  writeArb_io_chosen;
  wire [63:0] T_2765;
  wire [33:0] T_2766;
  wire  T_2768;
  wire  GEN_32;
  wire  T_2773;
  wire  GEN_33;
  wire [33:0] T_2775;
  wire [19:0] T_2778;
  wire  T_2779;
  wire  T_2781;
  wire  T_2783;
  wire  T_2785;
  wire  T_2791_0;
  wire  T_2791_1;
  wire  T_2791_2;
  wire  T_2791_3;
  wire [1:0] T_2793;
  wire [1:0] T_2794;
  wire [3:0] s1_tag_eq_way;
  wire  T_2795;
  wire  T_2796;
  wire  T_2797;
  wire  T_2798;
  wire  T_2799;
  wire  T_2800;
  wire  T_2801;
  wire  T_2802;
  wire  T_2803;
  wire  T_2804;
  wire  T_2805;
  wire  T_2806;
  wire  T_2812_0;
  wire  T_2812_1;
  wire  T_2812_2;
  wire  T_2812_3;
  wire [1:0] T_2814;
  wire [1:0] T_2815;
  wire [3:0] s1_tag_match_way;
  wire  T_2817;
  reg [3:0] s2_tag_match_way;
  reg [31:0] GEN_137;
  wire [3:0] GEN_34;
  wire [3:0] GEN_89;
  wire  s2_tag_match;
  reg [1:0] T_2822_state;
  reg [31:0] GEN_138;
  wire [1:0] GEN_35;
  reg [1:0] T_2847_state;
  reg [31:0] GEN_139;
  wire [1:0] GEN_36;
  reg [1:0] T_2872_state;
  reg [31:0] GEN_140;
  wire [1:0] GEN_37;
  reg [1:0] T_2897_state;
  reg [31:0] GEN_141;
  wire [1:0] GEN_38;
  wire [1:0] T_3119_0_state;
  wire [1:0] T_3119_1_state;
  wire [1:0] T_3119_2_state;
  wire [1:0] T_3119_3_state;
  wire  T_3241;
  wire  T_3242;
  wire  T_3243;
  wire  T_3244;
  wire [1:0] T_3246;
  wire [1:0] T_3248;
  wire [1:0] T_3250;
  wire [1:0] T_3252;
  wire [1:0] T_3278;
  wire [1:0] T_3279;
  wire [1:0] T_3280;
  wire [1:0] s2_hit_state_state;
  wire  T_3331;
  wire  T_3332;
  wire  T_3333;
  wire  T_3334;
  wire  T_3335;
  wire  T_3336;
  wire  T_3337;
  wire  T_3338;
  wire  T_3339;
  wire  T_3340;
  wire  T_3341;
  wire [1:0] T_3347_0;
  wire [1:0] T_3347_1;
  wire  T_3349;
  wire  T_3350;
  wire  T_3353;
  wire [1:0] T_3359_0;
  wire [1:0] T_3359_1;
  wire [1:0] T_3359_2;
  wire  T_3361;
  wire  T_3362;
  wire  T_3363;
  wire  T_3366;
  wire  T_3367;
  wire  T_3368;
  wire  T_3369;
  wire [1:0] T_3377;
  wire [1:0] T_3403_state;
  wire  T_3428;
  wire  s2_hit;
  reg [4:0] lrsc_count;
  reg [31:0] GEN_142;
  wire [4:0] GEN_90;
  wire  lrsc_valid;
  reg [33:0] lrsc_addr;
  reg [63:0] GEN_143;
  wire  T_3433;
  wire  s2_lrsc_addr_match;
  wire  T_3435;
  wire  s2_sc_fail;
  wire [4:0] GEN_91;
  wire [5:0] T_3437;
  wire [4:0] T_3438;
  wire [4:0] GEN_39;
  wire  T_3439;
  wire  T_3440;
  wire  T_3442;
  wire [4:0] GEN_40;
  wire [4:0] GEN_41;
  wire [33:0] GEN_42;
  wire [4:0] GEN_43;
  wire [4:0] GEN_44;
  wire [33:0] GEN_45;
  wire [4:0] GEN_46;
  wire [63:0] s2_data_0;
  wire [63:0] s2_data_1;
  wire [63:0] s2_data_2;
  wire [63:0] s2_data_3;
  reg [63:0] T_3460_0;
  reg [63:0] GEN_144;
  wire  T_3463;
  wire [63:0] T_3471;
  wire [63:0] GEN_47;
  reg [63:0] T_3478_0;
  reg [63:0] GEN_145;
  wire  T_3481;
  wire [63:0] T_3489;
  wire [63:0] GEN_48;
  reg [63:0] T_3496_0;
  reg [63:0] GEN_146;
  wire  T_3499;
  wire [63:0] T_3507;
  wire [63:0] GEN_49;
  reg [63:0] T_3514_0;
  reg [63:0] GEN_147;
  wire  T_3517;
  wire [63:0] T_3525;
  wire [63:0] GEN_50;
  wire [63:0] T_3531;
  wire [63:0] T_3533;
  wire [63:0] T_3535;
  wire [63:0] T_3537;
  wire [63:0] T_3539;
  wire [63:0] T_3540;
  wire [63:0] T_3541;
  wire [63:0] s2_data_muxed;
  wire [63:0] T_3548_0;
  wire [63:0] T_3555_0;
  wire  T_3563_0;
  wire  T_3565;
  wire  T_3569;
  wire  T_3570;
  wire  T_3578;
  wire  amoalu_clk;
  wire  amoalu_reset;
  wire [5:0] amoalu_io_addr;
  wire [4:0] amoalu_io_cmd;
  wire [2:0] amoalu_io_typ;
  wire [63:0] amoalu_io_lhs;
  wire [63:0] amoalu_io_rhs;
  wire [63:0] amoalu_io_out;
  wire  T_3579;
  wire  T_3587;
  wire  T_3588;
  wire [63:0] T_3589;
  wire [39:0] GEN_51;
  wire [8:0] GEN_52;
  wire [4:0] GEN_53;
  wire [2:0] GEN_54;
  wire  GEN_55;
  wire [63:0] GEN_56;
  wire [3:0] GEN_57;
  wire [1:0] GEN_92;
  wire [1:0] rowWMask;
  wire  T_3593;
  reg [15:0] T_3596;
  reg [31:0] GEN_148;
  wire  T_3597;
  wire  T_3598;
  wire  T_3599;
  wire  T_3600;
  wire  T_3601;
  wire  T_3602;
  wire  T_3603;
  wire [14:0] T_3604;
  wire [15:0] T_3605;
  wire [15:0] GEN_58;
  wire [1:0] T_3606;
  wire [3:0] s1_replaced_way_en;
  reg [1:0] T_3609;
  reg [31:0] GEN_149;
  wire [1:0] GEN_59;
  wire [3:0] s2_replaced_way_en;
  wire  T_3611;
  wire  T_3612;
  reg [19:0] T_3613_tag;
  reg [31:0] GEN_150;
  reg [1:0] T_3613_coh_state;
  reg [31:0] GEN_151;
  wire [19:0] GEN_60;
  wire [1:0] GEN_61;
  wire  T_3709;
  wire  T_3710;
  reg [19:0] T_3711_tag;
  reg [31:0] GEN_152;
  reg [1:0] T_3711_coh_state;
  reg [31:0] GEN_153;
  wire [19:0] GEN_62;
  wire [1:0] GEN_63;
  wire  T_3807;
  wire  T_3808;
  reg [19:0] T_3809_tag;
  reg [31:0] GEN_154;
  reg [1:0] T_3809_coh_state;
  reg [31:0] GEN_155;
  wire [19:0] GEN_64;
  wire [1:0] GEN_65;
  wire  T_3905;
  wire  T_3906;
  reg [19:0] T_3907_tag;
  reg [31:0] GEN_156;
  reg [1:0] T_3907_coh_state;
  reg [31:0] GEN_157;
  wire [19:0] GEN_66;
  wire [1:0] GEN_67;
  wire [19:0] T_4768_0_tag;
  wire [1:0] T_4768_0_coh_state;
  wire [19:0] T_4768_1_tag;
  wire [1:0] T_4768_1_coh_state;
  wire [19:0] T_4768_2_tag;
  wire [1:0] T_4768_2_coh_state;
  wire [19:0] T_4768_3_tag;
  wire [1:0] T_4768_3_coh_state;
  wire  T_5245;
  wire  T_5246;
  wire  T_5247;
  wire  T_5248;
  wire [21:0] T_5249;
  wire [21:0] T_5251;
  wire [21:0] T_5252;
  wire [21:0] T_5254;
  wire [21:0] T_5255;
  wire [21:0] T_5257;
  wire [21:0] T_5258;
  wire [21:0] T_5260;
  wire [21:0] T_5357;
  wire [21:0] T_5358;
  wire [21:0] T_5359;
  wire [19:0] s2_repl_meta_tag;
  wire [1:0] s2_repl_meta_coh_state;
  wire [1:0] T_5551;
  wire [19:0] T_5552;
  wire  T_5554;
  wire  T_5555;
  wire  T_5556;
  wire  T_5558;
  wire  T_5559;
  wire  T_5561;
  wire  T_5563;
  wire  T_5567;
  wire  T_5568;
  wire  T_5576;
  wire  T_5577;
  wire [19:0] T_5674_tag;
  wire [1:0] T_5674_coh_state;
  wire [19:0] T_5770_tag;
  wire [1:0] T_5770_coh_state;
  wire [3:0] T_5866;
  wire  T_5867;
  wire  T_5871;
  wire  releaseArb_clk;
  wire  releaseArb_reset;
  wire  releaseArb_io_in_0_ready;
  wire  releaseArb_io_in_0_valid;
  wire [2:0] releaseArb_io_in_0_bits_addr_beat;
  wire [25:0] releaseArb_io_in_0_bits_addr_block;
  wire [1:0] releaseArb_io_in_0_bits_client_xact_id;
  wire  releaseArb_io_in_0_bits_voluntary;
  wire [2:0] releaseArb_io_in_0_bits_r_type;
  wire [63:0] releaseArb_io_in_0_bits_data;
  wire  releaseArb_io_in_1_ready;
  wire  releaseArb_io_in_1_valid;
  wire [2:0] releaseArb_io_in_1_bits_addr_beat;
  wire [25:0] releaseArb_io_in_1_bits_addr_block;
  wire [1:0] releaseArb_io_in_1_bits_client_xact_id;
  wire  releaseArb_io_in_1_bits_voluntary;
  wire [2:0] releaseArb_io_in_1_bits_r_type;
  wire [63:0] releaseArb_io_in_1_bits_data;
  wire  releaseArb_io_out_ready;
  wire  releaseArb_io_out_valid;
  wire [2:0] releaseArb_io_out_bits_addr_beat;
  wire [25:0] releaseArb_io_out_bits_addr_block;
  wire [1:0] releaseArb_io_out_bits_client_xact_id;
  wire  releaseArb_io_out_bits_voluntary;
  wire [2:0] releaseArb_io_out_bits_r_type;
  wire [63:0] releaseArb_io_out_bits_data;
  wire  releaseArb_io_chosen;
  wire  T_5904;
  wire  T_5907;
  wire  FlowThroughSerializer_88_5908_clk;
  wire  FlowThroughSerializer_88_5908_reset;
  wire  FlowThroughSerializer_88_5908_io_in_ready;
  wire  FlowThroughSerializer_88_5908_io_in_valid;
  wire [2:0] FlowThroughSerializer_88_5908_io_in_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_88_5908_io_in_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_88_5908_io_in_bits_manager_xact_id;
  wire  FlowThroughSerializer_88_5908_io_in_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_88_5908_io_in_bits_g_type;
  wire [63:0] FlowThroughSerializer_88_5908_io_in_bits_data;
  wire  FlowThroughSerializer_88_5908_io_in_bits_manager_id;
  wire  FlowThroughSerializer_88_5908_io_out_ready;
  wire  FlowThroughSerializer_88_5908_io_out_valid;
  wire [2:0] FlowThroughSerializer_88_5908_io_out_bits_addr_beat;
  wire [1:0] FlowThroughSerializer_88_5908_io_out_bits_client_xact_id;
  wire [2:0] FlowThroughSerializer_88_5908_io_out_bits_manager_xact_id;
  wire  FlowThroughSerializer_88_5908_io_out_bits_is_builtin_type;
  wire [3:0] FlowThroughSerializer_88_5908_io_out_bits_g_type;
  wire [63:0] FlowThroughSerializer_88_5908_io_out_bits_data;
  wire  FlowThroughSerializer_88_5908_io_out_bits_manager_id;
  wire  FlowThroughSerializer_88_5908_io_cnt;
  wire  FlowThroughSerializer_88_5908_io_done;
  wire  T_5909;
  wire [2:0] T_5917_0;
  wire [2:0] T_5917_1;
  wire [3:0] GEN_95;
  wire  T_5919;
  wire [3:0] GEN_96;
  wire  T_5920;
  wire  T_5923;
  wire [1:0] T_5929_0;
  wire [1:0] T_5929_1;
  wire [3:0] GEN_97;
  wire  T_5931;
  wire [3:0] GEN_98;
  wire  T_5932;
  wire  T_5935;
  wire  T_5936;
  wire  T_5938;
  wire  T_5939;
  wire [2:0] T_5947_0;
  wire [2:0] T_5947_1;
  wire [3:0] GEN_99;
  wire  T_5949;
  wire [3:0] GEN_100;
  wire  T_5950;
  wire  T_5953;
  wire [1:0] T_5959_0;
  wire [1:0] T_5959_1;
  wire [3:0] GEN_101;
  wire  T_5961;
  wire [3:0] GEN_102;
  wire  T_5962;
  wire  T_5965;
  wire  T_5966;
  wire  T_5967;
  wire  T_5969;
  wire  T_5970;
  wire [63:0] T_5973;
  wire  T_5975;
  wire  T_5976;
  wire  wbArb_clk;
  wire  wbArb_reset;
  wire  wbArb_io_in_0_ready;
  wire  wbArb_io_in_0_valid;
  wire [2:0] wbArb_io_in_0_bits_addr_beat;
  wire [25:0] wbArb_io_in_0_bits_addr_block;
  wire [1:0] wbArb_io_in_0_bits_client_xact_id;
  wire  wbArb_io_in_0_bits_voluntary;
  wire [2:0] wbArb_io_in_0_bits_r_type;
  wire [63:0] wbArb_io_in_0_bits_data;
  wire [3:0] wbArb_io_in_0_bits_way_en;
  wire  wbArb_io_in_1_ready;
  wire  wbArb_io_in_1_valid;
  wire [2:0] wbArb_io_in_1_bits_addr_beat;
  wire [25:0] wbArb_io_in_1_bits_addr_block;
  wire [1:0] wbArb_io_in_1_bits_client_xact_id;
  wire  wbArb_io_in_1_bits_voluntary;
  wire [2:0] wbArb_io_in_1_bits_r_type;
  wire [63:0] wbArb_io_in_1_bits_data;
  wire [3:0] wbArb_io_in_1_bits_way_en;
  wire  wbArb_io_out_ready;
  wire  wbArb_io_out_valid;
  wire [2:0] wbArb_io_out_bits_addr_beat;
  wire [25:0] wbArb_io_out_bits_addr_block;
  wire [1:0] wbArb_io_out_bits_client_xact_id;
  wire  wbArb_io_out_bits_voluntary;
  wire [2:0] wbArb_io_out_bits_r_type;
  wire [63:0] wbArb_io_out_bits_data;
  wire [3:0] wbArb_io_out_bits_way_en;
  wire  wbArb_io_chosen;
  reg  s4_valid;
  reg [31:0] GEN_158;
  wire  T_6032;
  reg [39:0] s4_req_addr;
  reg [63:0] GEN_159;
  reg [8:0] s4_req_tag;
  reg [31:0] GEN_160;
  reg [4:0] s4_req_cmd;
  reg [31:0] GEN_161;
  reg [2:0] s4_req_typ;
  reg [31:0] GEN_162;
  reg  s4_req_phys;
  reg [31:0] GEN_163;
  reg [63:0] s4_req_data;
  reg [63:0] GEN_164;
  wire [39:0] GEN_69;
  wire [8:0] GEN_70;
  wire [4:0] GEN_71;
  wire [2:0] GEN_72;
  wire  GEN_73;
  wire [63:0] GEN_74;
  wire  T_6108;
  wire  T_6111;
  wire [28:0] T_6112;
  wire [36:0] T_6113;
  wire [36:0] GEN_103;
  wire  T_6114;
  wire  T_6115;
  wire  T_6123;
  wire [36:0] T_6125;
  wire  T_6126;
  wire  T_6127;
  wire  T_6128;
  wire  T_6129;
  wire  T_6130;
  wire  T_6131;
  wire  T_6132;
  wire  T_6133;
  wire  T_6134;
  wire  T_6135;
  wire [36:0] T_6137;
  wire  T_6138;
  wire  T_6139;
  wire  T_6140;
  wire  T_6141;
  wire  T_6142;
  wire  T_6143;
  wire  T_6144;
  wire  T_6145;
  wire  T_6146;
  wire  T_6147;
  reg [63:0] s2_store_bypass_data;
  reg [63:0] GEN_165;
  reg  s2_store_bypass;
  reg [31:0] GEN_166;
  wire  T_6151;
  wire  T_6152;
  wire [63:0] T_6153;
  wire [63:0] T_6154;
  wire [63:0] GEN_75;
  wire  GEN_77;
  wire [63:0] GEN_78;
  wire [63:0] s2_data_word_prebypass;
  wire [63:0] s2_data_word;
  wire [1:0] T_6158;
  wire [2:0] T_6159;
  wire  GEN_106;
  wire [2:0] GEN_107;
  wire  T_6161;
  wire  T_6162;
  wire [5:0] T_6163;
  wire  T_6164;
  wire  T_6166;
  wire  T_6167;
  wire  s1_nack;
  wire  T_6168;
  reg  s2_nack_hit;
  reg [31:0] GEN_167;
  wire  GEN_79;
  wire  GEN_80;
  wire  s2_nack_victim;
  wire  T_6173;
  wire  s2_nack_miss;
  wire  T_6174;
  wire  s2_nack;
  wire  T_6176;
  wire  T_6177;
  wire  T_6179;
  wire  s2_recycle_ecc;
  reg  s2_recycle_next;
  reg [31:0] GEN_168;
  wire  GEN_81;
  wire  T_6182;
  reg  block_miss;
  reg [31:0] GEN_169;
  wire  T_6184;
  wire  T_6185;
  wire  GEN_82;
  wire  cache_resp_valid;
  wire [39:0] cache_resp_bits_addr;
  wire [8:0] cache_resp_bits_tag;
  wire [4:0] cache_resp_bits_cmd;
  wire [2:0] cache_resp_bits_typ;
  wire [63:0] cache_resp_bits_data;
  wire  cache_resp_bits_replay;
  wire  cache_resp_bits_has_data;
  wire [63:0] cache_resp_bits_data_word_bypass;
  wire [63:0] cache_resp_bits_store_data;
  wire  T_6586;
  wire  T_6588;
  wire  T_6589;
  wire  T_6599;
  wire [31:0] T_6600;
  wire [31:0] T_6601;
  wire [31:0] T_6602;
  wire  T_6608;
  wire  T_6610;
  wire  T_6611;
  wire [31:0] GEN_108;
  wire [32:0] T_6613;
  wire [31:0] T_6614;
  wire [31:0] T_6616;
  wire [63:0] T_6617;
  wire  T_6618;
  wire [15:0] T_6619;
  wire [15:0] T_6620;
  wire [15:0] T_6621;
  wire  T_6627;
  wire  T_6629;
  wire  T_6630;
  wire [47:0] GEN_110;
  wire [48:0] T_6632;
  wire [47:0] T_6633;
  wire [47:0] T_6634;
  wire [47:0] T_6635;
  wire [63:0] T_6636;
  wire  T_6637;
  wire [7:0] T_6638;
  wire [7:0] T_6639;
  wire [7:0] T_6640;
  wire [7:0] T_6644;
  wire [1:0] GEN_111;
  wire  T_6646;
  wire  T_6647;
  wire  T_6648;
  wire  T_6649;
  wire [55:0] GEN_112;
  wire [56:0] T_6651;
  wire [55:0] T_6652;
  wire [55:0] T_6653;
  wire [55:0] T_6654;
  wire [63:0] T_6655;
  wire [63:0] GEN_113;
  wire [63:0] T_6656;
  wire  uncache_resp_valid;
  wire [39:0] uncache_resp_bits_addr;
  wire [8:0] uncache_resp_bits_tag;
  wire [4:0] uncache_resp_bits_cmd;
  wire [2:0] uncache_resp_bits_typ;
  wire [63:0] uncache_resp_bits_data;
  wire  uncache_resp_bits_replay;
  wire  uncache_resp_bits_has_data;
  wire [63:0] uncache_resp_bits_data_word_bypass;
  wire [63:0] uncache_resp_bits_store_data;
  wire  T_7057;
  reg  T_7058;
  reg [31:0] GEN_170;
  wire  T_7059;
  wire  T_7060_valid;
  wire [39:0] T_7060_bits_addr;
  wire [8:0] T_7060_bits_tag;
  wire [4:0] T_7060_bits_cmd;
  wire [2:0] T_7060_bits_typ;
  wire [63:0] T_7060_bits_data;
  wire  T_7060_bits_replay;
  wire  T_7060_bits_has_data;
  wire [63:0] T_7060_bits_store_data;
  wire  T_7241;
  wire  T_7243;
  wire  T_7244;
  wire  T_7245;
  wire  T_7246;
  reg [1:0] GEN_68;
  reg [31:0] GEN_171;
  reg [3:0] GEN_76;
  reg [31:0] GEN_172;
  reg [3:0] GEN_86;
  reg [31:0] GEN_173;
  reg [63:0] GEN_93;
  reg [63:0] GEN_174;
  WritebackUnit wb (
    .clk(wb_clk),
    .reset(wb_reset),
    .io_req_ready(wb_io_req_ready),
    .io_req_valid(wb_io_req_valid),
    .io_req_bits_addr_beat(wb_io_req_bits_addr_beat),
    .io_req_bits_addr_block(wb_io_req_bits_addr_block),
    .io_req_bits_client_xact_id(wb_io_req_bits_client_xact_id),
    .io_req_bits_voluntary(wb_io_req_bits_voluntary),
    .io_req_bits_r_type(wb_io_req_bits_r_type),
    .io_req_bits_data(wb_io_req_bits_data),
    .io_req_bits_way_en(wb_io_req_bits_way_en),
    .io_meta_read_ready(wb_io_meta_read_ready),
    .io_meta_read_valid(wb_io_meta_read_valid),
    .io_meta_read_bits_idx(wb_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(wb_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(wb_io_meta_read_bits_tag),
    .io_data_req_ready(wb_io_data_req_ready),
    .io_data_req_valid(wb_io_data_req_valid),
    .io_data_req_bits_way_en(wb_io_data_req_bits_way_en),
    .io_data_req_bits_addr(wb_io_data_req_bits_addr),
    .io_data_resp(wb_io_data_resp),
    .io_release_ready(wb_io_release_ready),
    .io_release_valid(wb_io_release_valid),
    .io_release_bits_addr_beat(wb_io_release_bits_addr_beat),
    .io_release_bits_addr_block(wb_io_release_bits_addr_block),
    .io_release_bits_client_xact_id(wb_io_release_bits_client_xact_id),
    .io_release_bits_voluntary(wb_io_release_bits_voluntary),
    .io_release_bits_r_type(wb_io_release_bits_r_type),
    .io_release_bits_data(wb_io_release_bits_data)
  );
  ProbeUnit prober (
    .clk(prober_clk),
    .reset(prober_reset),
    .io_req_ready(prober_io_req_ready),
    .io_req_valid(prober_io_req_valid),
    .io_req_bits_addr_block(prober_io_req_bits_addr_block),
    .io_req_bits_p_type(prober_io_req_bits_p_type),
    .io_req_bits_client_xact_id(prober_io_req_bits_client_xact_id),
    .io_rep_ready(prober_io_rep_ready),
    .io_rep_valid(prober_io_rep_valid),
    .io_rep_bits_addr_beat(prober_io_rep_bits_addr_beat),
    .io_rep_bits_addr_block(prober_io_rep_bits_addr_block),
    .io_rep_bits_client_xact_id(prober_io_rep_bits_client_xact_id),
    .io_rep_bits_voluntary(prober_io_rep_bits_voluntary),
    .io_rep_bits_r_type(prober_io_rep_bits_r_type),
    .io_rep_bits_data(prober_io_rep_bits_data),
    .io_meta_read_ready(prober_io_meta_read_ready),
    .io_meta_read_valid(prober_io_meta_read_valid),
    .io_meta_read_bits_idx(prober_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(prober_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(prober_io_meta_read_bits_tag),
    .io_meta_write_ready(prober_io_meta_write_ready),
    .io_meta_write_valid(prober_io_meta_write_valid),
    .io_meta_write_bits_idx(prober_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(prober_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(prober_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(prober_io_meta_write_bits_data_coh_state),
    .io_wb_req_ready(prober_io_wb_req_ready),
    .io_wb_req_valid(prober_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(prober_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(prober_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(prober_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(prober_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(prober_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(prober_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(prober_io_wb_req_bits_way_en),
    .io_way_en(prober_io_way_en),
    .io_mshr_rdy(prober_io_mshr_rdy),
    .io_block_state_state(prober_io_block_state_state)
  );
  MSHRFile mshrs (
    .clk(mshrs_clk),
    .reset(mshrs_reset),
    .io_req_ready(mshrs_io_req_ready),
    .io_req_valid(mshrs_io_req_valid),
    .io_req_bits_addr(mshrs_io_req_bits_addr),
    .io_req_bits_tag(mshrs_io_req_bits_tag),
    .io_req_bits_cmd(mshrs_io_req_bits_cmd),
    .io_req_bits_typ(mshrs_io_req_bits_typ),
    .io_req_bits_phys(mshrs_io_req_bits_phys),
    .io_req_bits_data(mshrs_io_req_bits_data),
    .io_req_bits_tag_match(mshrs_io_req_bits_tag_match),
    .io_req_bits_old_meta_tag(mshrs_io_req_bits_old_meta_tag),
    .io_req_bits_old_meta_coh_state(mshrs_io_req_bits_old_meta_coh_state),
    .io_req_bits_way_en(mshrs_io_req_bits_way_en),
    .io_resp_ready(mshrs_io_resp_ready),
    .io_resp_valid(mshrs_io_resp_valid),
    .io_resp_bits_addr(mshrs_io_resp_bits_addr),
    .io_resp_bits_tag(mshrs_io_resp_bits_tag),
    .io_resp_bits_cmd(mshrs_io_resp_bits_cmd),
    .io_resp_bits_typ(mshrs_io_resp_bits_typ),
    .io_resp_bits_data(mshrs_io_resp_bits_data),
    .io_resp_bits_replay(mshrs_io_resp_bits_replay),
    .io_resp_bits_has_data(mshrs_io_resp_bits_has_data),
    .io_resp_bits_data_word_bypass(mshrs_io_resp_bits_data_word_bypass),
    .io_resp_bits_store_data(mshrs_io_resp_bits_store_data),
    .io_secondary_miss(mshrs_io_secondary_miss),
    .io_mem_req_ready(mshrs_io_mem_req_ready),
    .io_mem_req_valid(mshrs_io_mem_req_valid),
    .io_mem_req_bits_addr_block(mshrs_io_mem_req_bits_addr_block),
    .io_mem_req_bits_client_xact_id(mshrs_io_mem_req_bits_client_xact_id),
    .io_mem_req_bits_addr_beat(mshrs_io_mem_req_bits_addr_beat),
    .io_mem_req_bits_is_builtin_type(mshrs_io_mem_req_bits_is_builtin_type),
    .io_mem_req_bits_a_type(mshrs_io_mem_req_bits_a_type),
    .io_mem_req_bits_union(mshrs_io_mem_req_bits_union),
    .io_mem_req_bits_data(mshrs_io_mem_req_bits_data),
    .io_refill_way_en(mshrs_io_refill_way_en),
    .io_refill_addr(mshrs_io_refill_addr),
    .io_meta_read_ready(mshrs_io_meta_read_ready),
    .io_meta_read_valid(mshrs_io_meta_read_valid),
    .io_meta_read_bits_idx(mshrs_io_meta_read_bits_idx),
    .io_meta_read_bits_way_en(mshrs_io_meta_read_bits_way_en),
    .io_meta_read_bits_tag(mshrs_io_meta_read_bits_tag),
    .io_meta_write_ready(mshrs_io_meta_write_ready),
    .io_meta_write_valid(mshrs_io_meta_write_valid),
    .io_meta_write_bits_idx(mshrs_io_meta_write_bits_idx),
    .io_meta_write_bits_way_en(mshrs_io_meta_write_bits_way_en),
    .io_meta_write_bits_data_tag(mshrs_io_meta_write_bits_data_tag),
    .io_meta_write_bits_data_coh_state(mshrs_io_meta_write_bits_data_coh_state),
    .io_replay_ready(mshrs_io_replay_ready),
    .io_replay_valid(mshrs_io_replay_valid),
    .io_replay_bits_addr(mshrs_io_replay_bits_addr),
    .io_replay_bits_tag(mshrs_io_replay_bits_tag),
    .io_replay_bits_cmd(mshrs_io_replay_bits_cmd),
    .io_replay_bits_typ(mshrs_io_replay_bits_typ),
    .io_replay_bits_phys(mshrs_io_replay_bits_phys),
    .io_replay_bits_data(mshrs_io_replay_bits_data),
    .io_mem_grant_valid(mshrs_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(mshrs_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(mshrs_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(mshrs_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(mshrs_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(mshrs_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(mshrs_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(mshrs_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(mshrs_io_mem_finish_ready),
    .io_mem_finish_valid(mshrs_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(mshrs_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(mshrs_io_mem_finish_bits_manager_id),
    .io_wb_req_ready(mshrs_io_wb_req_ready),
    .io_wb_req_valid(mshrs_io_wb_req_valid),
    .io_wb_req_bits_addr_beat(mshrs_io_wb_req_bits_addr_beat),
    .io_wb_req_bits_addr_block(mshrs_io_wb_req_bits_addr_block),
    .io_wb_req_bits_client_xact_id(mshrs_io_wb_req_bits_client_xact_id),
    .io_wb_req_bits_voluntary(mshrs_io_wb_req_bits_voluntary),
    .io_wb_req_bits_r_type(mshrs_io_wb_req_bits_r_type),
    .io_wb_req_bits_data(mshrs_io_wb_req_bits_data),
    .io_wb_req_bits_way_en(mshrs_io_wb_req_bits_way_en),
    .io_probe_rdy(mshrs_io_probe_rdy),
    .io_fence_rdy(mshrs_io_fence_rdy),
    .io_replay_next(mshrs_io_replay_next)
  );
  TLB dtlb (
    .clk(dtlb_clk),
    .reset(dtlb_reset),
    .io_req_ready(dtlb_io_req_ready),
    .io_req_valid(dtlb_io_req_valid),
    .io_req_bits_asid(dtlb_io_req_bits_asid),
    .io_req_bits_vpn(dtlb_io_req_bits_vpn),
    .io_req_bits_passthrough(dtlb_io_req_bits_passthrough),
    .io_req_bits_instruction(dtlb_io_req_bits_instruction),
    .io_req_bits_store(dtlb_io_req_bits_store),
    .io_resp_miss(dtlb_io_resp_miss),
    .io_resp_ppn(dtlb_io_resp_ppn),
    .io_resp_xcpt_ld(dtlb_io_resp_xcpt_ld),
    .io_resp_xcpt_st(dtlb_io_resp_xcpt_st),
    .io_resp_xcpt_if(dtlb_io_resp_xcpt_if),
    .io_resp_hit_idx(dtlb_io_resp_hit_idx),
    .io_ptw_req_ready(dtlb_io_ptw_req_ready),
    .io_ptw_req_valid(dtlb_io_ptw_req_valid),
    .io_ptw_req_bits_addr(dtlb_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(dtlb_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(dtlb_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(dtlb_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(dtlb_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(dtlb_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(dtlb_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(dtlb_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(dtlb_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(dtlb_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(dtlb_io_ptw_resp_bits_pte_v),
    .io_ptw_status_debug(dtlb_io_ptw_status_debug),
    .io_ptw_status_prv(dtlb_io_ptw_status_prv),
    .io_ptw_status_sd(dtlb_io_ptw_status_sd),
    .io_ptw_status_zero3(dtlb_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(dtlb_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(dtlb_io_ptw_status_zero2),
    .io_ptw_status_vm(dtlb_io_ptw_status_vm),
    .io_ptw_status_zero1(dtlb_io_ptw_status_zero1),
    .io_ptw_status_pum(dtlb_io_ptw_status_pum),
    .io_ptw_status_mprv(dtlb_io_ptw_status_mprv),
    .io_ptw_status_xs(dtlb_io_ptw_status_xs),
    .io_ptw_status_fs(dtlb_io_ptw_status_fs),
    .io_ptw_status_mpp(dtlb_io_ptw_status_mpp),
    .io_ptw_status_hpp(dtlb_io_ptw_status_hpp),
    .io_ptw_status_spp(dtlb_io_ptw_status_spp),
    .io_ptw_status_mpie(dtlb_io_ptw_status_mpie),
    .io_ptw_status_hpie(dtlb_io_ptw_status_hpie),
    .io_ptw_status_spie(dtlb_io_ptw_status_spie),
    .io_ptw_status_upie(dtlb_io_ptw_status_upie),
    .io_ptw_status_mie(dtlb_io_ptw_status_mie),
    .io_ptw_status_hie(dtlb_io_ptw_status_hie),
    .io_ptw_status_sie(dtlb_io_ptw_status_sie),
    .io_ptw_status_uie(dtlb_io_ptw_status_uie),
    .io_ptw_invalidate(dtlb_io_ptw_invalidate)
  );
  MetadataArray meta (
    .clk(meta_clk),
    .reset(meta_reset),
    .io_read_ready(meta_io_read_ready),
    .io_read_valid(meta_io_read_valid),
    .io_read_bits_idx(meta_io_read_bits_idx),
    .io_read_bits_way_en(meta_io_read_bits_way_en),
    .io_write_ready(meta_io_write_ready),
    .io_write_valid(meta_io_write_valid),
    .io_write_bits_idx(meta_io_write_bits_idx),
    .io_write_bits_way_en(meta_io_write_bits_way_en),
    .io_write_bits_data_tag(meta_io_write_bits_data_tag),
    .io_write_bits_data_coh_state(meta_io_write_bits_data_coh_state),
    .io_resp_0_tag(meta_io_resp_0_tag),
    .io_resp_0_coh_state(meta_io_resp_0_coh_state),
    .io_resp_1_tag(meta_io_resp_1_tag),
    .io_resp_1_coh_state(meta_io_resp_1_coh_state),
    .io_resp_2_tag(meta_io_resp_2_tag),
    .io_resp_2_coh_state(meta_io_resp_2_coh_state),
    .io_resp_3_tag(meta_io_resp_3_tag),
    .io_resp_3_coh_state(meta_io_resp_3_coh_state)
  );
  Arbiter_83 metaReadArb (
    .clk(metaReadArb_clk),
    .reset(metaReadArb_reset),
    .io_in_0_ready(metaReadArb_io_in_0_ready),
    .io_in_0_valid(metaReadArb_io_in_0_valid),
    .io_in_0_bits_idx(metaReadArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaReadArb_io_in_0_bits_way_en),
    .io_in_1_ready(metaReadArb_io_in_1_ready),
    .io_in_1_valid(metaReadArb_io_in_1_valid),
    .io_in_1_bits_idx(metaReadArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaReadArb_io_in_1_bits_way_en),
    .io_in_2_ready(metaReadArb_io_in_2_ready),
    .io_in_2_valid(metaReadArb_io_in_2_valid),
    .io_in_2_bits_idx(metaReadArb_io_in_2_bits_idx),
    .io_in_2_bits_way_en(metaReadArb_io_in_2_bits_way_en),
    .io_in_3_ready(metaReadArb_io_in_3_ready),
    .io_in_3_valid(metaReadArb_io_in_3_valid),
    .io_in_3_bits_idx(metaReadArb_io_in_3_bits_idx),
    .io_in_3_bits_way_en(metaReadArb_io_in_3_bits_way_en),
    .io_in_4_ready(metaReadArb_io_in_4_ready),
    .io_in_4_valid(metaReadArb_io_in_4_valid),
    .io_in_4_bits_idx(metaReadArb_io_in_4_bits_idx),
    .io_in_4_bits_way_en(metaReadArb_io_in_4_bits_way_en),
    .io_out_ready(metaReadArb_io_out_ready),
    .io_out_valid(metaReadArb_io_out_valid),
    .io_out_bits_idx(metaReadArb_io_out_bits_idx),
    .io_out_bits_way_en(metaReadArb_io_out_bits_way_en),
    .io_chosen(metaReadArb_io_chosen)
  );
  Arbiter_68 metaWriteArb (
    .clk(metaWriteArb_clk),
    .reset(metaWriteArb_reset),
    .io_in_0_ready(metaWriteArb_io_in_0_ready),
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_idx(metaWriteArb_io_in_0_bits_idx),
    .io_in_0_bits_way_en(metaWriteArb_io_in_0_bits_way_en),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_coh_state(metaWriteArb_io_in_0_bits_data_coh_state),
    .io_in_1_ready(metaWriteArb_io_in_1_ready),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_idx(metaWriteArb_io_in_1_bits_idx),
    .io_in_1_bits_way_en(metaWriteArb_io_in_1_bits_way_en),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_coh_state(metaWriteArb_io_in_1_bits_data_coh_state),
    .io_out_ready(metaWriteArb_io_out_ready),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_idx(metaWriteArb_io_out_bits_idx),
    .io_out_bits_way_en(metaWriteArb_io_out_bits_way_en),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_coh_state(metaWriteArb_io_out_bits_data_coh_state),
    .io_chosen(metaWriteArb_io_chosen)
  );
  DataArray data (
    .clk(data_clk),
    .reset(data_reset),
    .io_read_ready(data_io_read_ready),
    .io_read_valid(data_io_read_valid),
    .io_read_bits_way_en(data_io_read_bits_way_en),
    .io_read_bits_addr(data_io_read_bits_addr),
    .io_write_ready(data_io_write_ready),
    .io_write_valid(data_io_write_valid),
    .io_write_bits_way_en(data_io_write_bits_way_en),
    .io_write_bits_addr(data_io_write_bits_addr),
    .io_write_bits_wmask(data_io_write_bits_wmask),
    .io_write_bits_data(data_io_write_bits_data),
    .io_resp_0(data_io_resp_0),
    .io_resp_1(data_io_resp_1),
    .io_resp_2(data_io_resp_2),
    .io_resp_3(data_io_resp_3)
  );
  Arbiter_85 readArb (
    .clk(readArb_clk),
    .reset(readArb_reset),
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_way_en(readArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(readArb_io_in_0_bits_addr),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_way_en(readArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(readArb_io_in_1_bits_addr),
    .io_in_2_ready(readArb_io_in_2_ready),
    .io_in_2_valid(readArb_io_in_2_valid),
    .io_in_2_bits_way_en(readArb_io_in_2_bits_way_en),
    .io_in_2_bits_addr(readArb_io_in_2_bits_addr),
    .io_in_3_ready(readArb_io_in_3_ready),
    .io_in_3_valid(readArb_io_in_3_valid),
    .io_in_3_bits_way_en(readArb_io_in_3_bits_way_en),
    .io_in_3_bits_addr(readArb_io_in_3_bits_addr),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_way_en(readArb_io_out_bits_way_en),
    .io_out_bits_addr(readArb_io_out_bits_addr),
    .io_chosen(readArb_io_chosen)
  );
  Arbiter_86 writeArb (
    .clk(writeArb_clk),
    .reset(writeArb_reset),
    .io_in_0_ready(writeArb_io_in_0_ready),
    .io_in_0_valid(writeArb_io_in_0_valid),
    .io_in_0_bits_way_en(writeArb_io_in_0_bits_way_en),
    .io_in_0_bits_addr(writeArb_io_in_0_bits_addr),
    .io_in_0_bits_wmask(writeArb_io_in_0_bits_wmask),
    .io_in_0_bits_data(writeArb_io_in_0_bits_data),
    .io_in_1_ready(writeArb_io_in_1_ready),
    .io_in_1_valid(writeArb_io_in_1_valid),
    .io_in_1_bits_way_en(writeArb_io_in_1_bits_way_en),
    .io_in_1_bits_addr(writeArb_io_in_1_bits_addr),
    .io_in_1_bits_wmask(writeArb_io_in_1_bits_wmask),
    .io_in_1_bits_data(writeArb_io_in_1_bits_data),
    .io_out_ready(writeArb_io_out_ready),
    .io_out_valid(writeArb_io_out_valid),
    .io_out_bits_way_en(writeArb_io_out_bits_way_en),
    .io_out_bits_addr(writeArb_io_out_bits_addr),
    .io_out_bits_wmask(writeArb_io_out_bits_wmask),
    .io_out_bits_data(writeArb_io_out_bits_data),
    .io_chosen(writeArb_io_chosen)
  );
  AMOALU amoalu (
    .clk(amoalu_clk),
    .reset(amoalu_reset),
    .io_addr(amoalu_io_addr),
    .io_cmd(amoalu_io_cmd),
    .io_typ(amoalu_io_typ),
    .io_lhs(amoalu_io_lhs),
    .io_rhs(amoalu_io_rhs),
    .io_out(amoalu_io_out)
  );
  LockingArbiter_87 releaseArb (
    .clk(releaseArb_clk),
    .reset(releaseArb_reset),
    .io_in_0_ready(releaseArb_io_in_0_ready),
    .io_in_0_valid(releaseArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(releaseArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(releaseArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(releaseArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(releaseArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(releaseArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(releaseArb_io_in_0_bits_data),
    .io_in_1_ready(releaseArb_io_in_1_ready),
    .io_in_1_valid(releaseArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(releaseArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(releaseArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(releaseArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(releaseArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(releaseArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(releaseArb_io_in_1_bits_data),
    .io_out_ready(releaseArb_io_out_ready),
    .io_out_valid(releaseArb_io_out_valid),
    .io_out_bits_addr_beat(releaseArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(releaseArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(releaseArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(releaseArb_io_out_bits_voluntary),
    .io_out_bits_r_type(releaseArb_io_out_bits_r_type),
    .io_out_bits_data(releaseArb_io_out_bits_data),
    .io_chosen(releaseArb_io_chosen)
  );
  FlowThroughSerializer_88 FlowThroughSerializer_88_5908 (
    .clk(FlowThroughSerializer_88_5908_clk),
    .reset(FlowThroughSerializer_88_5908_reset),
    .io_in_ready(FlowThroughSerializer_88_5908_io_in_ready),
    .io_in_valid(FlowThroughSerializer_88_5908_io_in_valid),
    .io_in_bits_addr_beat(FlowThroughSerializer_88_5908_io_in_bits_addr_beat),
    .io_in_bits_client_xact_id(FlowThroughSerializer_88_5908_io_in_bits_client_xact_id),
    .io_in_bits_manager_xact_id(FlowThroughSerializer_88_5908_io_in_bits_manager_xact_id),
    .io_in_bits_is_builtin_type(FlowThroughSerializer_88_5908_io_in_bits_is_builtin_type),
    .io_in_bits_g_type(FlowThroughSerializer_88_5908_io_in_bits_g_type),
    .io_in_bits_data(FlowThroughSerializer_88_5908_io_in_bits_data),
    .io_in_bits_manager_id(FlowThroughSerializer_88_5908_io_in_bits_manager_id),
    .io_out_ready(FlowThroughSerializer_88_5908_io_out_ready),
    .io_out_valid(FlowThroughSerializer_88_5908_io_out_valid),
    .io_out_bits_addr_beat(FlowThroughSerializer_88_5908_io_out_bits_addr_beat),
    .io_out_bits_client_xact_id(FlowThroughSerializer_88_5908_io_out_bits_client_xact_id),
    .io_out_bits_manager_xact_id(FlowThroughSerializer_88_5908_io_out_bits_manager_xact_id),
    .io_out_bits_is_builtin_type(FlowThroughSerializer_88_5908_io_out_bits_is_builtin_type),
    .io_out_bits_g_type(FlowThroughSerializer_88_5908_io_out_bits_g_type),
    .io_out_bits_data(FlowThroughSerializer_88_5908_io_out_bits_data),
    .io_out_bits_manager_id(FlowThroughSerializer_88_5908_io_out_bits_manager_id),
    .io_cnt(FlowThroughSerializer_88_5908_io_cnt),
    .io_done(FlowThroughSerializer_88_5908_io_done)
  );
  Arbiter_70 wbArb (
    .clk(wbArb_clk),
    .reset(wbArb_reset),
    .io_in_0_ready(wbArb_io_in_0_ready),
    .io_in_0_valid(wbArb_io_in_0_valid),
    .io_in_0_bits_addr_beat(wbArb_io_in_0_bits_addr_beat),
    .io_in_0_bits_addr_block(wbArb_io_in_0_bits_addr_block),
    .io_in_0_bits_client_xact_id(wbArb_io_in_0_bits_client_xact_id),
    .io_in_0_bits_voluntary(wbArb_io_in_0_bits_voluntary),
    .io_in_0_bits_r_type(wbArb_io_in_0_bits_r_type),
    .io_in_0_bits_data(wbArb_io_in_0_bits_data),
    .io_in_0_bits_way_en(wbArb_io_in_0_bits_way_en),
    .io_in_1_ready(wbArb_io_in_1_ready),
    .io_in_1_valid(wbArb_io_in_1_valid),
    .io_in_1_bits_addr_beat(wbArb_io_in_1_bits_addr_beat),
    .io_in_1_bits_addr_block(wbArb_io_in_1_bits_addr_block),
    .io_in_1_bits_client_xact_id(wbArb_io_in_1_bits_client_xact_id),
    .io_in_1_bits_voluntary(wbArb_io_in_1_bits_voluntary),
    .io_in_1_bits_r_type(wbArb_io_in_1_bits_r_type),
    .io_in_1_bits_data(wbArb_io_in_1_bits_data),
    .io_in_1_bits_way_en(wbArb_io_in_1_bits_way_en),
    .io_out_ready(wbArb_io_out_ready),
    .io_out_valid(wbArb_io_out_valid),
    .io_out_bits_addr_beat(wbArb_io_out_bits_addr_beat),
    .io_out_bits_addr_block(wbArb_io_out_bits_addr_block),
    .io_out_bits_client_xact_id(wbArb_io_out_bits_client_xact_id),
    .io_out_bits_voluntary(wbArb_io_out_bits_voluntary),
    .io_out_bits_r_type(wbArb_io_out_bits_r_type),
    .io_out_bits_data(wbArb_io_out_bits_data),
    .io_out_bits_way_en(wbArb_io_out_bits_way_en),
    .io_chosen(wbArb_io_chosen)
  );
  assign io_cpu_req_ready = GEN_82;
  assign io_cpu_s2_nack = T_7059;
  assign io_cpu_resp_valid = T_7060_valid;
  assign io_cpu_resp_bits_addr = T_7060_bits_addr;
  assign io_cpu_resp_bits_tag = T_7060_bits_tag;
  assign io_cpu_resp_bits_cmd = T_7060_bits_cmd;
  assign io_cpu_resp_bits_typ = T_7060_bits_typ;
  assign io_cpu_resp_bits_data = T_7060_bits_data;
  assign io_cpu_resp_bits_replay = T_7060_bits_replay;
  assign io_cpu_resp_bits_has_data = T_7060_bits_has_data;
  assign io_cpu_resp_bits_data_word_bypass = T_6617;
  assign io_cpu_resp_bits_store_data = T_7060_bits_store_data;
  assign io_cpu_replay_next = T_7246;
  assign io_cpu_xcpt_ma_ld = T_2361;
  assign io_cpu_xcpt_ma_st = T_2362;
  assign io_cpu_xcpt_pf_ld = T_2363;
  assign io_cpu_xcpt_pf_st = T_2364;
  assign io_cpu_ordered = T_7244;
  assign io_ptw_req_valid = dtlb_io_ptw_req_valid;
  assign io_ptw_req_bits_addr = dtlb_io_ptw_req_bits_addr;
  assign io_ptw_req_bits_prv = dtlb_io_ptw_req_bits_prv;
  assign io_ptw_req_bits_store = dtlb_io_ptw_req_bits_store;
  assign io_ptw_req_bits_fetch = dtlb_io_ptw_req_bits_fetch;
  assign io_mem_acquire_valid = mshrs_io_mem_req_valid;
  assign io_mem_acquire_bits_addr_block = mshrs_io_mem_req_bits_addr_block;
  assign io_mem_acquire_bits_client_xact_id = mshrs_io_mem_req_bits_client_xact_id;
  assign io_mem_acquire_bits_addr_beat = mshrs_io_mem_req_bits_addr_beat;
  assign io_mem_acquire_bits_is_builtin_type = mshrs_io_mem_req_bits_is_builtin_type;
  assign io_mem_acquire_bits_a_type = mshrs_io_mem_req_bits_a_type;
  assign io_mem_acquire_bits_union = mshrs_io_mem_req_bits_union;
  assign io_mem_acquire_bits_data = mshrs_io_mem_req_bits_data;
  assign io_mem_probe_ready = T_5907;
  assign io_mem_release_valid = releaseArb_io_out_valid;
  assign io_mem_release_bits_addr_beat = releaseArb_io_out_bits_addr_beat;
  assign io_mem_release_bits_addr_block = releaseArb_io_out_bits_addr_block;
  assign io_mem_release_bits_client_xact_id = releaseArb_io_out_bits_client_xact_id;
  assign io_mem_release_bits_voluntary = releaseArb_io_out_bits_voluntary;
  assign io_mem_release_bits_r_type = releaseArb_io_out_bits_r_type;
  assign io_mem_release_bits_data = releaseArb_io_out_bits_data;
  assign io_mem_grant_ready = FlowThroughSerializer_88_5908_io_in_ready;
  assign io_mem_finish_valid = mshrs_io_mem_finish_valid;
  assign io_mem_finish_bits_manager_xact_id = mshrs_io_mem_finish_bits_manager_xact_id;
  assign io_mem_finish_bits_manager_id = mshrs_io_mem_finish_bits_manager_id;
  assign wb_clk = clk;
  assign wb_reset = reset;
  assign wb_io_req_valid = wbArb_io_out_valid;
  assign wb_io_req_bits_addr_beat = wbArb_io_out_bits_addr_beat;
  assign wb_io_req_bits_addr_block = wbArb_io_out_bits_addr_block;
  assign wb_io_req_bits_client_xact_id = wbArb_io_out_bits_client_xact_id;
  assign wb_io_req_bits_voluntary = wbArb_io_out_bits_voluntary;
  assign wb_io_req_bits_r_type = wbArb_io_out_bits_r_type;
  assign wb_io_req_bits_data = wbArb_io_out_bits_data;
  assign wb_io_req_bits_way_en = wbArb_io_out_bits_way_en;
  assign wb_io_meta_read_ready = metaReadArb_io_in_3_ready;
  assign wb_io_data_req_ready = readArb_io_in_2_ready;
  assign wb_io_data_resp = T_3548_0;
  assign wb_io_release_ready = releaseArb_io_in_0_ready;
  assign prober_clk = clk;
  assign prober_reset = reset;
  assign prober_io_req_valid = T_5904;
  assign prober_io_req_bits_addr_block = io_mem_probe_bits_addr_block;
  assign prober_io_req_bits_p_type = io_mem_probe_bits_p_type;
  assign prober_io_req_bits_client_xact_id = GEN_68;
  assign prober_io_rep_ready = releaseArb_io_in_1_ready;
  assign prober_io_meta_read_ready = metaReadArb_io_in_2_ready;
  assign prober_io_meta_write_ready = metaWriteArb_io_in_1_ready;
  assign prober_io_wb_req_ready = wbArb_io_in_0_ready;
  assign prober_io_way_en = s2_tag_match_way;
  assign prober_io_mshr_rdy = mshrs_io_probe_rdy;
  assign prober_io_block_state_state = s2_hit_state_state;
  assign mshrs_clk = clk;
  assign mshrs_reset = reset;
  assign mshrs_io_req_valid = GEN_80;
  assign mshrs_io_req_bits_addr = s2_req_addr;
  assign mshrs_io_req_bits_tag = s2_req_tag;
  assign mshrs_io_req_bits_cmd = s2_req_cmd;
  assign mshrs_io_req_bits_typ = s2_req_typ;
  assign mshrs_io_req_bits_phys = s2_req_phys;
  assign mshrs_io_req_bits_data = s2_req_data;
  assign mshrs_io_req_bits_tag_match = s2_tag_match;
  assign mshrs_io_req_bits_old_meta_tag = T_5770_tag;
  assign mshrs_io_req_bits_old_meta_coh_state = T_5770_coh_state;
  assign mshrs_io_req_bits_way_en = T_5866;
  assign mshrs_io_resp_ready = T_7058;
  assign mshrs_io_mem_req_ready = io_mem_acquire_ready;
  assign mshrs_io_meta_read_ready = metaReadArb_io_in_1_ready;
  assign mshrs_io_meta_write_ready = metaWriteArb_io_in_0_ready;
  assign mshrs_io_replay_ready = readArb_io_in_1_ready;
  assign mshrs_io_mem_grant_valid = T_5909;
  assign mshrs_io_mem_grant_bits_addr_beat = FlowThroughSerializer_88_5908_io_out_bits_addr_beat;
  assign mshrs_io_mem_grant_bits_client_xact_id = FlowThroughSerializer_88_5908_io_out_bits_client_xact_id;
  assign mshrs_io_mem_grant_bits_manager_xact_id = FlowThroughSerializer_88_5908_io_out_bits_manager_xact_id;
  assign mshrs_io_mem_grant_bits_is_builtin_type = FlowThroughSerializer_88_5908_io_out_bits_is_builtin_type;
  assign mshrs_io_mem_grant_bits_g_type = FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign mshrs_io_mem_grant_bits_data = FlowThroughSerializer_88_5908_io_out_bits_data;
  assign mshrs_io_mem_grant_bits_manager_id = FlowThroughSerializer_88_5908_io_out_bits_manager_id;
  assign mshrs_io_mem_finish_ready = io_mem_finish_ready;
  assign mshrs_io_wb_req_ready = wbArb_io_in_1_ready;
  assign T_2075 = io_cpu_req_ready & io_cpu_req_valid;
  assign T_2153 = io_cpu_s1_kill == 1'h0;
  assign s1_valid_masked = s1_valid & T_2153;
  assign T_2234 = s2_req_cmd != 5'h5;
  assign s2_replay = T_2233 & T_2234;
  assign s2_recycle = T_6182;
  assign s2_valid_masked = T_6177;
  assign GEN_0 = s1_clk_en ? s2_recycle : s1_recycled;
  assign T_2315 = s1_req_cmd == 5'h0;
  assign T_2316 = s1_req_cmd == 5'h6;
  assign T_2317 = T_2315 | T_2316;
  assign T_2318 = s1_req_cmd == 5'h7;
  assign T_2319 = T_2317 | T_2318;
  assign T_2320 = s1_req_cmd[3];
  assign T_2321 = s1_req_cmd == 5'h4;
  assign T_2322 = T_2320 | T_2321;
  assign s1_read = T_2319 | T_2322;
  assign T_2323 = s1_req_cmd == 5'h1;
  assign T_2325 = T_2323 | T_2318;
  assign s1_write = T_2325 | T_2322;
  assign T_2329 = s1_read | s1_write;
  assign T_2330 = s1_req_cmd == 5'h2;
  assign T_2331 = s1_req_cmd == 5'h3;
  assign T_2332 = T_2330 | T_2331;
  assign s1_readwrite = T_2329 | T_2332;
  assign dtlb_clk = clk;
  assign dtlb_reset = reset;
  assign dtlb_io_req_valid = T_2333;
  assign dtlb_io_req_bits_asid = {{6'd0}, 1'h0};
  assign dtlb_io_req_bits_vpn = T_2335;
  assign dtlb_io_req_bits_passthrough = s1_req_phys;
  assign dtlb_io_req_bits_instruction = 1'h0;
  assign dtlb_io_req_bits_store = s1_write;
  assign dtlb_io_ptw_req_ready = io_ptw_req_ready;
  assign dtlb_io_ptw_resp_valid = io_ptw_resp_valid;
  assign dtlb_io_ptw_resp_bits_pte_ppn = io_ptw_resp_bits_pte_ppn;
  assign dtlb_io_ptw_resp_bits_pte_reserved_for_software = io_ptw_resp_bits_pte_reserved_for_software;
  assign dtlb_io_ptw_resp_bits_pte_d = io_ptw_resp_bits_pte_d;
  assign dtlb_io_ptw_resp_bits_pte_r = io_ptw_resp_bits_pte_r;
  assign dtlb_io_ptw_resp_bits_pte_typ = io_ptw_resp_bits_pte_typ;
  assign dtlb_io_ptw_resp_bits_pte_v = io_ptw_resp_bits_pte_v;
  assign dtlb_io_ptw_status_debug = io_ptw_status_debug;
  assign dtlb_io_ptw_status_prv = io_ptw_status_prv;
  assign dtlb_io_ptw_status_sd = io_ptw_status_sd;
  assign dtlb_io_ptw_status_zero3 = io_ptw_status_zero3;
  assign dtlb_io_ptw_status_sd_rv32 = io_ptw_status_sd_rv32;
  assign dtlb_io_ptw_status_zero2 = io_ptw_status_zero2;
  assign dtlb_io_ptw_status_vm = io_ptw_status_vm;
  assign dtlb_io_ptw_status_zero1 = io_ptw_status_zero1;
  assign dtlb_io_ptw_status_pum = io_ptw_status_pum;
  assign dtlb_io_ptw_status_mprv = io_ptw_status_mprv;
  assign dtlb_io_ptw_status_xs = io_ptw_status_xs;
  assign dtlb_io_ptw_status_fs = io_ptw_status_fs;
  assign dtlb_io_ptw_status_mpp = io_ptw_status_mpp;
  assign dtlb_io_ptw_status_hpp = io_ptw_status_hpp;
  assign dtlb_io_ptw_status_spp = io_ptw_status_spp;
  assign dtlb_io_ptw_status_mpie = io_ptw_status_mpie;
  assign dtlb_io_ptw_status_hpie = io_ptw_status_hpie;
  assign dtlb_io_ptw_status_spie = io_ptw_status_spie;
  assign dtlb_io_ptw_status_upie = io_ptw_status_upie;
  assign dtlb_io_ptw_status_mie = io_ptw_status_mie;
  assign dtlb_io_ptw_status_hie = io_ptw_status_hie;
  assign dtlb_io_ptw_status_sie = io_ptw_status_sie;
  assign dtlb_io_ptw_status_uie = io_ptw_status_uie;
  assign dtlb_io_ptw_invalidate = io_ptw_invalidate;
  assign T_2333 = s1_valid_masked & s1_readwrite;
  assign T_2335 = s1_req_addr[39:12];
  assign T_2338 = dtlb_io_req_ready == 1'h0;
  assign T_2340 = io_cpu_req_bits_phys == 1'h0;
  assign T_2341 = T_2338 & T_2340;
  assign GEN_1 = T_2341 ? 1'h0 : 1'h1;
  assign GEN_2 = io_cpu_req_valid ? io_cpu_req_bits_addr : s1_req_addr;
  assign GEN_3 = io_cpu_req_valid ? io_cpu_req_bits_tag : s1_req_tag;
  assign GEN_4 = io_cpu_req_valid ? io_cpu_req_bits_cmd : s1_req_cmd;
  assign GEN_5 = io_cpu_req_valid ? io_cpu_req_bits_typ : s1_req_typ;
  assign GEN_6 = io_cpu_req_valid ? io_cpu_req_bits_phys : s1_req_phys;
  assign GEN_7 = io_cpu_req_valid ? io_cpu_req_bits_data : s1_req_data;
  assign T_2343 = {wb_io_meta_read_bits_tag,wb_io_meta_read_bits_idx};
  assign GEN_83 = {{6'd0}, T_2343};
  assign T_2344 = GEN_83 << 6;
  assign GEN_8 = wb_io_meta_read_valid ? {{8'd0}, T_2344} : GEN_2;
  assign GEN_9 = wb_io_meta_read_valid ? 1'h1 : GEN_6;
  assign T_2346 = {prober_io_meta_read_bits_tag,prober_io_meta_read_bits_idx};
  assign GEN_84 = {{6'd0}, T_2346};
  assign T_2347 = GEN_84 << 6;
  assign GEN_10 = prober_io_meta_read_valid ? {{8'd0}, T_2347} : GEN_8;
  assign GEN_11 = prober_io_meta_read_valid ? 1'h1 : GEN_9;
  assign GEN_12 = mshrs_io_replay_valid ? mshrs_io_replay_bits_addr : GEN_10;
  assign GEN_13 = mshrs_io_replay_valid ? mshrs_io_replay_bits_tag : GEN_3;
  assign GEN_14 = mshrs_io_replay_valid ? mshrs_io_replay_bits_cmd : GEN_4;
  assign GEN_15 = mshrs_io_replay_valid ? mshrs_io_replay_bits_typ : GEN_5;
  assign GEN_16 = mshrs_io_replay_valid ? mshrs_io_replay_bits_phys : GEN_11;
  assign GEN_17 = mshrs_io_replay_valid ? mshrs_io_replay_bits_data : GEN_7;
  assign GEN_18 = s2_recycle ? s2_req_addr : GEN_12;
  assign GEN_19 = s2_recycle ? s2_req_tag : GEN_13;
  assign GEN_20 = s2_recycle ? s2_req_cmd : GEN_14;
  assign GEN_21 = s2_recycle ? s2_req_typ : GEN_15;
  assign GEN_22 = s2_recycle ? s2_req_phys : GEN_16;
  assign GEN_23 = s2_recycle ? s2_req_data : GEN_17;
  assign T_2349 = s1_req_addr[11:0];
  assign s1_addr = {dtlb_io_resp_ppn,T_2349};
  assign T_2350 = s1_replay ? mshrs_io_replay_bits_data : io_cpu_s1_data;
  assign GEN_24 = s1_write ? T_2350 : s2_req_data;
  assign GEN_25 = s1_recycled ? s1_req_data : GEN_24;
  assign GEN_26 = s1_clk_en ? s1_req_typ : s2_req_typ;
  assign GEN_27 = s1_clk_en ? s1_req_phys : s2_req_phys;
  assign GEN_28 = s1_clk_en ? {{8'd0}, s1_addr} : s2_req_addr;
  assign GEN_29 = s1_clk_en ? GEN_25 : s2_req_data;
  assign GEN_30 = s1_clk_en ? s1_req_tag : s2_req_tag;
  assign GEN_31 = s1_clk_en ? s1_req_cmd : s2_req_cmd;
  assign T_2352 = s1_req_typ[1:0];
  assign GEN_85 = {{3'd0}, 1'h1};
  assign T_2354 = GEN_85 << T_2352;
  assign T_2356 = T_2354 - GEN_85;
  assign T_2357 = T_2356[3:0];
  assign T_2358 = T_2357[2:0];
  assign GEN_87 = {{37'd0}, T_2358};
  assign T_2359 = s1_req_addr & GEN_87;
  assign GEN_88 = {{39'd0}, 1'h0};
  assign misaligned = T_2359 != GEN_88;
  assign T_2361 = s1_read & misaligned;
  assign T_2362 = s1_write & misaligned;
  assign T_2363 = s1_read & dtlb_io_resp_xcpt_ld;
  assign T_2364 = s1_write & dtlb_io_resp_xcpt_st;
  assign T_2365 = io_cpu_xcpt_ma_ld | io_cpu_xcpt_ma_st;
  assign T_2366 = T_2365 | io_cpu_xcpt_pf_ld;
  assign T_2367 = T_2366 | io_cpu_xcpt_pf_st;
  assign T_2369 = T_2368 & s2_valid_masked;
  assign T_2371 = T_2369 == 1'h0;
  assign T_2372 = T_2371 | reset;
  assign T_2374 = T_2372 == 1'h0;
  assign meta_clk = clk;
  assign meta_reset = reset;
  assign meta_io_read_valid = metaReadArb_io_out_valid;
  assign meta_io_read_bits_idx = metaReadArb_io_out_bits_idx;
  assign meta_io_read_bits_way_en = metaReadArb_io_out_bits_way_en;
  assign meta_io_write_valid = metaWriteArb_io_out_valid;
  assign meta_io_write_bits_idx = metaWriteArb_io_out_bits_idx;
  assign meta_io_write_bits_way_en = metaWriteArb_io_out_bits_way_en;
  assign meta_io_write_bits_data_tag = metaWriteArb_io_out_bits_data_tag;
  assign meta_io_write_bits_data_coh_state = metaWriteArb_io_out_bits_data_coh_state;
  assign metaReadArb_clk = clk;
  assign metaReadArb_reset = reset;
  assign metaReadArb_io_in_0_valid = s2_recycle;
  assign metaReadArb_io_in_0_bits_idx = T_2775[5:0];
  assign metaReadArb_io_in_0_bits_way_en = GEN_76;
  assign metaReadArb_io_in_1_valid = mshrs_io_meta_read_valid;
  assign metaReadArb_io_in_1_bits_idx = mshrs_io_meta_read_bits_idx;
  assign metaReadArb_io_in_1_bits_way_en = mshrs_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_2_valid = prober_io_meta_read_valid;
  assign metaReadArb_io_in_2_bits_idx = prober_io_meta_read_bits_idx;
  assign metaReadArb_io_in_2_bits_way_en = prober_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_3_valid = wb_io_meta_read_valid;
  assign metaReadArb_io_in_3_bits_idx = wb_io_meta_read_bits_idx;
  assign metaReadArb_io_in_3_bits_way_en = wb_io_meta_read_bits_way_en;
  assign metaReadArb_io_in_4_valid = io_cpu_req_valid;
  assign metaReadArb_io_in_4_bits_idx = T_2766[5:0];
  assign metaReadArb_io_in_4_bits_way_en = GEN_86;
  assign metaReadArb_io_out_ready = meta_io_read_ready;
  assign metaWriteArb_clk = clk;
  assign metaWriteArb_reset = reset;
  assign metaWriteArb_io_in_0_valid = mshrs_io_meta_write_valid;
  assign metaWriteArb_io_in_0_bits_idx = mshrs_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_0_bits_way_en = mshrs_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_0_bits_data_tag = mshrs_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_0_bits_data_coh_state = mshrs_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_in_1_valid = prober_io_meta_write_valid;
  assign metaWriteArb_io_in_1_bits_idx = prober_io_meta_write_bits_idx;
  assign metaWriteArb_io_in_1_bits_way_en = prober_io_meta_write_bits_way_en;
  assign metaWriteArb_io_in_1_bits_data_tag = prober_io_meta_write_bits_data_tag;
  assign metaWriteArb_io_in_1_bits_data_coh_state = prober_io_meta_write_bits_data_coh_state;
  assign metaWriteArb_io_out_ready = meta_io_write_ready;
  assign data_clk = clk;
  assign data_reset = reset;
  assign data_io_read_valid = readArb_io_out_valid;
  assign data_io_read_bits_way_en = readArb_io_out_bits_way_en;
  assign data_io_read_bits_addr = readArb_io_out_bits_addr;
  assign data_io_write_valid = writeArb_io_out_valid;
  assign data_io_write_bits_way_en = writeArb_io_out_bits_way_en;
  assign data_io_write_bits_addr = writeArb_io_out_bits_addr;
  assign data_io_write_bits_wmask = writeArb_io_out_bits_wmask;
  assign data_io_write_bits_data = T_2765;
  assign readArb_clk = clk;
  assign readArb_reset = reset;
  assign readArb_io_in_0_valid = s2_recycle;
  assign readArb_io_in_0_bits_way_en = 4'hf;
  assign readArb_io_in_0_bits_addr = s2_req_addr[11:0];
  assign readArb_io_in_1_valid = mshrs_io_replay_valid;
  assign readArb_io_in_1_bits_way_en = 4'hf;
  assign readArb_io_in_1_bits_addr = mshrs_io_replay_bits_addr[11:0];
  assign readArb_io_in_2_valid = wb_io_data_req_valid;
  assign readArb_io_in_2_bits_way_en = wb_io_data_req_bits_way_en;
  assign readArb_io_in_2_bits_addr = wb_io_data_req_bits_addr;
  assign readArb_io_in_3_valid = io_cpu_req_valid;
  assign readArb_io_in_3_bits_way_en = 4'hf;
  assign readArb_io_in_3_bits_addr = io_cpu_req_bits_addr[11:0];
  assign readArb_io_out_ready = T_5976;
  assign writeArb_clk = clk;
  assign writeArb_reset = reset;
  assign writeArb_io_in_0_valid = s3_valid;
  assign writeArb_io_in_0_bits_way_en = s3_way;
  assign writeArb_io_in_0_bits_addr = s3_req_addr[11:0];
  assign writeArb_io_in_0_bits_wmask = rowWMask[0];
  assign writeArb_io_in_0_bits_data = s3_req_data;
  assign writeArb_io_in_1_valid = T_5970;
  assign writeArb_io_in_1_bits_way_en = mshrs_io_refill_way_en;
  assign writeArb_io_in_1_bits_addr = mshrs_io_refill_addr;
  assign writeArb_io_in_1_bits_wmask = 1'h1;
  assign writeArb_io_in_1_bits_data = T_5973;
  assign writeArb_io_out_ready = data_io_write_ready;
  assign T_2765 = writeArb_io_out_bits_data;
  assign T_2766 = io_cpu_req_bits_addr[39:6];
  assign T_2768 = metaReadArb_io_in_4_ready == 1'h0;
  assign GEN_32 = T_2768 ? 1'h0 : GEN_1;
  assign T_2773 = readArb_io_in_3_ready == 1'h0;
  assign GEN_33 = T_2773 ? 1'h0 : GEN_32;
  assign T_2775 = s2_req_addr[39:6];
  assign T_2778 = s1_addr[31:12];
  assign T_2779 = meta_io_resp_0_tag == T_2778;
  assign T_2781 = meta_io_resp_1_tag == T_2778;
  assign T_2783 = meta_io_resp_2_tag == T_2778;
  assign T_2785 = meta_io_resp_3_tag == T_2778;
  assign T_2791_0 = T_2779;
  assign T_2791_1 = T_2781;
  assign T_2791_2 = T_2783;
  assign T_2791_3 = T_2785;
  assign T_2793 = {T_2791_1,T_2791_0};
  assign T_2794 = {T_2791_3,T_2791_2};
  assign s1_tag_eq_way = {T_2794,T_2793};
  assign T_2795 = s1_tag_eq_way[0];
  assign T_2796 = meta_io_resp_0_coh_state != 2'h0;
  assign T_2797 = T_2795 & T_2796;
  assign T_2798 = s1_tag_eq_way[1];
  assign T_2799 = meta_io_resp_1_coh_state != 2'h0;
  assign T_2800 = T_2798 & T_2799;
  assign T_2801 = s1_tag_eq_way[2];
  assign T_2802 = meta_io_resp_2_coh_state != 2'h0;
  assign T_2803 = T_2801 & T_2802;
  assign T_2804 = s1_tag_eq_way[3];
  assign T_2805 = meta_io_resp_3_coh_state != 2'h0;
  assign T_2806 = T_2804 & T_2805;
  assign T_2812_0 = T_2797;
  assign T_2812_1 = T_2800;
  assign T_2812_2 = T_2803;
  assign T_2812_3 = T_2806;
  assign T_2814 = {T_2812_1,T_2812_0};
  assign T_2815 = {T_2812_3,T_2812_2};
  assign s1_tag_match_way = {T_2815,T_2814};
  assign T_2817 = s1_valid == 1'h0;
  assign GEN_34 = s1_clk_en ? s1_tag_match_way : s2_tag_match_way;
  assign GEN_89 = {{3'd0}, 1'h0};
  assign s2_tag_match = s2_tag_match_way != GEN_89;
  assign GEN_35 = s1_clk_en ? meta_io_resp_0_coh_state : T_2822_state;
  assign GEN_36 = s1_clk_en ? meta_io_resp_1_coh_state : T_2847_state;
  assign GEN_37 = s1_clk_en ? meta_io_resp_2_coh_state : T_2872_state;
  assign GEN_38 = s1_clk_en ? meta_io_resp_3_coh_state : T_2897_state;
  assign T_3119_0_state = T_2822_state;
  assign T_3119_1_state = T_2847_state;
  assign T_3119_2_state = T_2872_state;
  assign T_3119_3_state = T_2897_state;
  assign T_3241 = s2_tag_match_way[0];
  assign T_3242 = s2_tag_match_way[1];
  assign T_3243 = s2_tag_match_way[2];
  assign T_3244 = s2_tag_match_way[3];
  assign T_3246 = T_3241 ? T_3119_0_state : {{1'd0}, 1'h0};
  assign T_3248 = T_3242 ? T_3119_1_state : {{1'd0}, 1'h0};
  assign T_3250 = T_3243 ? T_3119_2_state : {{1'd0}, 1'h0};
  assign T_3252 = T_3244 ? T_3119_3_state : {{1'd0}, 1'h0};
  assign T_3278 = T_3246 | T_3248;
  assign T_3279 = T_3278 | T_3250;
  assign T_3280 = T_3279 | T_3252;
  assign s2_hit_state_state = T_3280;
  assign T_3331 = s2_req_cmd == 5'h1;
  assign T_3332 = s2_req_cmd == 5'h7;
  assign T_3333 = T_3331 | T_3332;
  assign T_3334 = s2_req_cmd[3];
  assign T_3335 = s2_req_cmd == 5'h4;
  assign T_3336 = T_3334 | T_3335;
  assign T_3337 = T_3333 | T_3336;
  assign T_3338 = s2_req_cmd == 5'h3;
  assign T_3339 = T_3337 | T_3338;
  assign T_3340 = s2_req_cmd == 5'h6;
  assign T_3341 = T_3339 | T_3340;
  assign T_3347_0 = 2'h2;
  assign T_3347_1 = 2'h3;
  assign T_3349 = T_3347_0 == s2_hit_state_state;
  assign T_3350 = T_3347_1 == s2_hit_state_state;
  assign T_3353 = T_3349 | T_3350;
  assign T_3359_0 = 2'h1;
  assign T_3359_1 = 2'h2;
  assign T_3359_2 = 2'h3;
  assign T_3361 = T_3359_0 == s2_hit_state_state;
  assign T_3362 = T_3359_1 == s2_hit_state_state;
  assign T_3363 = T_3359_2 == s2_hit_state_state;
  assign T_3366 = T_3361 | T_3362;
  assign T_3367 = T_3366 | T_3363;
  assign T_3368 = T_3341 ? T_3353 : T_3367;
  assign T_3369 = s2_tag_match & T_3368;
  assign T_3377 = T_3337 ? 2'h3 : s2_hit_state_state;
  assign T_3403_state = T_3377;
  assign T_3428 = s2_hit_state_state == T_3403_state;
  assign s2_hit = T_3369 & T_3428;
  assign GEN_90 = {{4'd0}, 1'h0};
  assign lrsc_valid = lrsc_count != GEN_90;
  assign T_3433 = lrsc_addr == T_2775;
  assign s2_lrsc_addr_match = lrsc_valid & T_3433;
  assign T_3435 = s2_lrsc_addr_match == 1'h0;
  assign s2_sc_fail = T_3332 & T_3435;
  assign GEN_91 = {{4'd0}, 1'h1};
  assign T_3437 = lrsc_count - GEN_91;
  assign T_3438 = T_3437[4:0];
  assign GEN_39 = lrsc_valid ? T_3438 : lrsc_count;
  assign T_3439 = s2_valid_masked & s2_hit;
  assign T_3440 = T_3439 | s2_replay;
  assign T_3442 = lrsc_valid == 1'h0;
  assign GEN_40 = T_3442 ? 5'h1f : GEN_39;
  assign GEN_41 = T_3340 ? GEN_40 : GEN_39;
  assign GEN_42 = T_3340 ? T_2775 : lrsc_addr;
  assign GEN_43 = T_3332 ? {{4'd0}, 1'h0} : GEN_41;
  assign GEN_44 = T_3440 ? GEN_43 : GEN_39;
  assign GEN_45 = T_3440 ? GEN_42 : lrsc_addr;
  assign GEN_46 = io_cpu_invalidate_lr ? {{4'd0}, 1'h0} : GEN_44;
  assign s2_data_0 = T_3460_0;
  assign s2_data_1 = T_3478_0;
  assign s2_data_2 = T_3496_0;
  assign s2_data_3 = T_3514_0;
  assign T_3463 = s1_clk_en & T_2795;
  assign T_3471 = data_io_resp_0;
  assign GEN_47 = T_3463 ? T_3471 : T_3460_0;
  assign T_3481 = s1_clk_en & T_2798;
  assign T_3489 = data_io_resp_1;
  assign GEN_48 = T_3481 ? T_3489 : T_3478_0;
  assign T_3499 = s1_clk_en & T_2801;
  assign T_3507 = data_io_resp_2;
  assign GEN_49 = T_3499 ? T_3507 : T_3496_0;
  assign T_3517 = s1_clk_en & T_2804;
  assign T_3525 = data_io_resp_3;
  assign GEN_50 = T_3517 ? T_3525 : T_3514_0;
  assign T_3531 = T_3241 ? s2_data_0 : {{63'd0}, 1'h0};
  assign T_3533 = T_3242 ? s2_data_1 : {{63'd0}, 1'h0};
  assign T_3535 = T_3243 ? s2_data_2 : {{63'd0}, 1'h0};
  assign T_3537 = T_3244 ? s2_data_3 : {{63'd0}, 1'h0};
  assign T_3539 = T_3531 | T_3533;
  assign T_3540 = T_3539 | T_3535;
  assign T_3541 = T_3540 | T_3537;
  assign s2_data_muxed = T_3541;
  assign T_3548_0 = s2_data_muxed;
  assign T_3555_0 = s2_data_muxed;
  assign T_3563_0 = 1'h0;
  assign T_3565 = T_3563_0 >> 1'h0;
  assign T_3569 = s2_sc_fail == 1'h0;
  assign T_3570 = T_3440 & T_3569;
  assign T_3578 = T_3570 & T_3337;
  assign amoalu_clk = clk;
  assign amoalu_reset = reset;
  assign amoalu_io_addr = s2_req_addr[5:0];
  assign amoalu_io_cmd = s2_req_cmd;
  assign amoalu_io_typ = s2_req_typ;
  assign amoalu_io_lhs = s2_data_word;
  assign amoalu_io_rhs = s2_req_data;
  assign T_3579 = s2_valid | s2_replay;
  assign T_3587 = T_3337 | T_3565;
  assign T_3588 = T_3579 & T_3587;
  assign T_3589 = T_3565 ? T_3548_0 : amoalu_io_out;
  assign GEN_51 = T_3588 ? s2_req_addr : s3_req_addr;
  assign GEN_52 = T_3588 ? s2_req_tag : s3_req_tag;
  assign GEN_53 = T_3588 ? s2_req_cmd : s3_req_cmd;
  assign GEN_54 = T_3588 ? s2_req_typ : s3_req_typ;
  assign GEN_55 = T_3588 ? s2_req_phys : s3_req_phys;
  assign GEN_56 = T_3588 ? T_3589 : s3_req_data;
  assign GEN_57 = T_3588 ? s2_tag_match_way : s3_way;
  assign GEN_92 = {{1'd0}, 1'h1};
  assign rowWMask = GEN_92 << 1'h0;
  assign T_3593 = T_5867;
  assign T_3597 = T_3596[0];
  assign T_3598 = T_3596[2];
  assign T_3599 = T_3597 ^ T_3598;
  assign T_3600 = T_3596[3];
  assign T_3601 = T_3599 ^ T_3600;
  assign T_3602 = T_3596[5];
  assign T_3603 = T_3601 ^ T_3602;
  assign T_3604 = T_3596[15:1];
  assign T_3605 = {T_3603,T_3604};
  assign GEN_58 = T_3593 ? T_3605 : T_3596;
  assign T_3606 = T_3596[1:0];
  assign s1_replaced_way_en = GEN_85 << T_3606;
  assign GEN_59 = s1_clk_en ? T_3606 : T_3609;
  assign s2_replaced_way_en = GEN_85 << T_3609;
  assign T_3611 = s1_replaced_way_en[0];
  assign T_3612 = s1_clk_en & T_3611;
  assign GEN_60 = T_3612 ? meta_io_resp_0_tag : T_3613_tag;
  assign GEN_61 = T_3612 ? meta_io_resp_0_coh_state : T_3613_coh_state;
  assign T_3709 = s1_replaced_way_en[1];
  assign T_3710 = s1_clk_en & T_3709;
  assign GEN_62 = T_3710 ? meta_io_resp_1_tag : T_3711_tag;
  assign GEN_63 = T_3710 ? meta_io_resp_1_coh_state : T_3711_coh_state;
  assign T_3807 = s1_replaced_way_en[2];
  assign T_3808 = s1_clk_en & T_3807;
  assign GEN_64 = T_3808 ? meta_io_resp_2_tag : T_3809_tag;
  assign GEN_65 = T_3808 ? meta_io_resp_2_coh_state : T_3809_coh_state;
  assign T_3905 = s1_replaced_way_en[3];
  assign T_3906 = s1_clk_en & T_3905;
  assign GEN_66 = T_3906 ? meta_io_resp_3_tag : T_3907_tag;
  assign GEN_67 = T_3906 ? meta_io_resp_3_coh_state : T_3907_coh_state;
  assign T_4768_0_tag = T_3613_tag;
  assign T_4768_0_coh_state = T_3613_coh_state;
  assign T_4768_1_tag = T_3711_tag;
  assign T_4768_1_coh_state = T_3711_coh_state;
  assign T_4768_2_tag = T_3809_tag;
  assign T_4768_2_coh_state = T_3809_coh_state;
  assign T_4768_3_tag = T_3907_tag;
  assign T_4768_3_coh_state = T_3907_coh_state;
  assign T_5245 = s2_replaced_way_en[0];
  assign T_5246 = s2_replaced_way_en[1];
  assign T_5247 = s2_replaced_way_en[2];
  assign T_5248 = s2_replaced_way_en[3];
  assign T_5249 = {T_4768_0_tag,T_4768_0_coh_state};
  assign T_5251 = T_5245 ? T_5249 : {{21'd0}, 1'h0};
  assign T_5252 = {T_4768_1_tag,T_4768_1_coh_state};
  assign T_5254 = T_5246 ? T_5252 : {{21'd0}, 1'h0};
  assign T_5255 = {T_4768_2_tag,T_4768_2_coh_state};
  assign T_5257 = T_5247 ? T_5255 : {{21'd0}, 1'h0};
  assign T_5258 = {T_4768_3_tag,T_4768_3_coh_state};
  assign T_5260 = T_5248 ? T_5258 : {{21'd0}, 1'h0};
  assign T_5357 = T_5251 | T_5254;
  assign T_5358 = T_5357 | T_5257;
  assign T_5359 = T_5358 | T_5260;
  assign s2_repl_meta_tag = T_5552;
  assign s2_repl_meta_coh_state = T_5551;
  assign T_5551 = T_5359[1:0];
  assign T_5552 = T_5359[21:2];
  assign T_5554 = s2_hit == 1'h0;
  assign T_5555 = s2_valid_masked & T_5554;
  assign T_5556 = s2_req_cmd == 5'h2;
  assign T_5558 = T_5556 | T_3338;
  assign T_5559 = s2_req_cmd == 5'h0;
  assign T_5561 = T_5559 | T_3340;
  assign T_5563 = T_5561 | T_3332;
  assign T_5567 = T_5563 | T_3336;
  assign T_5568 = T_5558 | T_5567;
  assign T_5576 = T_5568 | T_3337;
  assign T_5577 = T_5555 & T_5576;
  assign T_5674_tag = s2_repl_meta_tag;
  assign T_5674_coh_state = s2_hit_state_state;
  assign T_5770_tag = s2_tag_match ? T_5674_tag : s2_repl_meta_tag;
  assign T_5770_coh_state = s2_tag_match ? T_5674_coh_state : s2_repl_meta_coh_state;
  assign T_5866 = s2_tag_match ? s2_tag_match_way : s2_replaced_way_en;
  assign T_5867 = mshrs_io_req_ready & mshrs_io_req_valid;
  assign T_5871 = mshrs_io_replay_valid & readArb_io_in_1_ready;
  assign releaseArb_clk = clk;
  assign releaseArb_reset = reset;
  assign releaseArb_io_in_0_valid = wb_io_release_valid;
  assign releaseArb_io_in_0_bits_addr_beat = wb_io_release_bits_addr_beat;
  assign releaseArb_io_in_0_bits_addr_block = wb_io_release_bits_addr_block;
  assign releaseArb_io_in_0_bits_client_xact_id = wb_io_release_bits_client_xact_id;
  assign releaseArb_io_in_0_bits_voluntary = wb_io_release_bits_voluntary;
  assign releaseArb_io_in_0_bits_r_type = wb_io_release_bits_r_type;
  assign releaseArb_io_in_0_bits_data = wb_io_release_bits_data;
  assign releaseArb_io_in_1_valid = prober_io_rep_valid;
  assign releaseArb_io_in_1_bits_addr_beat = prober_io_rep_bits_addr_beat;
  assign releaseArb_io_in_1_bits_addr_block = prober_io_rep_bits_addr_block;
  assign releaseArb_io_in_1_bits_client_xact_id = prober_io_rep_bits_client_xact_id;
  assign releaseArb_io_in_1_bits_voluntary = prober_io_rep_bits_voluntary;
  assign releaseArb_io_in_1_bits_r_type = prober_io_rep_bits_r_type;
  assign releaseArb_io_in_1_bits_data = prober_io_rep_bits_data;
  assign releaseArb_io_out_ready = io_mem_release_ready;
  assign T_5904 = io_mem_probe_valid & T_3442;
  assign T_5907 = prober_io_req_ready & T_3442;
  assign FlowThroughSerializer_88_5908_clk = clk;
  assign FlowThroughSerializer_88_5908_reset = reset;
  assign FlowThroughSerializer_88_5908_io_in_valid = io_mem_grant_valid;
  assign FlowThroughSerializer_88_5908_io_in_bits_addr_beat = io_mem_grant_bits_addr_beat;
  assign FlowThroughSerializer_88_5908_io_in_bits_client_xact_id = io_mem_grant_bits_client_xact_id;
  assign FlowThroughSerializer_88_5908_io_in_bits_manager_xact_id = io_mem_grant_bits_manager_xact_id;
  assign FlowThroughSerializer_88_5908_io_in_bits_is_builtin_type = io_mem_grant_bits_is_builtin_type;
  assign FlowThroughSerializer_88_5908_io_in_bits_g_type = io_mem_grant_bits_g_type;
  assign FlowThroughSerializer_88_5908_io_in_bits_data = io_mem_grant_bits_data;
  assign FlowThroughSerializer_88_5908_io_in_bits_manager_id = io_mem_grant_bits_manager_id;
  assign FlowThroughSerializer_88_5908_io_out_ready = T_5939;
  assign T_5909 = FlowThroughSerializer_88_5908_io_out_ready & FlowThroughSerializer_88_5908_io_out_valid;
  assign T_5917_0 = 3'h5;
  assign T_5917_1 = 3'h4;
  assign GEN_95 = {{1'd0}, T_5917_0};
  assign T_5919 = GEN_95 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign GEN_96 = {{1'd0}, T_5917_1};
  assign T_5920 = GEN_96 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign T_5923 = T_5919 | T_5920;
  assign T_5929_0 = 2'h0;
  assign T_5929_1 = 2'h1;
  assign GEN_97 = {{2'd0}, T_5929_0};
  assign T_5931 = GEN_97 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign GEN_98 = {{2'd0}, T_5929_1};
  assign T_5932 = GEN_98 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign T_5935 = T_5931 | T_5932;
  assign T_5936 = FlowThroughSerializer_88_5908_io_out_bits_is_builtin_type ? T_5923 : T_5935;
  assign T_5938 = T_5936 == 1'h0;
  assign T_5939 = writeArb_io_in_1_ready | T_5938;
  assign T_5947_0 = 3'h5;
  assign T_5947_1 = 3'h4;
  assign GEN_99 = {{1'd0}, T_5947_0};
  assign T_5949 = GEN_99 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign GEN_100 = {{1'd0}, T_5947_1};
  assign T_5950 = GEN_100 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign T_5953 = T_5949 | T_5950;
  assign T_5959_0 = 2'h0;
  assign T_5959_1 = 2'h1;
  assign GEN_101 = {{2'd0}, T_5959_0};
  assign T_5961 = GEN_101 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign GEN_102 = {{2'd0}, T_5959_1};
  assign T_5962 = GEN_102 == FlowThroughSerializer_88_5908_io_out_bits_g_type;
  assign T_5965 = T_5961 | T_5962;
  assign T_5966 = FlowThroughSerializer_88_5908_io_out_bits_is_builtin_type ? T_5953 : T_5965;
  assign T_5967 = FlowThroughSerializer_88_5908_io_out_valid & T_5966;
  assign T_5969 = FlowThroughSerializer_88_5908_io_out_bits_client_xact_id < 2'h2;
  assign T_5970 = T_5967 & T_5969;
  assign T_5973 = FlowThroughSerializer_88_5908_io_out_bits_data;
  assign T_5975 = FlowThroughSerializer_88_5908_io_out_valid == 1'h0;
  assign T_5976 = T_5975 | FlowThroughSerializer_88_5908_io_out_ready;
  assign wbArb_clk = clk;
  assign wbArb_reset = reset;
  assign wbArb_io_in_0_valid = prober_io_wb_req_valid;
  assign wbArb_io_in_0_bits_addr_beat = prober_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_0_bits_addr_block = prober_io_wb_req_bits_addr_block;
  assign wbArb_io_in_0_bits_client_xact_id = prober_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_0_bits_voluntary = prober_io_wb_req_bits_voluntary;
  assign wbArb_io_in_0_bits_r_type = prober_io_wb_req_bits_r_type;
  assign wbArb_io_in_0_bits_data = prober_io_wb_req_bits_data;
  assign wbArb_io_in_0_bits_way_en = prober_io_wb_req_bits_way_en;
  assign wbArb_io_in_1_valid = mshrs_io_wb_req_valid;
  assign wbArb_io_in_1_bits_addr_beat = mshrs_io_wb_req_bits_addr_beat;
  assign wbArb_io_in_1_bits_addr_block = mshrs_io_wb_req_bits_addr_block;
  assign wbArb_io_in_1_bits_client_xact_id = mshrs_io_wb_req_bits_client_xact_id;
  assign wbArb_io_in_1_bits_voluntary = mshrs_io_wb_req_bits_voluntary;
  assign wbArb_io_in_1_bits_r_type = mshrs_io_wb_req_bits_r_type;
  assign wbArb_io_in_1_bits_data = mshrs_io_wb_req_bits_data;
  assign wbArb_io_in_1_bits_way_en = mshrs_io_wb_req_bits_way_en;
  assign wbArb_io_out_ready = wb_io_req_ready;
  assign T_6032 = s3_valid & metaReadArb_io_out_valid;
  assign GEN_69 = T_6032 ? s3_req_addr : s4_req_addr;
  assign GEN_70 = T_6032 ? s3_req_tag : s4_req_tag;
  assign GEN_71 = T_6032 ? s3_req_cmd : s4_req_cmd;
  assign GEN_72 = T_6032 ? s3_req_typ : s4_req_typ;
  assign GEN_73 = T_6032 ? s3_req_phys : s4_req_phys;
  assign GEN_74 = T_6032 ? s3_req_data : s4_req_data;
  assign T_6108 = s2_valid_masked | s2_replay;
  assign T_6111 = T_6108 & T_3569;
  assign T_6112 = s1_addr[31:3];
  assign T_6113 = s2_req_addr[39:3];
  assign GEN_103 = {{8'd0}, T_6112};
  assign T_6114 = GEN_103 == T_6113;
  assign T_6115 = T_6111 & T_6114;
  assign T_6123 = T_6115 & T_3337;
  assign T_6125 = s3_req_addr[39:3];
  assign T_6126 = GEN_103 == T_6125;
  assign T_6127 = s3_valid & T_6126;
  assign T_6128 = s3_req_cmd == 5'h1;
  assign T_6129 = s3_req_cmd == 5'h7;
  assign T_6130 = T_6128 | T_6129;
  assign T_6131 = s3_req_cmd[3];
  assign T_6132 = s3_req_cmd == 5'h4;
  assign T_6133 = T_6131 | T_6132;
  assign T_6134 = T_6130 | T_6133;
  assign T_6135 = T_6127 & T_6134;
  assign T_6137 = s4_req_addr[39:3];
  assign T_6138 = GEN_103 == T_6137;
  assign T_6139 = s4_valid & T_6138;
  assign T_6140 = s4_req_cmd == 5'h1;
  assign T_6141 = s4_req_cmd == 5'h7;
  assign T_6142 = T_6140 | T_6141;
  assign T_6143 = s4_req_cmd[3];
  assign T_6144 = s4_req_cmd == 5'h4;
  assign T_6145 = T_6143 | T_6144;
  assign T_6146 = T_6142 | T_6145;
  assign T_6147 = T_6139 & T_6146;
  assign T_6151 = T_6123 | T_6135;
  assign T_6152 = T_6151 | T_6147;
  assign T_6153 = T_6135 ? s3_req_data : s4_req_data;
  assign T_6154 = T_6123 ? amoalu_io_out : T_6153;
  assign GEN_75 = T_6152 ? T_6154 : s2_store_bypass_data;
  assign GEN_77 = s1_clk_en ? T_6152 : s2_store_bypass;
  assign GEN_78 = s1_clk_en ? GEN_75 : s2_store_bypass_data;
  assign s2_data_word_prebypass = T_3555_0 >> 7'h0;
  assign s2_data_word = s2_store_bypass ? s2_store_bypass_data : s2_data_word_prebypass;
  assign T_6158 = s2_req_typ[1:0];
  assign T_6159 = $signed(s2_req_typ);
  assign GEN_106 = $signed(1'h0);
  assign GEN_107 = {3{GEN_106}};
  assign T_6161 = $signed(T_6159) >= $signed(GEN_107);
  assign T_6162 = dtlb_io_req_valid & dtlb_io_resp_miss;
  assign T_6163 = s1_req_addr[11:6];
  assign T_6164 = T_6163 == prober_io_meta_write_bits_idx;
  assign T_6166 = prober_io_req_ready == 1'h0;
  assign T_6167 = T_6164 & T_6166;
  assign s1_nack = T_6162 | T_6167;
  assign T_6168 = s1_valid | s1_replay;
  assign GEN_79 = T_6168 ? s1_nack : s2_nack_hit;
  assign GEN_80 = s2_nack_hit ? 1'h0 : T_5577;
  assign s2_nack_victim = s2_hit & mshrs_io_secondary_miss;
  assign T_6173 = mshrs_io_req_ready == 1'h0;
  assign s2_nack_miss = T_5554 & T_6173;
  assign T_6174 = s2_nack_hit | s2_nack_victim;
  assign s2_nack = T_6174 | s2_nack_miss;
  assign T_6176 = s2_nack == 1'h0;
  assign T_6177 = s2_valid & T_6176;
  assign T_6179 = T_3579 & s2_hit;
  assign s2_recycle_ecc = T_6179 & T_3565;
  assign GEN_81 = T_6168 ? s2_recycle_ecc : s2_recycle_next;
  assign T_6182 = s2_recycle_ecc | s2_recycle_next;
  assign T_6184 = s2_valid | block_miss;
  assign T_6185 = T_6184 & s2_nack_miss;
  assign GEN_82 = block_miss ? 1'h0 : GEN_33;
  assign cache_resp_valid = T_6589;
  assign cache_resp_bits_addr = s2_req_addr;
  assign cache_resp_bits_tag = s2_req_tag;
  assign cache_resp_bits_cmd = s2_req_cmd;
  assign cache_resp_bits_typ = s2_req_typ;
  assign cache_resp_bits_data = T_6656;
  assign cache_resp_bits_replay = s2_replay;
  assign cache_resp_bits_has_data = T_5567;
  assign cache_resp_bits_data_word_bypass = GEN_93;
  assign cache_resp_bits_store_data = s2_req_data;
  assign T_6586 = s2_replay | T_3439;
  assign T_6588 = T_3565 == 1'h0;
  assign T_6589 = T_6586 & T_6588;
  assign T_6599 = s2_req_addr[2];
  assign T_6600 = s2_data_word[63:32];
  assign T_6601 = s2_data_word[31:0];
  assign T_6602 = T_6599 ? T_6600 : T_6601;
  assign T_6608 = T_6158 == 2'h2;
  assign T_6610 = T_6602[31];
  assign T_6611 = T_6161 & T_6610;
  assign GEN_108 = {{31'd0}, T_6611};
  assign T_6613 = 32'h0 - GEN_108;
  assign T_6614 = T_6613[31:0];
  assign T_6616 = T_6608 ? T_6614 : T_6600;
  assign T_6617 = {T_6616,T_6602};
  assign T_6618 = s2_req_addr[1];
  assign T_6619 = T_6617[31:16];
  assign T_6620 = T_6617[15:0];
  assign T_6621 = T_6618 ? T_6619 : T_6620;
  assign T_6627 = T_6158 == GEN_92;
  assign T_6629 = T_6621[15];
  assign T_6630 = T_6161 & T_6629;
  assign GEN_110 = {{47'd0}, T_6630};
  assign T_6632 = 48'h0 - GEN_110;
  assign T_6633 = T_6632[47:0];
  assign T_6634 = T_6617[63:16];
  assign T_6635 = T_6627 ? T_6633 : T_6634;
  assign T_6636 = {T_6635,T_6621};
  assign T_6637 = s2_req_addr[0];
  assign T_6638 = T_6636[15:8];
  assign T_6639 = T_6636[7:0];
  assign T_6640 = T_6637 ? T_6638 : T_6639;
  assign T_6644 = T_3332 ? {{7'd0}, 1'h0} : T_6640;
  assign GEN_111 = {{1'd0}, 1'h0};
  assign T_6646 = T_6158 == GEN_111;
  assign T_6647 = T_6646 | T_3332;
  assign T_6648 = T_6644[7];
  assign T_6649 = T_6161 & T_6648;
  assign GEN_112 = {{55'd0}, T_6649};
  assign T_6651 = 56'h0 - GEN_112;
  assign T_6652 = T_6651[55:0];
  assign T_6653 = T_6636[63:8];
  assign T_6654 = T_6647 ? T_6652 : T_6653;
  assign T_6655 = {T_6654,T_6644};
  assign GEN_113 = {{63'd0}, s2_sc_fail};
  assign T_6656 = T_6655 | GEN_113;
  assign uncache_resp_valid = mshrs_io_resp_valid;
  assign uncache_resp_bits_addr = mshrs_io_resp_bits_addr;
  assign uncache_resp_bits_tag = mshrs_io_resp_bits_tag;
  assign uncache_resp_bits_cmd = mshrs_io_resp_bits_cmd;
  assign uncache_resp_bits_typ = mshrs_io_resp_bits_typ;
  assign uncache_resp_bits_data = mshrs_io_resp_bits_data;
  assign uncache_resp_bits_replay = mshrs_io_resp_bits_replay;
  assign uncache_resp_bits_has_data = mshrs_io_resp_bits_has_data;
  assign uncache_resp_bits_data_word_bypass = mshrs_io_resp_bits_data_word_bypass;
  assign uncache_resp_bits_store_data = mshrs_io_resp_bits_store_data;
  assign T_7057 = T_6168 == 1'h0;
  assign T_7059 = s2_valid & s2_nack;
  assign T_7060_valid = mshrs_io_resp_ready ? uncache_resp_valid : cache_resp_valid;
  assign T_7060_bits_addr = mshrs_io_resp_ready ? uncache_resp_bits_addr : cache_resp_bits_addr;
  assign T_7060_bits_tag = mshrs_io_resp_ready ? uncache_resp_bits_tag : cache_resp_bits_tag;
  assign T_7060_bits_cmd = mshrs_io_resp_ready ? uncache_resp_bits_cmd : cache_resp_bits_cmd;
  assign T_7060_bits_typ = mshrs_io_resp_ready ? uncache_resp_bits_typ : cache_resp_bits_typ;
  assign T_7060_bits_data = mshrs_io_resp_ready ? uncache_resp_bits_data : cache_resp_bits_data;
  assign T_7060_bits_replay = mshrs_io_resp_ready ? uncache_resp_bits_replay : cache_resp_bits_replay;
  assign T_7060_bits_has_data = mshrs_io_resp_ready ? uncache_resp_bits_has_data : cache_resp_bits_has_data;
  assign T_7060_bits_store_data = mshrs_io_resp_ready ? uncache_resp_bits_store_data : cache_resp_bits_store_data;
  assign T_7241 = mshrs_io_fence_rdy & T_2817;
  assign T_7243 = s2_valid == 1'h0;
  assign T_7244 = T_7241 & T_7243;
  assign T_7245 = s1_replay & s1_read;
  assign T_7246 = T_7245 | mshrs_io_replay_next;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_94 = {1{$random}};
  s1_valid = GEN_94[0:0];
  GEN_104 = {2{$random}};
  s1_req_addr = GEN_104[39:0];
  GEN_105 = {1{$random}};
  s1_req_tag = GEN_105[8:0];
  GEN_109 = {1{$random}};
  s1_req_cmd = GEN_109[4:0];
  GEN_114 = {1{$random}};
  s1_req_typ = GEN_114[2:0];
  GEN_115 = {1{$random}};
  s1_req_phys = GEN_115[0:0];
  GEN_116 = {2{$random}};
  s1_req_data = GEN_116[63:0];
  GEN_117 = {1{$random}};
  s1_replay = GEN_117[0:0];
  GEN_118 = {1{$random}};
  s1_clk_en = GEN_118[0:0];
  GEN_119 = {1{$random}};
  s2_valid = GEN_119[0:0];
  GEN_120 = {2{$random}};
  s2_req_addr = GEN_120[39:0];
  GEN_121 = {1{$random}};
  s2_req_tag = GEN_121[8:0];
  GEN_122 = {1{$random}};
  s2_req_cmd = GEN_122[4:0];
  GEN_123 = {1{$random}};
  s2_req_typ = GEN_123[2:0];
  GEN_124 = {1{$random}};
  s2_req_phys = GEN_124[0:0];
  GEN_125 = {2{$random}};
  s2_req_data = GEN_125[63:0];
  GEN_126 = {1{$random}};
  T_2233 = GEN_126[0:0];
  GEN_127 = {1{$random}};
  s3_valid = GEN_127[0:0];
  GEN_128 = {2{$random}};
  s3_req_addr = GEN_128[39:0];
  GEN_129 = {1{$random}};
  s3_req_tag = GEN_129[8:0];
  GEN_130 = {1{$random}};
  s3_req_cmd = GEN_130[4:0];
  GEN_131 = {1{$random}};
  s3_req_typ = GEN_131[2:0];
  GEN_132 = {1{$random}};
  s3_req_phys = GEN_132[0:0];
  GEN_133 = {2{$random}};
  s3_req_data = GEN_133[63:0];
  GEN_134 = {1{$random}};
  s3_way = GEN_134[3:0];
  GEN_135 = {1{$random}};
  s1_recycled = GEN_135[0:0];
  GEN_136 = {1{$random}};
  T_2368 = GEN_136[0:0];
  GEN_137 = {1{$random}};
  s2_tag_match_way = GEN_137[3:0];
  GEN_138 = {1{$random}};
  T_2822_state = GEN_138[1:0];
  GEN_139 = {1{$random}};
  T_2847_state = GEN_139[1:0];
  GEN_140 = {1{$random}};
  T_2872_state = GEN_140[1:0];
  GEN_141 = {1{$random}};
  T_2897_state = GEN_141[1:0];
  GEN_142 = {1{$random}};
  lrsc_count = GEN_142[4:0];
  GEN_143 = {2{$random}};
  lrsc_addr = GEN_143[33:0];
  GEN_144 = {2{$random}};
  T_3460_0 = GEN_144[63:0];
  GEN_145 = {2{$random}};
  T_3478_0 = GEN_145[63:0];
  GEN_146 = {2{$random}};
  T_3496_0 = GEN_146[63:0];
  GEN_147 = {2{$random}};
  T_3514_0 = GEN_147[63:0];
  GEN_148 = {1{$random}};
  T_3596 = GEN_148[15:0];
  GEN_149 = {1{$random}};
  T_3609 = GEN_149[1:0];
  GEN_150 = {1{$random}};
  T_3613_tag = GEN_150[19:0];
  GEN_151 = {1{$random}};
  T_3613_coh_state = GEN_151[1:0];
  GEN_152 = {1{$random}};
  T_3711_tag = GEN_152[19:0];
  GEN_153 = {1{$random}};
  T_3711_coh_state = GEN_153[1:0];
  GEN_154 = {1{$random}};
  T_3809_tag = GEN_154[19:0];
  GEN_155 = {1{$random}};
  T_3809_coh_state = GEN_155[1:0];
  GEN_156 = {1{$random}};
  T_3907_tag = GEN_156[19:0];
  GEN_157 = {1{$random}};
  T_3907_coh_state = GEN_157[1:0];
  GEN_158 = {1{$random}};
  s4_valid = GEN_158[0:0];
  GEN_159 = {2{$random}};
  s4_req_addr = GEN_159[39:0];
  GEN_160 = {1{$random}};
  s4_req_tag = GEN_160[8:0];
  GEN_161 = {1{$random}};
  s4_req_cmd = GEN_161[4:0];
  GEN_162 = {1{$random}};
  s4_req_typ = GEN_162[2:0];
  GEN_163 = {1{$random}};
  s4_req_phys = GEN_163[0:0];
  GEN_164 = {2{$random}};
  s4_req_data = GEN_164[63:0];
  GEN_165 = {2{$random}};
  s2_store_bypass_data = GEN_165[63:0];
  GEN_166 = {1{$random}};
  s2_store_bypass = GEN_166[0:0];
  GEN_167 = {1{$random}};
  s2_nack_hit = GEN_167[0:0];
  GEN_168 = {1{$random}};
  s2_recycle_next = GEN_168[0:0];
  GEN_169 = {1{$random}};
  block_miss = GEN_169[0:0];
  GEN_170 = {1{$random}};
  T_7058 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  GEN_68 = GEN_171[1:0];
  GEN_172 = {1{$random}};
  GEN_76 = GEN_172[3:0];
  GEN_173 = {1{$random}};
  GEN_86 = GEN_173[3:0];
  GEN_174 = {2{$random}};
  GEN_93 = GEN_174[63:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      s1_valid <= 1'h0;
    end else begin
      s1_valid <= T_2075;
    end
    if(1'h0) begin
    end else begin
      s1_req_addr <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      s1_req_tag <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      s1_req_cmd <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      s1_req_typ <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      s1_req_phys <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      s1_req_data <= GEN_23;
    end
    if(reset) begin
      s1_replay <= 1'h0;
    end else begin
      s1_replay <= T_5871;
    end
    if(1'h0) begin
    end else begin
      s1_clk_en <= metaReadArb_io_out_valid;
    end
    if(reset) begin
      s2_valid <= 1'h0;
    end else begin
      s2_valid <= s1_valid_masked;
    end
    if(1'h0) begin
    end else begin
      s2_req_addr <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      s2_req_tag <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      s2_req_cmd <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      s2_req_typ <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      s2_req_phys <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      s2_req_data <= GEN_29;
    end
    if(reset) begin
      T_2233 <= 1'h0;
    end else begin
      T_2233 <= s1_replay;
    end
    if(reset) begin
      s3_valid <= 1'h0;
    end else begin
      s3_valid <= T_3578;
    end
    if(1'h0) begin
    end else begin
      s3_req_addr <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      s3_req_tag <= GEN_52;
    end
    if(1'h0) begin
    end else begin
      s3_req_cmd <= GEN_53;
    end
    if(1'h0) begin
    end else begin
      s3_req_typ <= GEN_54;
    end
    if(1'h0) begin
    end else begin
      s3_req_phys <= GEN_55;
    end
    if(1'h0) begin
    end else begin
      s3_req_data <= GEN_56;
    end
    if(1'h0) begin
    end else begin
      s3_way <= GEN_57;
    end
    if(reset) begin
      s1_recycled <= 1'h0;
    end else begin
      s1_recycled <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      T_2368 <= T_2367;
    end
    if(1'h0) begin
    end else begin
      s2_tag_match_way <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      T_2822_state <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      T_2847_state <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      T_2872_state <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      T_2897_state <= GEN_38;
    end
    if(reset) begin
      lrsc_count <= {{4'd0}, 1'h0};
    end else begin
      lrsc_count <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      lrsc_addr <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      T_3460_0 <= GEN_47;
    end
    if(1'h0) begin
    end else begin
      T_3478_0 <= GEN_48;
    end
    if(1'h0) begin
    end else begin
      T_3496_0 <= GEN_49;
    end
    if(1'h0) begin
    end else begin
      T_3514_0 <= GEN_50;
    end
    if(reset) begin
      T_3596 <= 16'h1;
    end else begin
      T_3596 <= GEN_58;
    end
    if(1'h0) begin
    end else begin
      T_3609 <= GEN_59;
    end
    if(1'h0) begin
    end else begin
      T_3613_tag <= GEN_60;
    end
    if(1'h0) begin
    end else begin
      T_3613_coh_state <= GEN_61;
    end
    if(1'h0) begin
    end else begin
      T_3711_tag <= GEN_62;
    end
    if(1'h0) begin
    end else begin
      T_3711_coh_state <= GEN_63;
    end
    if(1'h0) begin
    end else begin
      T_3809_tag <= GEN_64;
    end
    if(1'h0) begin
    end else begin
      T_3809_coh_state <= GEN_65;
    end
    if(1'h0) begin
    end else begin
      T_3907_tag <= GEN_66;
    end
    if(1'h0) begin
    end else begin
      T_3907_coh_state <= GEN_67;
    end
    if(reset) begin
      s4_valid <= 1'h0;
    end else begin
      s4_valid <= s3_valid;
    end
    if(1'h0) begin
    end else begin
      s4_req_addr <= GEN_69;
    end
    if(1'h0) begin
    end else begin
      s4_req_tag <= GEN_70;
    end
    if(1'h0) begin
    end else begin
      s4_req_cmd <= GEN_71;
    end
    if(1'h0) begin
    end else begin
      s4_req_typ <= GEN_72;
    end
    if(1'h0) begin
    end else begin
      s4_req_phys <= GEN_73;
    end
    if(1'h0) begin
    end else begin
      s4_req_data <= GEN_74;
    end
    if(1'h0) begin
    end else begin
      s2_store_bypass_data <= GEN_78;
    end
    if(1'h0) begin
    end else begin
      s2_store_bypass <= GEN_77;
    end
    if(1'h0) begin
    end else begin
      s2_nack_hit <= GEN_79;
    end
    if(reset) begin
      s2_recycle_next <= 1'h0;
    end else begin
      s2_recycle_next <= GEN_81;
    end
    if(reset) begin
      block_miss <= 1'h0;
    end else begin
      block_miss <= T_6185;
    end
    if(1'h0) begin
    end else begin
      T_7058 <= T_7057;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2374) begin
          $fwrite(32'h80000002,"Assertion failed: DCache exception occurred - cache response not killed.\n    at nbdcache.scala:863 assert (!(Reg(next=\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_2374) begin
          $fdisplay(32'h80000002,"1");$finish;
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
  end
endmodule
module FPUDecoder(
  input   clk,
  input   reset,
  input  [31:0] io_inst,
  output [4:0] io_sigs_cmd,
  output  io_sigs_ldst,
  output  io_sigs_wen,
  output  io_sigs_ren1,
  output  io_sigs_ren2,
  output  io_sigs_ren3,
  output  io_sigs_swap12,
  output  io_sigs_swap23,
  output  io_sigs_single,
  output  io_sigs_fromint,
  output  io_sigs_toint,
  output  io_sigs_fastpipe,
  output  io_sigs_fma,
  output  io_sigs_div,
  output  io_sigs_sqrt,
  output  io_sigs_round,
  output  io_sigs_wflags
);
  wire [31:0] T_37;
  wire  T_39;
  wire [31:0] T_41;
  wire  T_43;
  wire  T_46;
  wire [31:0] T_48;
  wire  T_50;
  wire [31:0] T_52;
  wire  T_54;
  wire  T_57;
  wire [31:0] T_59;
  wire  T_61;
  wire [31:0] T_63;
  wire  T_65;
  wire  T_68;
  wire [31:0] T_70;
  wire  T_72;
  wire  T_75;
  wire [31:0] T_77;
  wire  T_79;
  wire [1:0] T_82;
  wire [2:0] T_83;
  wire [3:0] T_84;
  wire [4:0] T_85;
  wire [31:0] T_89;
  wire  T_91;
  wire [31:0] T_93;
  wire  T_95;
  wire [31:0] T_97;
  wire  T_99;
  wire  T_102;
  wire  T_103;
  wire [31:0] T_105;
  wire  T_107;
  wire [31:0] T_109;
  wire  T_111;
  wire [31:0] T_113;
  wire  T_115;
  wire  T_118;
  wire  T_119;
  wire [31:0] T_121;
  wire  T_123;
  wire [31:0] T_125;
  wire  T_127;
  wire  T_130;
  wire  T_131;
  wire [31:0] T_135;
  wire  T_137;
  wire  T_140;
  wire [31:0] T_142;
  wire  T_144;
  wire [31:0] T_148;
  wire  T_150;
  wire [31:0] T_152;
  wire  T_154;
  wire  T_157;
  wire [31:0] T_159;
  wire  T_161;
  wire  T_167;
  wire  T_170;
  wire [31:0] T_172;
  wire  T_174;
  wire [31:0] T_176;
  wire  T_178;
  wire  T_181;
  wire [31:0] T_183;
  wire  T_185;
  wire [31:0] T_187;
  wire  T_189;
  wire  T_192;
  wire  T_193;
  wire [31:0] T_195;
  wire  T_197;
  wire  T_203;
  wire [31:0] T_207;
  wire  T_209;
  wire [31:0] T_211;
  wire  T_213;
  wire  T_216;
  wire  T_217;
  wire [31:0] T_219;
  wire  T_221;
  wire [31:0] T_223;
  wire  T_225;
  wire  T_229;
  wire  T_230;
  assign io_sigs_cmd = T_85;
  assign io_sigs_ldst = T_61;
  assign io_sigs_wen = T_103;
  assign io_sigs_ren1 = T_119;
  assign io_sigs_ren2 = T_131;
  assign io_sigs_ren3 = T_115;
  assign io_sigs_swap12 = T_140;
  assign io_sigs_swap23 = T_144;
  assign io_sigs_single = T_157;
  assign io_sigs_fromint = T_161;
  assign io_sigs_toint = T_170;
  assign io_sigs_fastpipe = T_181;
  assign io_sigs_fma = T_193;
  assign io_sigs_div = T_197;
  assign io_sigs_sqrt = T_203;
  assign io_sigs_round = T_217;
  assign io_sigs_wflags = T_230;
  assign T_37 = io_inst & 32'h4;
  assign T_39 = T_37 == 32'h4;
  assign T_41 = io_inst & 32'h8000010;
  assign T_43 = T_41 == 32'h8000010;
  assign T_46 = T_39 | T_43;
  assign T_48 = io_inst & 32'h8;
  assign T_50 = T_48 == 32'h8;
  assign T_52 = io_inst & 32'h10000010;
  assign T_54 = T_52 == 32'h10000010;
  assign T_57 = T_50 | T_54;
  assign T_59 = io_inst & 32'h40;
  assign T_61 = T_59 == 32'h0;
  assign T_63 = io_inst & 32'h20000000;
  assign T_65 = T_63 == 32'h20000000;
  assign T_68 = T_61 | T_65;
  assign T_70 = io_inst & 32'h40000000;
  assign T_72 = T_70 == 32'h40000000;
  assign T_75 = T_61 | T_72;
  assign T_77 = io_inst & 32'h10;
  assign T_79 = T_77 == 32'h0;
  assign T_82 = {T_57,T_46};
  assign T_83 = {T_68,T_82};
  assign T_84 = {T_75,T_83};
  assign T_85 = {T_79,T_84};
  assign T_89 = io_inst & 32'h80000020;
  assign T_91 = T_89 == 32'h0;
  assign T_93 = io_inst & 32'h30;
  assign T_95 = T_93 == 32'h0;
  assign T_97 = io_inst & 32'h10000020;
  assign T_99 = T_97 == 32'h10000000;
  assign T_102 = T_91 | T_95;
  assign T_103 = T_102 | T_99;
  assign T_105 = io_inst & 32'h80000004;
  assign T_107 = T_105 == 32'h0;
  assign T_109 = io_inst & 32'h10000004;
  assign T_111 = T_109 == 32'h0;
  assign T_113 = io_inst & 32'h50;
  assign T_115 = T_113 == 32'h40;
  assign T_118 = T_107 | T_111;
  assign T_119 = T_118 | T_115;
  assign T_121 = io_inst & 32'h40000004;
  assign T_123 = T_121 == 32'h0;
  assign T_125 = io_inst & 32'h20;
  assign T_127 = T_125 == 32'h20;
  assign T_130 = T_123 | T_127;
  assign T_131 = T_130 | T_115;
  assign T_135 = io_inst & 32'h50000010;
  assign T_137 = T_135 == 32'h50000010;
  assign T_140 = T_61 | T_137;
  assign T_142 = io_inst & 32'h30000010;
  assign T_144 = T_142 == 32'h10;
  assign T_148 = io_inst & 32'h1040;
  assign T_150 = T_148 == 32'h0;
  assign T_152 = io_inst & 32'h2000040;
  assign T_154 = T_152 == 32'h40;
  assign T_157 = T_150 | T_154;
  assign T_159 = io_inst & 32'h90000010;
  assign T_161 = T_159 == 32'h90000010;
  assign T_167 = T_159 == 32'h80000010;
  assign T_170 = T_127 | T_167;
  assign T_172 = io_inst & 32'ha0000010;
  assign T_174 = T_172 == 32'h20000010;
  assign T_176 = io_inst & 32'hd0000010;
  assign T_178 = T_176 == 32'h40000010;
  assign T_181 = T_174 | T_178;
  assign T_183 = io_inst & 32'h70000004;
  assign T_185 = T_183 == 32'h0;
  assign T_187 = io_inst & 32'h68000004;
  assign T_189 = T_187 == 32'h0;
  assign T_192 = T_185 | T_189;
  assign T_193 = T_192 | T_115;
  assign T_195 = io_inst & 32'h58000010;
  assign T_197 = T_195 == 32'h18000010;
  assign T_203 = T_176 == 32'h50000010;
  assign T_207 = io_inst & 32'h20000004;
  assign T_209 = T_207 == 32'h0;
  assign T_211 = io_inst & 32'h40002000;
  assign T_213 = T_211 == 32'h40000000;
  assign T_216 = T_209 | T_115;
  assign T_217 = T_216 | T_213;
  assign T_219 = io_inst & 32'h8002000;
  assign T_221 = T_219 == 32'h8000000;
  assign T_223 = io_inst & 32'hc0000004;
  assign T_225 = T_223 == 32'h80000000;
  assign T_229 = T_216 | T_221;
  assign T_230 = T_229 | T_225;
endmodule
module MulAddRecFN_preMul(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [1:0] io_roundingMode,
  output [23:0] io_mulAddA,
  output [23:0] io_mulAddB,
  output [47:0] io_mulAddC,
  output [2:0] io_toPostMul_highExpA,
  output  io_toPostMul_isNaN_isQuietNaNA,
  output [2:0] io_toPostMul_highExpB,
  output  io_toPostMul_isNaN_isQuietNaNB,
  output  io_toPostMul_signProd,
  output  io_toPostMul_isZeroProd,
  output  io_toPostMul_opSignC,
  output [2:0] io_toPostMul_highExpC,
  output  io_toPostMul_isNaN_isQuietNaNC,
  output  io_toPostMul_isCDominant,
  output  io_toPostMul_CAlignDist_0,
  output [6:0] io_toPostMul_CAlignDist,
  output  io_toPostMul_bit0AlignedNegSigC,
  output [25:0] io_toPostMul_highAlignedNegSigC,
  output [10:0] io_toPostMul_sExpSum,
  output [1:0] io_toPostMul_roundingMode
);
  wire  signA;
  wire [8:0] expA;
  wire [22:0] fractA;
  wire [2:0] T_42;
  wire [2:0] GEN_0;
  wire  isZeroA;
  wire  T_45;
  wire [23:0] sigA;
  wire  signB;
  wire [8:0] expB;
  wire [22:0] fractB;
  wire [2:0] T_46;
  wire  isZeroB;
  wire  T_49;
  wire [23:0] sigB;
  wire  T_50;
  wire  T_51;
  wire  opSignC;
  wire [8:0] expC;
  wire [22:0] fractC;
  wire [2:0] T_52;
  wire  isZeroC;
  wire  T_55;
  wire [23:0] sigC;
  wire  T_56;
  wire  T_57;
  wire  signProd;
  wire  isZeroProd;
  wire  T_58;
  wire  T_60;
  wire [2:0] GEN_3;
  wire [3:0] T_62;
  wire [2:0] T_63;
  wire [7:0] T_64;
  wire [10:0] T_65;
  wire [10:0] GEN_4;
  wire [11:0] T_66;
  wire [10:0] T_67;
  wire [10:0] GEN_5;
  wire [11:0] T_69;
  wire [10:0] sExpAlignedProd;
  wire  doSubMags;
  wire [10:0] GEN_6;
  wire [11:0] T_70;
  wire [10:0] sNatCAlignDist;
  wire  T_71;
  wire  CAlignDist_floor;
  wire [9:0] T_72;
  wire [9:0] GEN_7;
  wire  T_74;
  wire  CAlignDist_0;
  wire [9:0] GEN_8;
  wire  T_79;
  wire  T_80;
  wire  isCDominant;
  wire [9:0] GEN_9;
  wire  T_84;
  wire [6:0] T_85;
  wire [6:0] T_87;
  wire [6:0] CAlignDist;
  wire [10:0] sExpSum;
  wire [128:0] GEN_10;
  wire [128:0] T_89;
  wire [23:0] T_90;
  wire [15:0] T_91;
  wire [7:0] T_96;
  wire [15:0] GEN_11;
  wire [15:0] T_97;
  wire [7:0] T_98;
  wire [15:0] GEN_12;
  wire [15:0] T_99;
  wire [15:0] T_101;
  wire [15:0] T_102;
  wire [11:0] T_106;
  wire [15:0] GEN_13;
  wire [15:0] T_107;
  wire [11:0] T_108;
  wire [15:0] GEN_14;
  wire [15:0] T_109;
  wire [15:0] T_111;
  wire [15:0] T_112;
  wire [13:0] T_116;
  wire [15:0] GEN_15;
  wire [15:0] T_117;
  wire [13:0] T_118;
  wire [15:0] GEN_16;
  wire [15:0] T_119;
  wire [15:0] T_121;
  wire [15:0] T_122;
  wire [14:0] T_126;
  wire [15:0] GEN_17;
  wire [15:0] T_127;
  wire [14:0] T_128;
  wire [15:0] GEN_18;
  wire [15:0] T_129;
  wire [15:0] T_131;
  wire [15:0] T_132;
  wire [7:0] T_133;
  wire [3:0] T_138;
  wire [7:0] GEN_19;
  wire [7:0] T_139;
  wire [3:0] T_140;
  wire [7:0] GEN_20;
  wire [7:0] T_141;
  wire [7:0] T_143;
  wire [7:0] T_144;
  wire [5:0] T_148;
  wire [7:0] GEN_21;
  wire [7:0] T_149;
  wire [5:0] T_150;
  wire [7:0] GEN_22;
  wire [7:0] T_151;
  wire [7:0] T_153;
  wire [7:0] T_154;
  wire [6:0] T_158;
  wire [7:0] GEN_23;
  wire [7:0] T_159;
  wire [6:0] T_160;
  wire [7:0] GEN_24;
  wire [7:0] T_161;
  wire [7:0] T_163;
  wire [7:0] T_164;
  wire [23:0] CExtraMask;
  wire [23:0] T_165;
  wire [23:0] negSigC;
  wire [49:0] GEN_25;
  wire [50:0] T_167;
  wire [49:0] T_168;
  wire [24:0] T_169;
  wire [74:0] T_170;
  wire [74:0] T_171;
  wire [74:0] T_172;
  wire [23:0] T_173;
  wire [23:0] GEN_26;
  wire  T_175;
  wire  T_176;
  wire [74:0] T_177;
  wire [75:0] T_178;
  wire [74:0] alignedNegSigC;
  wire [47:0] T_179;
  wire  T_181;
  wire  T_183;
  wire  T_185;
  wire  T_186;
  wire [25:0] T_187;
  assign io_mulAddA = sigA;
  assign io_mulAddB = sigB;
  assign io_mulAddC = T_179;
  assign io_toPostMul_highExpA = T_42;
  assign io_toPostMul_isNaN_isQuietNaNA = T_181;
  assign io_toPostMul_highExpB = T_46;
  assign io_toPostMul_isNaN_isQuietNaNB = T_183;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_highExpC = T_52;
  assign io_toPostMul_isNaN_isQuietNaNC = T_185;
  assign io_toPostMul_isCDominant = isCDominant;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_bit0AlignedNegSigC = T_186;
  assign io_toPostMul_highAlignedNegSigC = T_187;
  assign io_toPostMul_sExpSum = sExpSum;
  assign io_toPostMul_roundingMode = io_roundingMode;
  assign signA = io_a[32];
  assign expA = io_a[31:23];
  assign fractA = io_a[22:0];
  assign T_42 = expA[8:6];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZeroA = T_42 == GEN_0;
  assign T_45 = isZeroA == 1'h0;
  assign sigA = {T_45,fractA};
  assign signB = io_b[32];
  assign expB = io_b[31:23];
  assign fractB = io_b[22:0];
  assign T_46 = expB[8:6];
  assign isZeroB = T_46 == GEN_0;
  assign T_49 = isZeroB == 1'h0;
  assign sigB = {T_49,fractB};
  assign T_50 = io_c[32];
  assign T_51 = io_op[0];
  assign opSignC = T_50 ^ T_51;
  assign expC = io_c[31:23];
  assign fractC = io_c[22:0];
  assign T_52 = expC[8:6];
  assign isZeroC = T_52 == GEN_0;
  assign T_55 = isZeroC == 1'h0;
  assign sigC = {T_55,fractC};
  assign T_56 = signA ^ signB;
  assign T_57 = io_op[1];
  assign signProd = T_56 ^ T_57;
  assign isZeroProd = isZeroA | isZeroB;
  assign T_58 = expB[8];
  assign T_60 = T_58 == 1'h0;
  assign GEN_3 = {{2'd0}, T_60};
  assign T_62 = 3'h0 - GEN_3;
  assign T_63 = T_62[2:0];
  assign T_64 = expB[7:0];
  assign T_65 = {T_63,T_64};
  assign GEN_4 = {{2'd0}, expA};
  assign T_66 = GEN_4 + T_65;
  assign T_67 = T_66[10:0];
  assign GEN_5 = {{6'd0}, 5'h1b};
  assign T_69 = T_67 + GEN_5;
  assign sExpAlignedProd = T_69[10:0];
  assign doSubMags = signProd ^ opSignC;
  assign GEN_6 = {{2'd0}, expC};
  assign T_70 = sExpAlignedProd - GEN_6;
  assign sNatCAlignDist = T_70[10:0];
  assign T_71 = sNatCAlignDist[10];
  assign CAlignDist_floor = isZeroProd | T_71;
  assign T_72 = sNatCAlignDist[9:0];
  assign GEN_7 = {{9'd0}, 1'h0};
  assign T_74 = T_72 == GEN_7;
  assign CAlignDist_0 = CAlignDist_floor | T_74;
  assign GEN_8 = {{5'd0}, 5'h19};
  assign T_79 = T_72 < GEN_8;
  assign T_80 = CAlignDist_floor | T_79;
  assign isCDominant = T_55 & T_80;
  assign GEN_9 = {{3'd0}, 7'h4a};
  assign T_84 = T_72 < GEN_9;
  assign T_85 = sNatCAlignDist[6:0];
  assign T_87 = T_84 ? T_85 : 7'h4a;
  assign CAlignDist = CAlignDist_floor ? {{6'd0}, 1'h0} : T_87;
  assign sExpSum = CAlignDist_floor ? {{2'd0}, expC} : sExpAlignedProd;
  assign GEN_10 = $signed(129'h100000000000000000000000000000000);
  assign T_89 = $signed(GEN_10) >>> CAlignDist;
  assign T_90 = T_89[77:54];
  assign T_91 = T_90[15:0];
  assign T_96 = T_91[15:8];
  assign GEN_11 = {{8'd0}, T_96};
  assign T_97 = GEN_11 & 16'hff;
  assign T_98 = T_91[7:0];
  assign GEN_12 = {{8'd0}, T_98};
  assign T_99 = GEN_12 << 8;
  assign T_101 = T_99 & 16'hff00;
  assign T_102 = T_97 | T_101;
  assign T_106 = T_102[15:4];
  assign GEN_13 = {{4'd0}, T_106};
  assign T_107 = GEN_13 & 16'hf0f;
  assign T_108 = T_102[11:0];
  assign GEN_14 = {{4'd0}, T_108};
  assign T_109 = GEN_14 << 4;
  assign T_111 = T_109 & 16'hf0f0;
  assign T_112 = T_107 | T_111;
  assign T_116 = T_112[15:2];
  assign GEN_15 = {{2'd0}, T_116};
  assign T_117 = GEN_15 & 16'h3333;
  assign T_118 = T_112[13:0];
  assign GEN_16 = {{2'd0}, T_118};
  assign T_119 = GEN_16 << 2;
  assign T_121 = T_119 & 16'hcccc;
  assign T_122 = T_117 | T_121;
  assign T_126 = T_122[15:1];
  assign GEN_17 = {{1'd0}, T_126};
  assign T_127 = GEN_17 & 16'h5555;
  assign T_128 = T_122[14:0];
  assign GEN_18 = {{1'd0}, T_128};
  assign T_129 = GEN_18 << 1;
  assign T_131 = T_129 & 16'haaaa;
  assign T_132 = T_127 | T_131;
  assign T_133 = T_90[23:16];
  assign T_138 = T_133[7:4];
  assign GEN_19 = {{4'd0}, T_138};
  assign T_139 = GEN_19 & 8'hf;
  assign T_140 = T_133[3:0];
  assign GEN_20 = {{4'd0}, T_140};
  assign T_141 = GEN_20 << 4;
  assign T_143 = T_141 & 8'hf0;
  assign T_144 = T_139 | T_143;
  assign T_148 = T_144[7:2];
  assign GEN_21 = {{2'd0}, T_148};
  assign T_149 = GEN_21 & 8'h33;
  assign T_150 = T_144[5:0];
  assign GEN_22 = {{2'd0}, T_150};
  assign T_151 = GEN_22 << 2;
  assign T_153 = T_151 & 8'hcc;
  assign T_154 = T_149 | T_153;
  assign T_158 = T_154[7:1];
  assign GEN_23 = {{1'd0}, T_158};
  assign T_159 = GEN_23 & 8'h55;
  assign T_160 = T_154[6:0];
  assign GEN_24 = {{1'd0}, T_160};
  assign T_161 = GEN_24 << 1;
  assign T_163 = T_161 & 8'haa;
  assign T_164 = T_159 | T_163;
  assign CExtraMask = {T_132,T_164};
  assign T_165 = ~ sigC;
  assign negSigC = doSubMags ? T_165 : sigC;
  assign GEN_25 = {{49'd0}, doSubMags};
  assign T_167 = 50'h0 - GEN_25;
  assign T_168 = T_167[49:0];
  assign T_169 = {doSubMags,negSigC};
  assign T_170 = {T_169,T_168};
  assign T_171 = $signed(T_170);
  assign T_172 = $signed(T_171) >>> CAlignDist;
  assign T_173 = sigC & CExtraMask;
  assign GEN_26 = {{23'd0}, 1'h0};
  assign T_175 = T_173 != GEN_26;
  assign T_176 = T_175 ^ doSubMags;
  assign T_177 = $unsigned(T_172);
  assign T_178 = {T_177,T_176};
  assign alignedNegSigC = T_178[74:0];
  assign T_179 = alignedNegSigC[48:1];
  assign T_181 = fractA[22];
  assign T_183 = fractB[22];
  assign T_185 = fractC[22];
  assign T_186 = alignedNegSigC[0];
  assign T_187 = alignedNegSigC[74:49];
endmodule
module MulAddRecFN_postMul(
  input   clk,
  input   reset,
  input  [2:0] io_fromPreMul_highExpA,
  input   io_fromPreMul_isNaN_isQuietNaNA,
  input  [2:0] io_fromPreMul_highExpB,
  input   io_fromPreMul_isNaN_isQuietNaNB,
  input   io_fromPreMul_signProd,
  input   io_fromPreMul_isZeroProd,
  input   io_fromPreMul_opSignC,
  input  [2:0] io_fromPreMul_highExpC,
  input   io_fromPreMul_isNaN_isQuietNaNC,
  input   io_fromPreMul_isCDominant,
  input   io_fromPreMul_CAlignDist_0,
  input  [6:0] io_fromPreMul_CAlignDist,
  input   io_fromPreMul_bit0AlignedNegSigC,
  input  [25:0] io_fromPreMul_highAlignedNegSigC,
  input  [10:0] io_fromPreMul_sExpSum,
  input  [1:0] io_fromPreMul_roundingMode,
  input  [48:0] io_mulAddResult,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [2:0] GEN_0;
  wire  isZeroA;
  wire [1:0] T_38;
  wire  isSpecialA;
  wire  T_40;
  wire  T_42;
  wire  isInfA;
  wire  isNaNA;
  wire  T_45;
  wire  isSigNaNA;
  wire  isZeroB;
  wire [1:0] T_47;
  wire  isSpecialB;
  wire  T_49;
  wire  T_51;
  wire  isInfB;
  wire  isNaNB;
  wire  T_54;
  wire  isSigNaNB;
  wire  isZeroC;
  wire [1:0] T_56;
  wire  isSpecialC;
  wire  T_58;
  wire  T_60;
  wire  isInfC;
  wire  isNaNC;
  wire  T_63;
  wire  isSigNaNC;
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  doSubMags;
  wire  T_70;
  wire [25:0] GEN_3;
  wire [26:0] T_72;
  wire [25:0] T_73;
  wire [25:0] T_74;
  wire [47:0] T_75;
  wire [73:0] T_76;
  wire [74:0] sigSum;
  wire [49:0] T_78;
  wire [50:0] GEN_4;
  wire [50:0] T_81;
  wire [50:0] T_82;
  wire [49:0] T_84;
  wire  T_85;
  wire  T_87;
  wire  T_89;
  wire  T_91;
  wire  T_93;
  wire  T_95;
  wire  T_97;
  wire  T_99;
  wire  T_101;
  wire  T_103;
  wire  T_105;
  wire  T_107;
  wire  T_109;
  wire  T_111;
  wire  T_113;
  wire  T_115;
  wire  T_117;
  wire  T_119;
  wire  T_121;
  wire  T_123;
  wire  T_125;
  wire  T_127;
  wire  T_129;
  wire  T_131;
  wire  T_133;
  wire  T_135;
  wire  T_137;
  wire  T_139;
  wire  T_141;
  wire  T_143;
  wire  T_145;
  wire  T_147;
  wire  T_149;
  wire  T_151;
  wire  T_153;
  wire  T_155;
  wire  T_157;
  wire  T_159;
  wire  T_161;
  wire  T_163;
  wire  T_165;
  wire  T_167;
  wire  T_169;
  wire  T_171;
  wire  T_173;
  wire  T_175;
  wire  T_177;
  wire  T_179;
  wire  T_181;
  wire [1:0] T_183;
  wire [1:0] T_184;
  wire [2:0] T_185;
  wire [2:0] T_186;
  wire [2:0] T_187;
  wire [2:0] T_188;
  wire [3:0] T_189;
  wire [3:0] T_190;
  wire [3:0] T_191;
  wire [3:0] T_192;
  wire [3:0] T_193;
  wire [3:0] T_194;
  wire [3:0] T_195;
  wire [3:0] T_196;
  wire [4:0] T_197;
  wire [4:0] T_198;
  wire [4:0] T_199;
  wire [4:0] T_200;
  wire [4:0] T_201;
  wire [4:0] T_202;
  wire [4:0] T_203;
  wire [4:0] T_204;
  wire [4:0] T_205;
  wire [4:0] T_206;
  wire [4:0] T_207;
  wire [4:0] T_208;
  wire [4:0] T_209;
  wire [4:0] T_210;
  wire [4:0] T_211;
  wire [4:0] T_212;
  wire [5:0] T_213;
  wire [5:0] T_214;
  wire [5:0] T_215;
  wire [5:0] T_216;
  wire [5:0] T_217;
  wire [5:0] T_218;
  wire [5:0] T_219;
  wire [5:0] T_220;
  wire [5:0] T_221;
  wire [5:0] T_222;
  wire [5:0] T_223;
  wire [5:0] T_224;
  wire [5:0] T_225;
  wire [5:0] T_226;
  wire [5:0] T_227;
  wire [5:0] T_228;
  wire [5:0] T_229;
  wire [5:0] T_230;
  wire [6:0] GEN_6;
  wire [7:0] T_231;
  wire [6:0] estNormPos_dist;
  wire [15:0] T_232;
  wire [15:0] GEN_7;
  wire  T_234;
  wire [17:0] T_235;
  wire [17:0] GEN_8;
  wire  T_237;
  wire [1:0] firstReduceSigSum;
  wire [74:0] complSigSum;
  wire [15:0] T_238;
  wire  T_240;
  wire [17:0] T_241;
  wire  T_243;
  wire [1:0] firstReduceComplSigSum;
  wire  T_244;
  wire [6:0] GEN_11;
  wire [7:0] T_246;
  wire [6:0] T_247;
  wire [4:0] T_248;
  wire [6:0] CDom_estNormDist;
  wire  T_250;
  wire  T_251;
  wire  T_253;
  wire  T_254;
  wire [40:0] T_255;
  wire [1:0] GEN_12;
  wire  T_257;
  wire [41:0] T_258;
  wire [41:0] T_260;
  wire  T_264;
  wire [40:0] T_265;
  wire  T_266;
  wire [41:0] T_267;
  wire [41:0] T_269;
  wire [41:0] T_270;
  wire  T_274;
  wire [40:0] T_275;
  wire  T_277;
  wire [41:0] T_278;
  wire [41:0] T_280;
  wire [41:0] T_281;
  wire  T_283;
  wire [40:0] T_284;
  wire  T_285;
  wire [41:0] T_286;
  wire [41:0] T_288;
  wire [41:0] CDom_firstNormAbsSigSum;
  wire [32:0] T_289;
  wire  T_292;
  wire  T_294;
  wire [33:0] T_295;
  wire [41:0] T_296;
  wire  T_297;
  wire  T_298;
  wire [25:0] T_299;
  wire [15:0] GEN_14;
  wire [16:0] T_301;
  wire [15:0] T_302;
  wire [41:0] T_303;
  wire [41:0] T_304;
  wire [9:0] T_306;
  wire [31:0] GEN_15;
  wire [32:0] T_308;
  wire [31:0] T_309;
  wire [41:0] T_310;
  wire [41:0] T_311;
  wire [41:0] notCDom_pos_firstNormAbsSigSum;
  wire [31:0] T_312;
  wire [32:0] T_314;
  wire [41:0] T_315;
  wire [26:0] T_318;
  wire [42:0] GEN_16;
  wire [42:0] T_319;
  wire [42:0] T_320;
  wire [10:0] T_322;
  wire [42:0] GEN_17;
  wire [42:0] T_323;
  wire [42:0] T_324;
  wire [42:0] notCDom_neg_cFirstNormAbsSigSum;
  wire  notCDom_signSigSum;
  wire  T_326;
  wire  T_327;
  wire  doNegSignSum;
  wire [6:0] estNormDist;
  wire [42:0] T_329;
  wire [41:0] T_330;
  wire [42:0] cFirstNormAbsSigSum;
  wire  T_332;
  wire  T_334;
  wire  T_335;
  wire  doIncrSig;
  wire [3:0] estNormDist_5;
  wire [3:0] normTo2ShiftDist;
  wire [16:0] GEN_18;
  wire [16:0] T_337;
  wire [14:0] T_338;
  wire [7:0] T_339;
  wire [3:0] T_344;
  wire [7:0] GEN_19;
  wire [7:0] T_345;
  wire [3:0] T_346;
  wire [7:0] GEN_20;
  wire [7:0] T_347;
  wire [7:0] T_349;
  wire [7:0] T_350;
  wire [5:0] T_354;
  wire [7:0] GEN_21;
  wire [7:0] T_355;
  wire [5:0] T_356;
  wire [7:0] GEN_22;
  wire [7:0] T_357;
  wire [7:0] T_359;
  wire [7:0] T_360;
  wire [6:0] T_364;
  wire [7:0] GEN_23;
  wire [7:0] T_365;
  wire [6:0] T_366;
  wire [7:0] GEN_24;
  wire [7:0] T_367;
  wire [7:0] T_369;
  wire [7:0] T_370;
  wire [6:0] T_371;
  wire [3:0] T_372;
  wire [1:0] T_373;
  wire  T_374;
  wire  T_375;
  wire [1:0] T_376;
  wire [1:0] T_377;
  wire  T_378;
  wire  T_379;
  wire [1:0] T_380;
  wire [3:0] T_381;
  wire [2:0] T_382;
  wire [1:0] T_383;
  wire  T_384;
  wire  T_385;
  wire [1:0] T_386;
  wire  T_387;
  wire [2:0] T_388;
  wire [6:0] T_389;
  wire [14:0] T_390;
  wire [15:0] absSigSumExtraMask;
  wire [41:0] T_392;
  wire [41:0] T_393;
  wire [15:0] T_394;
  wire [15:0] T_395;
  wire [15:0] T_396;
  wire  T_398;
  wire [15:0] T_400;
  wire  T_402;
  wire  T_403;
  wire [42:0] T_404;
  wire [27:0] sigX3;
  wire [1:0] T_405;
  wire  sigX3Shift1;
  wire [10:0] GEN_28;
  wire [11:0] T_407;
  wire [10:0] sExpX3;
  wire [2:0] T_408;
  wire  isZeroY;
  wire  T_410;
  wire  signY;
  wire [9:0] sExpX3_13;
  wire  T_411;
  wire [26:0] GEN_30;
  wire [27:0] T_413;
  wire [26:0] T_414;
  wire [9:0] T_415;
  wire [1024:0] GEN_31;
  wire [1024:0] T_417;
  wire [24:0] T_418;
  wire [15:0] T_419;
  wire [7:0] T_424;
  wire [15:0] GEN_32;
  wire [15:0] T_425;
  wire [7:0] T_426;
  wire [15:0] GEN_33;
  wire [15:0] T_427;
  wire [15:0] T_429;
  wire [15:0] T_430;
  wire [11:0] T_434;
  wire [15:0] GEN_34;
  wire [15:0] T_435;
  wire [11:0] T_436;
  wire [15:0] GEN_35;
  wire [15:0] T_437;
  wire [15:0] T_439;
  wire [15:0] T_440;
  wire [13:0] T_444;
  wire [15:0] GEN_36;
  wire [15:0] T_445;
  wire [13:0] T_446;
  wire [15:0] GEN_37;
  wire [15:0] T_447;
  wire [15:0] T_449;
  wire [15:0] T_450;
  wire [14:0] T_454;
  wire [15:0] GEN_38;
  wire [15:0] T_455;
  wire [14:0] T_456;
  wire [15:0] GEN_39;
  wire [15:0] T_457;
  wire [15:0] T_459;
  wire [15:0] T_460;
  wire [8:0] T_461;
  wire [7:0] T_462;
  wire [3:0] T_467;
  wire [7:0] GEN_40;
  wire [7:0] T_468;
  wire [3:0] T_469;
  wire [7:0] GEN_41;
  wire [7:0] T_470;
  wire [7:0] T_472;
  wire [7:0] T_473;
  wire [5:0] T_477;
  wire [7:0] GEN_42;
  wire [7:0] T_478;
  wire [5:0] T_479;
  wire [7:0] GEN_43;
  wire [7:0] T_480;
  wire [7:0] T_482;
  wire [7:0] T_483;
  wire [6:0] T_487;
  wire [7:0] GEN_44;
  wire [7:0] T_488;
  wire [6:0] T_489;
  wire [7:0] GEN_45;
  wire [7:0] T_490;
  wire [7:0] T_492;
  wire [7:0] T_493;
  wire  T_494;
  wire [8:0] T_495;
  wire [24:0] T_496;
  wire  T_497;
  wire [24:0] GEN_46;
  wire [24:0] T_498;
  wire [26:0] T_500;
  wire [26:0] roundMask;
  wire [25:0] T_501;
  wire [25:0] T_502;
  wire [26:0] GEN_47;
  wire [26:0] roundPosMask;
  wire [27:0] GEN_48;
  wire [27:0] T_503;
  wire [27:0] GEN_49;
  wire  roundPosBit;
  wire [27:0] GEN_50;
  wire [27:0] T_506;
  wire  anyRoundExtra;
  wire [27:0] T_508;
  wire [27:0] T_510;
  wire  allRoundExtra;
  wire  anyRound;
  wire  allRound;
  wire  roundDirectUp;
  wire  T_513;
  wire  T_514;
  wire  T_515;
  wire  T_516;
  wire  T_519;
  wire  T_520;
  wire  T_521;
  wire  T_522;
  wire  T_523;
  wire  T_524;
  wire  T_525;
  wire  T_526;
  wire  T_527;
  wire  roundUp;
  wire  T_531;
  wire  T_532;
  wire  T_533;
  wire  T_534;
  wire  T_536;
  wire  T_537;
  wire  roundEven;
  wire  T_539;
  wire  roundInexact;
  wire [27:0] GEN_54;
  wire [27:0] T_540;
  wire [25:0] T_541;
  wire [26:0] T_543;
  wire [25:0] T_544;
  wire  T_546;
  wire  T_548;
  wire  T_549;
  wire [26:0] T_550;
  wire [27:0] GEN_56;
  wire [27:0] T_551;
  wire [25:0] T_552;
  wire [25:0] T_554;
  wire [25:0] T_556;
  wire [25:0] T_557;
  wire [25:0] T_560;
  wire [25:0] T_562;
  wire [25:0] sigY3;
  wire  T_563;
  wire [10:0] GEN_57;
  wire [11:0] T_565;
  wire [10:0] T_566;
  wire [10:0] T_568;
  wire  T_569;
  wire [10:0] T_571;
  wire [10:0] T_572;
  wire [1:0] T_573;
  wire  T_575;
  wire [11:0] T_577;
  wire [10:0] T_578;
  wire [10:0] T_580;
  wire [10:0] sExpY;
  wire [8:0] expY;
  wire [22:0] T_581;
  wire [22:0] T_582;
  wire [22:0] fractY;
  wire [2:0] T_583;
  wire [2:0] GEN_60;
  wire  overflowY;
  wire  T_586;
  wire  T_587;
  wire [8:0] GEN_61;
  wire  T_590;
  wire  T_591;
  wire  totalUnderflowY;
  wire [7:0] T_595;
  wire [9:0] GEN_62;
  wire  T_596;
  wire  T_597;
  wire  underflowY;
  wire  T_598;
  wire  T_600;
  wire  T_601;
  wire  roundMagUp;
  wire  overflowY_roundMagUp;
  wire  mulSpecial;
  wire  addSpecial;
  wire  notSpecial_addZeros;
  wire  T_603;
  wire  T_605;
  wire  commonCase;
  wire  T_606;
  wire  T_607;
  wire  T_608;
  wire  T_610;
  wire  T_612;
  wire  T_613;
  wire  T_614;
  wire  T_615;
  wire  T_616;
  wire  T_617;
  wire  notSigNaN_invalid;
  wire  T_618;
  wire  T_619;
  wire  invalid;
  wire  overflow;
  wire  underflow;
  wire  T_620;
  wire  inexact;
  wire  T_621;
  wire  notSpecial_isZeroOut;
  wire  T_622;
  wire  pegMinFiniteMagOut;
  wire  T_624;
  wire  pegMaxFiniteMagOut;
  wire  T_626;
  wire  T_627;
  wire  notNaN_isInfOut;
  wire  T_628;
  wire  T_629;
  wire  isNaNOut;
  wire  T_632;
  wire  T_634;
  wire  T_635;
  wire  T_636;
  wire  T_637;
  wire  T_639;
  wire  T_640;
  wire  T_641;
  wire  T_642;
  wire  T_645;
  wire  T_646;
  wire  T_647;
  wire  uncommonCaseSignOut;
  wire  T_649;
  wire  T_650;
  wire  T_651;
  wire  signOut;
  wire [8:0] T_654;
  wire [8:0] T_655;
  wire [8:0] T_656;
  wire [8:0] T_660;
  wire [8:0] T_661;
  wire [8:0] T_662;
  wire [8:0] T_665;
  wire [8:0] T_666;
  wire [8:0] T_667;
  wire [8:0] T_670;
  wire [8:0] T_671;
  wire [8:0] T_672;
  wire [8:0] T_675;
  wire [8:0] T_676;
  wire [8:0] T_679;
  wire [8:0] T_680;
  wire [8:0] T_683;
  wire [8:0] T_684;
  wire [8:0] T_687;
  wire [8:0] expOut;
  wire  T_688;
  wire  T_689;
  wire [22:0] T_693;
  wire [22:0] T_694;
  wire [22:0] GEN_63;
  wire [23:0] T_696;
  wire [22:0] T_697;
  wire [22:0] fractOut;
  wire [9:0] T_698;
  wire [32:0] T_699;
  wire [1:0] T_701;
  wire [1:0] T_702;
  wire [2:0] T_703;
  wire [4:0] T_704;
  assign io_out = T_699;
  assign io_exceptionFlags = T_704;
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZeroA = io_fromPreMul_highExpA == GEN_0;
  assign T_38 = io_fromPreMul_highExpA[2:1];
  assign isSpecialA = T_38 == 2'h3;
  assign T_40 = io_fromPreMul_highExpA[0];
  assign T_42 = T_40 == 1'h0;
  assign isInfA = isSpecialA & T_42;
  assign isNaNA = isSpecialA & T_40;
  assign T_45 = io_fromPreMul_isNaN_isQuietNaNA == 1'h0;
  assign isSigNaNA = isNaNA & T_45;
  assign isZeroB = io_fromPreMul_highExpB == GEN_0;
  assign T_47 = io_fromPreMul_highExpB[2:1];
  assign isSpecialB = T_47 == 2'h3;
  assign T_49 = io_fromPreMul_highExpB[0];
  assign T_51 = T_49 == 1'h0;
  assign isInfB = isSpecialB & T_51;
  assign isNaNB = isSpecialB & T_49;
  assign T_54 = io_fromPreMul_isNaN_isQuietNaNB == 1'h0;
  assign isSigNaNB = isNaNB & T_54;
  assign isZeroC = io_fromPreMul_highExpC == GEN_0;
  assign T_56 = io_fromPreMul_highExpC[2:1];
  assign isSpecialC = T_56 == 2'h3;
  assign T_58 = io_fromPreMul_highExpC[0];
  assign T_60 = T_58 == 1'h0;
  assign isInfC = isSpecialC & T_60;
  assign isNaNC = isSpecialC & T_58;
  assign T_63 = io_fromPreMul_isNaN_isQuietNaNC == 1'h0;
  assign isSigNaNC = isNaNC & T_63;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T_70 = io_mulAddResult[48];
  assign GEN_3 = {{25'd0}, 1'h1};
  assign T_72 = io_fromPreMul_highAlignedNegSigC + GEN_3;
  assign T_73 = T_72[25:0];
  assign T_74 = T_70 ? T_73 : io_fromPreMul_highAlignedNegSigC;
  assign T_75 = io_mulAddResult[47:0];
  assign T_76 = {T_74,T_75};
  assign sigSum = {T_76,io_fromPreMul_bit0AlignedNegSigC};
  assign T_78 = sigSum[50:1];
  assign GEN_4 = {{1'd0}, T_78};
  assign T_81 = GEN_4 << 1;
  assign T_82 = GEN_4 ^ T_81;
  assign T_84 = T_82[49:0];
  assign T_85 = T_84[49];
  assign T_87 = T_84[48];
  assign T_89 = T_84[47];
  assign T_91 = T_84[46];
  assign T_93 = T_84[45];
  assign T_95 = T_84[44];
  assign T_97 = T_84[43];
  assign T_99 = T_84[42];
  assign T_101 = T_84[41];
  assign T_103 = T_84[40];
  assign T_105 = T_84[39];
  assign T_107 = T_84[38];
  assign T_109 = T_84[37];
  assign T_111 = T_84[36];
  assign T_113 = T_84[35];
  assign T_115 = T_84[34];
  assign T_117 = T_84[33];
  assign T_119 = T_84[32];
  assign T_121 = T_84[31];
  assign T_123 = T_84[30];
  assign T_125 = T_84[29];
  assign T_127 = T_84[28];
  assign T_129 = T_84[27];
  assign T_131 = T_84[26];
  assign T_133 = T_84[25];
  assign T_135 = T_84[24];
  assign T_137 = T_84[23];
  assign T_139 = T_84[22];
  assign T_141 = T_84[21];
  assign T_143 = T_84[20];
  assign T_145 = T_84[19];
  assign T_147 = T_84[18];
  assign T_149 = T_84[17];
  assign T_151 = T_84[16];
  assign T_153 = T_84[15];
  assign T_155 = T_84[14];
  assign T_157 = T_84[13];
  assign T_159 = T_84[12];
  assign T_161 = T_84[11];
  assign T_163 = T_84[10];
  assign T_165 = T_84[9];
  assign T_167 = T_84[8];
  assign T_169 = T_84[7];
  assign T_171 = T_84[6];
  assign T_173 = T_84[5];
  assign T_175 = T_84[4];
  assign T_177 = T_84[3];
  assign T_179 = T_84[2];
  assign T_181 = T_84[1];
  assign T_183 = T_179 ? 2'h2 : {{1'd0}, T_181};
  assign T_184 = T_177 ? 2'h3 : T_183;
  assign T_185 = T_175 ? 3'h4 : {{1'd0}, T_184};
  assign T_186 = T_173 ? 3'h5 : T_185;
  assign T_187 = T_171 ? 3'h6 : T_186;
  assign T_188 = T_169 ? 3'h7 : T_187;
  assign T_189 = T_167 ? 4'h8 : {{1'd0}, T_188};
  assign T_190 = T_165 ? 4'h9 : T_189;
  assign T_191 = T_163 ? 4'ha : T_190;
  assign T_192 = T_161 ? 4'hb : T_191;
  assign T_193 = T_159 ? 4'hc : T_192;
  assign T_194 = T_157 ? 4'hd : T_193;
  assign T_195 = T_155 ? 4'he : T_194;
  assign T_196 = T_153 ? 4'hf : T_195;
  assign T_197 = T_151 ? 5'h10 : {{1'd0}, T_196};
  assign T_198 = T_149 ? 5'h11 : T_197;
  assign T_199 = T_147 ? 5'h12 : T_198;
  assign T_200 = T_145 ? 5'h13 : T_199;
  assign T_201 = T_143 ? 5'h14 : T_200;
  assign T_202 = T_141 ? 5'h15 : T_201;
  assign T_203 = T_139 ? 5'h16 : T_202;
  assign T_204 = T_137 ? 5'h17 : T_203;
  assign T_205 = T_135 ? 5'h18 : T_204;
  assign T_206 = T_133 ? 5'h19 : T_205;
  assign T_207 = T_131 ? 5'h1a : T_206;
  assign T_208 = T_129 ? 5'h1b : T_207;
  assign T_209 = T_127 ? 5'h1c : T_208;
  assign T_210 = T_125 ? 5'h1d : T_209;
  assign T_211 = T_123 ? 5'h1e : T_210;
  assign T_212 = T_121 ? 5'h1f : T_211;
  assign T_213 = T_119 ? 6'h20 : {{1'd0}, T_212};
  assign T_214 = T_117 ? 6'h21 : T_213;
  assign T_215 = T_115 ? 6'h22 : T_214;
  assign T_216 = T_113 ? 6'h23 : T_215;
  assign T_217 = T_111 ? 6'h24 : T_216;
  assign T_218 = T_109 ? 6'h25 : T_217;
  assign T_219 = T_107 ? 6'h26 : T_218;
  assign T_220 = T_105 ? 6'h27 : T_219;
  assign T_221 = T_103 ? 6'h28 : T_220;
  assign T_222 = T_101 ? 6'h29 : T_221;
  assign T_223 = T_99 ? 6'h2a : T_222;
  assign T_224 = T_97 ? 6'h2b : T_223;
  assign T_225 = T_95 ? 6'h2c : T_224;
  assign T_226 = T_93 ? 6'h2d : T_225;
  assign T_227 = T_91 ? 6'h2e : T_226;
  assign T_228 = T_89 ? 6'h2f : T_227;
  assign T_229 = T_87 ? 6'h30 : T_228;
  assign T_230 = T_85 ? 6'h31 : T_229;
  assign GEN_6 = {{1'd0}, T_230};
  assign T_231 = 7'h49 - GEN_6;
  assign estNormPos_dist = T_231[6:0];
  assign T_232 = sigSum[33:18];
  assign GEN_7 = {{15'd0}, 1'h0};
  assign T_234 = T_232 != GEN_7;
  assign T_235 = sigSum[17:0];
  assign GEN_8 = {{17'd0}, 1'h0};
  assign T_237 = T_235 != GEN_8;
  assign firstReduceSigSum = {T_234,T_237};
  assign complSigSum = ~ sigSum;
  assign T_238 = complSigSum[33:18];
  assign T_240 = T_238 != GEN_7;
  assign T_241 = complSigSum[17:0];
  assign T_243 = T_241 != GEN_8;
  assign firstReduceComplSigSum = {T_240,T_243};
  assign T_244 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign GEN_11 = {{6'd0}, 1'h1};
  assign T_246 = io_fromPreMul_CAlignDist - GEN_11;
  assign T_247 = T_246[6:0];
  assign T_248 = T_247[4:0];
  assign CDom_estNormDist = T_244 ? io_fromPreMul_CAlignDist : {{2'd0}, T_248};
  assign T_250 = doSubMags == 1'h0;
  assign T_251 = CDom_estNormDist[4];
  assign T_253 = T_251 == 1'h0;
  assign T_254 = T_250 & T_253;
  assign T_255 = sigSum[74:34];
  assign GEN_12 = {{1'd0}, 1'h0};
  assign T_257 = firstReduceSigSum != GEN_12;
  assign T_258 = {T_255,T_257};
  assign T_260 = T_254 ? T_258 : {{41'd0}, 1'h0};
  assign T_264 = T_250 & T_251;
  assign T_265 = sigSum[58:18];
  assign T_266 = firstReduceSigSum[0];
  assign T_267 = {T_265,T_266};
  assign T_269 = T_264 ? T_267 : {{41'd0}, 1'h0};
  assign T_270 = T_260 | T_269;
  assign T_274 = doSubMags & T_253;
  assign T_275 = complSigSum[74:34];
  assign T_277 = firstReduceComplSigSum != GEN_12;
  assign T_278 = {T_275,T_277};
  assign T_280 = T_274 ? T_278 : {{41'd0}, 1'h0};
  assign T_281 = T_270 | T_280;
  assign T_283 = doSubMags & T_251;
  assign T_284 = complSigSum[58:18];
  assign T_285 = firstReduceComplSigSum[0];
  assign T_286 = {T_284,T_285};
  assign T_288 = T_283 ? T_286 : {{41'd0}, 1'h0};
  assign CDom_firstNormAbsSigSum = T_281 | T_288;
  assign T_289 = sigSum[50:18];
  assign T_292 = T_285 == 1'h0;
  assign T_294 = doSubMags ? T_292 : T_266;
  assign T_295 = {T_289,T_294};
  assign T_296 = sigSum[42:1];
  assign T_297 = estNormPos_dist[5];
  assign T_298 = estNormPos_dist[4];
  assign T_299 = sigSum[26:1];
  assign GEN_14 = {{15'd0}, doSubMags};
  assign T_301 = 16'h0 - GEN_14;
  assign T_302 = T_301[15:0];
  assign T_303 = {T_299,T_302};
  assign T_304 = T_298 ? T_303 : T_296;
  assign T_306 = sigSum[10:1];
  assign GEN_15 = {{31'd0}, doSubMags};
  assign T_308 = 32'h0 - GEN_15;
  assign T_309 = T_308[31:0];
  assign T_310 = {T_306,T_309};
  assign T_311 = T_298 ? {{8'd0}, T_295} : T_310;
  assign notCDom_pos_firstNormAbsSigSum = T_297 ? T_304 : T_311;
  assign T_312 = complSigSum[49:18];
  assign T_314 = {T_312,T_285};
  assign T_315 = complSigSum[42:1];
  assign T_318 = complSigSum[27:1];
  assign GEN_16 = {{16'd0}, T_318};
  assign T_319 = GEN_16 << 16;
  assign T_320 = T_298 ? T_319 : {{1'd0}, T_315};
  assign T_322 = complSigSum[11:1];
  assign GEN_17 = {{32'd0}, T_322};
  assign T_323 = GEN_17 << 32;
  assign T_324 = T_298 ? {{10'd0}, T_314} : T_323;
  assign notCDom_neg_cFirstNormAbsSigSum = T_297 ? T_320 : T_324;
  assign notCDom_signSigSum = sigSum[51];
  assign T_326 = isZeroC == 1'h0;
  assign T_327 = doSubMags & T_326;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T_327 : notCDom_signSigSum;
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : estNormPos_dist;
  assign T_329 = io_fromPreMul_isCDominant ? {{1'd0}, CDom_firstNormAbsSigSum} : notCDom_neg_cFirstNormAbsSigSum;
  assign T_330 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T_329 : {{1'd0}, T_330};
  assign T_332 = io_fromPreMul_isCDominant == 1'h0;
  assign T_334 = notCDom_signSigSum == 1'h0;
  assign T_335 = T_332 & T_334;
  assign doIncrSig = T_335 & doSubMags;
  assign estNormDist_5 = estNormDist[3:0];
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign GEN_18 = $signed(17'h10000);
  assign T_337 = $signed(GEN_18) >>> normTo2ShiftDist;
  assign T_338 = T_337[15:1];
  assign T_339 = T_338[7:0];
  assign T_344 = T_339[7:4];
  assign GEN_19 = {{4'd0}, T_344};
  assign T_345 = GEN_19 & 8'hf;
  assign T_346 = T_339[3:0];
  assign GEN_20 = {{4'd0}, T_346};
  assign T_347 = GEN_20 << 4;
  assign T_349 = T_347 & 8'hf0;
  assign T_350 = T_345 | T_349;
  assign T_354 = T_350[7:2];
  assign GEN_21 = {{2'd0}, T_354};
  assign T_355 = GEN_21 & 8'h33;
  assign T_356 = T_350[5:0];
  assign GEN_22 = {{2'd0}, T_356};
  assign T_357 = GEN_22 << 2;
  assign T_359 = T_357 & 8'hcc;
  assign T_360 = T_355 | T_359;
  assign T_364 = T_360[7:1];
  assign GEN_23 = {{1'd0}, T_364};
  assign T_365 = GEN_23 & 8'h55;
  assign T_366 = T_360[6:0];
  assign GEN_24 = {{1'd0}, T_366};
  assign T_367 = GEN_24 << 1;
  assign T_369 = T_367 & 8'haa;
  assign T_370 = T_365 | T_369;
  assign T_371 = T_338[14:8];
  assign T_372 = T_371[3:0];
  assign T_373 = T_372[1:0];
  assign T_374 = T_373[0];
  assign T_375 = T_373[1];
  assign T_376 = {T_374,T_375};
  assign T_377 = T_372[3:2];
  assign T_378 = T_377[0];
  assign T_379 = T_377[1];
  assign T_380 = {T_378,T_379};
  assign T_381 = {T_376,T_380};
  assign T_382 = T_371[6:4];
  assign T_383 = T_382[1:0];
  assign T_384 = T_383[0];
  assign T_385 = T_383[1];
  assign T_386 = {T_384,T_385};
  assign T_387 = T_382[2];
  assign T_388 = {T_386,T_387};
  assign T_389 = {T_381,T_388};
  assign T_390 = {T_370,T_389};
  assign absSigSumExtraMask = {T_390,1'h1};
  assign T_392 = cFirstNormAbsSigSum[42:1];
  assign T_393 = T_392 >> normTo2ShiftDist;
  assign T_394 = cFirstNormAbsSigSum[15:0];
  assign T_395 = ~ T_394;
  assign T_396 = T_395 & absSigSumExtraMask;
  assign T_398 = T_396 == GEN_7;
  assign T_400 = T_394 & absSigSumExtraMask;
  assign T_402 = T_400 != GEN_7;
  assign T_403 = doIncrSig ? T_398 : T_402;
  assign T_404 = {T_393,T_403};
  assign sigX3 = T_404[27:0];
  assign T_405 = sigX3[27:26];
  assign sigX3Shift1 = T_405 == GEN_12;
  assign GEN_28 = {{4'd0}, estNormDist};
  assign T_407 = io_fromPreMul_sExpSum - GEN_28;
  assign sExpX3 = T_407[10:0];
  assign T_408 = sigX3[27:25];
  assign isZeroY = T_408 == GEN_0;
  assign T_410 = io_fromPreMul_signProd ^ doNegSignSum;
  assign signY = isZeroY ? roundingMode_min : T_410;
  assign sExpX3_13 = sExpX3[9:0];
  assign T_411 = sExpX3[10];
  assign GEN_30 = {{26'd0}, T_411};
  assign T_413 = 27'h0 - GEN_30;
  assign T_414 = T_413[26:0];
  assign T_415 = ~ sExpX3_13;
  assign GEN_31 = $signed(1025'h10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign T_417 = $signed(GEN_31) >>> T_415;
  assign T_418 = T_417[131:107];
  assign T_419 = T_418[15:0];
  assign T_424 = T_419[15:8];
  assign GEN_32 = {{8'd0}, T_424};
  assign T_425 = GEN_32 & 16'hff;
  assign T_426 = T_419[7:0];
  assign GEN_33 = {{8'd0}, T_426};
  assign T_427 = GEN_33 << 8;
  assign T_429 = T_427 & 16'hff00;
  assign T_430 = T_425 | T_429;
  assign T_434 = T_430[15:4];
  assign GEN_34 = {{4'd0}, T_434};
  assign T_435 = GEN_34 & 16'hf0f;
  assign T_436 = T_430[11:0];
  assign GEN_35 = {{4'd0}, T_436};
  assign T_437 = GEN_35 << 4;
  assign T_439 = T_437 & 16'hf0f0;
  assign T_440 = T_435 | T_439;
  assign T_444 = T_440[15:2];
  assign GEN_36 = {{2'd0}, T_444};
  assign T_445 = GEN_36 & 16'h3333;
  assign T_446 = T_440[13:0];
  assign GEN_37 = {{2'd0}, T_446};
  assign T_447 = GEN_37 << 2;
  assign T_449 = T_447 & 16'hcccc;
  assign T_450 = T_445 | T_449;
  assign T_454 = T_450[15:1];
  assign GEN_38 = {{1'd0}, T_454};
  assign T_455 = GEN_38 & 16'h5555;
  assign T_456 = T_450[14:0];
  assign GEN_39 = {{1'd0}, T_456};
  assign T_457 = GEN_39 << 1;
  assign T_459 = T_457 & 16'haaaa;
  assign T_460 = T_455 | T_459;
  assign T_461 = T_418[24:16];
  assign T_462 = T_461[7:0];
  assign T_467 = T_462[7:4];
  assign GEN_40 = {{4'd0}, T_467};
  assign T_468 = GEN_40 & 8'hf;
  assign T_469 = T_462[3:0];
  assign GEN_41 = {{4'd0}, T_469};
  assign T_470 = GEN_41 << 4;
  assign T_472 = T_470 & 8'hf0;
  assign T_473 = T_468 | T_472;
  assign T_477 = T_473[7:2];
  assign GEN_42 = {{2'd0}, T_477};
  assign T_478 = GEN_42 & 8'h33;
  assign T_479 = T_473[5:0];
  assign GEN_43 = {{2'd0}, T_479};
  assign T_480 = GEN_43 << 2;
  assign T_482 = T_480 & 8'hcc;
  assign T_483 = T_478 | T_482;
  assign T_487 = T_483[7:1];
  assign GEN_44 = {{1'd0}, T_487};
  assign T_488 = GEN_44 & 8'h55;
  assign T_489 = T_483[6:0];
  assign GEN_45 = {{1'd0}, T_489};
  assign T_490 = GEN_45 << 1;
  assign T_492 = T_490 & 8'haa;
  assign T_493 = T_488 | T_492;
  assign T_494 = T_461[8];
  assign T_495 = {T_493,T_494};
  assign T_496 = {T_460,T_495};
  assign T_497 = sigX3[26];
  assign GEN_46 = {{24'd0}, T_497};
  assign T_498 = T_496 | GEN_46;
  assign T_500 = {T_498,2'h3};
  assign roundMask = T_414 | T_500;
  assign T_501 = roundMask[26:1];
  assign T_502 = ~ T_501;
  assign GEN_47 = {{1'd0}, T_502};
  assign roundPosMask = GEN_47 & roundMask;
  assign GEN_48 = {{1'd0}, roundPosMask};
  assign T_503 = sigX3 & GEN_48;
  assign GEN_49 = {{27'd0}, 1'h0};
  assign roundPosBit = T_503 != GEN_49;
  assign GEN_50 = {{2'd0}, T_501};
  assign T_506 = sigX3 & GEN_50;
  assign anyRoundExtra = T_506 != GEN_49;
  assign T_508 = ~ sigX3;
  assign T_510 = T_508 & GEN_50;
  assign allRoundExtra = T_510 == GEN_49;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign allRound = roundPosBit & allRoundExtra;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign T_513 = doIncrSig == 1'h0;
  assign T_514 = T_513 & roundingMode_nearest_even;
  assign T_515 = T_514 & roundPosBit;
  assign T_516 = T_515 & anyRoundExtra;
  assign T_519 = T_513 & roundDirectUp;
  assign T_520 = T_519 & anyRound;
  assign T_521 = T_516 | T_520;
  assign T_522 = doIncrSig & allRound;
  assign T_523 = T_521 | T_522;
  assign T_524 = doIncrSig & roundingMode_nearest_even;
  assign T_525 = T_524 & roundPosBit;
  assign T_526 = T_523 | T_525;
  assign T_527 = doIncrSig & roundDirectUp;
  assign roundUp = T_526 | T_527;
  assign T_531 = roundPosBit == 1'h0;
  assign T_532 = roundingMode_nearest_even & T_531;
  assign T_533 = T_532 & allRoundExtra;
  assign T_534 = roundingMode_nearest_even & roundPosBit;
  assign T_536 = anyRoundExtra == 1'h0;
  assign T_537 = T_534 & T_536;
  assign roundEven = doIncrSig ? T_533 : T_537;
  assign T_539 = allRound == 1'h0;
  assign roundInexact = doIncrSig ? T_539 : anyRound;
  assign GEN_54 = {{1'd0}, roundMask};
  assign T_540 = sigX3 | GEN_54;
  assign T_541 = T_540[27:2];
  assign T_543 = T_541 + GEN_3;
  assign T_544 = T_543[25:0];
  assign T_546 = roundUp == 1'h0;
  assign T_548 = roundEven == 1'h0;
  assign T_549 = T_546 & T_548;
  assign T_550 = ~ roundMask;
  assign GEN_56 = {{1'd0}, T_550};
  assign T_551 = sigX3 & GEN_56;
  assign T_552 = T_551[27:2];
  assign T_554 = T_549 ? T_552 : {{25'd0}, 1'h0};
  assign T_556 = roundUp ? T_544 : {{25'd0}, 1'h0};
  assign T_557 = T_554 | T_556;
  assign T_560 = T_544 & T_502;
  assign T_562 = roundEven ? T_560 : {{25'd0}, 1'h0};
  assign sigY3 = T_557 | T_562;
  assign T_563 = sigY3[25];
  assign GEN_57 = {{10'd0}, 1'h1};
  assign T_565 = sExpX3 + GEN_57;
  assign T_566 = T_565[10:0];
  assign T_568 = T_563 ? T_566 : {{10'd0}, 1'h0};
  assign T_569 = sigY3[24];
  assign T_571 = T_569 ? sExpX3 : {{10'd0}, 1'h0};
  assign T_572 = T_568 | T_571;
  assign T_573 = sigY3[25:24];
  assign T_575 = T_573 == GEN_12;
  assign T_577 = sExpX3 - GEN_57;
  assign T_578 = T_577[10:0];
  assign T_580 = T_575 ? T_578 : {{10'd0}, 1'h0};
  assign sExpY = T_572 | T_580;
  assign expY = sExpY[8:0];
  assign T_581 = sigY3[22:0];
  assign T_582 = sigY3[23:1];
  assign fractY = sigX3Shift1 ? T_581 : T_582;
  assign T_583 = sExpY[9:7];
  assign GEN_60 = {{1'd0}, 2'h3};
  assign overflowY = T_583 == GEN_60;
  assign T_586 = isZeroY == 1'h0;
  assign T_587 = sExpY[9];
  assign GEN_61 = {{2'd0}, 7'h6b};
  assign T_590 = expY < GEN_61;
  assign T_591 = T_587 | T_590;
  assign totalUnderflowY = T_586 & T_591;
  assign T_595 = sigX3Shift1 ? 8'h82 : 8'h81;
  assign GEN_62 = {{2'd0}, T_595};
  assign T_596 = sExpX3_13 <= GEN_62;
  assign T_597 = T_411 | T_596;
  assign underflowY = roundInexact & T_597;
  assign T_598 = roundingMode_min & signY;
  assign T_600 = signY == 1'h0;
  assign T_601 = roundingMode_max & T_600;
  assign roundMagUp = T_598 | T_601;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign mulSpecial = isSpecialA | isSpecialB;
  assign addSpecial = mulSpecial | isSpecialC;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign T_603 = addSpecial == 1'h0;
  assign T_605 = notSpecial_addZeros == 1'h0;
  assign commonCase = T_603 & T_605;
  assign T_606 = isInfA & isZeroB;
  assign T_607 = isZeroA & isInfB;
  assign T_608 = T_606 | T_607;
  assign T_610 = isNaNA == 1'h0;
  assign T_612 = isNaNB == 1'h0;
  assign T_613 = T_610 & T_612;
  assign T_614 = isInfA | isInfB;
  assign T_615 = T_613 & T_614;
  assign T_616 = T_615 & isInfC;
  assign T_617 = T_616 & doSubMags;
  assign notSigNaN_invalid = T_608 | T_617;
  assign T_618 = isSigNaNA | isSigNaNB;
  assign T_619 = T_618 | isSigNaNC;
  assign invalid = T_619 | notSigNaN_invalid;
  assign overflow = commonCase & overflowY;
  assign underflow = commonCase & underflowY;
  assign T_620 = commonCase & roundInexact;
  assign inexact = overflow | T_620;
  assign T_621 = notSpecial_addZeros | isZeroY;
  assign notSpecial_isZeroOut = T_621 | totalUnderflowY;
  assign T_622 = commonCase & totalUnderflowY;
  assign pegMinFiniteMagOut = T_622 & roundMagUp;
  assign T_624 = overflowY_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = overflow & T_624;
  assign T_626 = T_614 | isInfC;
  assign T_627 = overflow & overflowY_roundMagUp;
  assign notNaN_isInfOut = T_626 | T_627;
  assign T_628 = isNaNA | isNaNB;
  assign T_629 = T_628 | isNaNC;
  assign isNaNOut = T_629 | notSigNaN_invalid;
  assign T_632 = T_250 & io_fromPreMul_opSignC;
  assign T_634 = isSpecialC == 1'h0;
  assign T_635 = mulSpecial & T_634;
  assign T_636 = T_635 & io_fromPreMul_signProd;
  assign T_637 = T_632 | T_636;
  assign T_639 = mulSpecial == 1'h0;
  assign T_640 = T_639 & isSpecialC;
  assign T_641 = T_640 & io_fromPreMul_opSignC;
  assign T_642 = T_637 | T_641;
  assign T_645 = T_639 & notSpecial_addZeros;
  assign T_646 = T_645 & doSubMags;
  assign T_647 = T_646 & roundingMode_min;
  assign uncommonCaseSignOut = T_642 | T_647;
  assign T_649 = isNaNOut == 1'h0;
  assign T_650 = T_649 & uncommonCaseSignOut;
  assign T_651 = commonCase & signY;
  assign signOut = T_650 | T_651;
  assign T_654 = notSpecial_isZeroOut ? 9'h1c0 : 9'h0;
  assign T_655 = ~ T_654;
  assign T_656 = expY & T_655;
  assign T_660 = pegMinFiniteMagOut ? 9'h194 : 9'h0;
  assign T_661 = ~ T_660;
  assign T_662 = T_656 & T_661;
  assign T_665 = pegMaxFiniteMagOut ? 9'h80 : 9'h0;
  assign T_666 = ~ T_665;
  assign T_667 = T_662 & T_666;
  assign T_670 = notNaN_isInfOut ? {{2'd0}, 7'h40} : 9'h0;
  assign T_671 = ~ T_670;
  assign T_672 = T_667 & T_671;
  assign T_675 = pegMinFiniteMagOut ? {{2'd0}, 7'h6b} : 9'h0;
  assign T_676 = T_672 | T_675;
  assign T_679 = pegMaxFiniteMagOut ? 9'h17f : 9'h0;
  assign T_680 = T_676 | T_679;
  assign T_683 = notNaN_isInfOut ? 9'h180 : 9'h0;
  assign T_684 = T_680 | T_683;
  assign T_687 = isNaNOut ? 9'h1c0 : 9'h0;
  assign expOut = T_684 | T_687;
  assign T_688 = totalUnderflowY & roundMagUp;
  assign T_689 = T_688 | isNaNOut;
  assign T_693 = isNaNOut ? 23'h400000 : {{22'd0}, 1'h0};
  assign T_694 = T_689 ? T_693 : fractY;
  assign GEN_63 = {{22'd0}, pegMaxFiniteMagOut};
  assign T_696 = 23'h0 - GEN_63;
  assign T_697 = T_696[22:0];
  assign fractOut = T_694 | T_697;
  assign T_698 = {signOut,expOut};
  assign T_699 = {T_698,fractOut};
  assign T_701 = {underflow,inexact};
  assign T_702 = {invalid,1'h0};
  assign T_703 = {T_702,overflow};
  assign T_704 = {T_703,T_701};
endmodule
module MulAddRecFN(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [32:0] io_a,
  input  [32:0] io_b,
  input  [32:0] io_c,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  mulAddRecFN_preMul_clk;
  wire  mulAddRecFN_preMul_reset;
  wire [1:0] mulAddRecFN_preMul_io_op;
  wire [32:0] mulAddRecFN_preMul_io_a;
  wire [32:0] mulAddRecFN_preMul_io_b;
  wire [32:0] mulAddRecFN_preMul_io_c;
  wire [1:0] mulAddRecFN_preMul_io_roundingMode;
  wire [23:0] mulAddRecFN_preMul_io_mulAddA;
  wire [23:0] mulAddRecFN_preMul_io_mulAddB;
  wire [47:0] mulAddRecFN_preMul_io_mulAddC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_preMul_io_toPostMul_signProd;
  wire  mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire  mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire  mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire [6:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire  mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire [25:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire [10:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire [1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire  mulAddRecFN_postMul_clk;
  wire  mulAddRecFN_postMul_reset;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpA;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpB;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_postMul_io_fromPreMul_signProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_isZeroProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_opSignC;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isCDominant;
  wire  mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0;
  wire [6:0] mulAddRecFN_postMul_io_fromPreMul_CAlignDist;
  wire  mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC;
  wire [25:0] mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC;
  wire [10:0] mulAddRecFN_postMul_io_fromPreMul_sExpSum;
  wire [1:0] mulAddRecFN_postMul_io_fromPreMul_roundingMode;
  wire [48:0] mulAddRecFN_postMul_io_mulAddResult;
  wire [32:0] mulAddRecFN_postMul_io_out;
  wire [4:0] mulAddRecFN_postMul_io_exceptionFlags;
  wire [47:0] T_7;
  wire [48:0] T_9;
  wire [48:0] GEN_0;
  wire [49:0] T_10;
  wire [48:0] T_11;
  MulAddRecFN_preMul mulAddRecFN_preMul (
    .clk(mulAddRecFN_preMul_clk),
    .reset(mulAddRecFN_preMul_reset),
    .io_op(mulAddRecFN_preMul_io_op),
    .io_a(mulAddRecFN_preMul_io_a),
    .io_b(mulAddRecFN_preMul_io_b),
    .io_c(mulAddRecFN_preMul_io_c),
    .io_roundingMode(mulAddRecFN_preMul_io_roundingMode),
    .io_mulAddA(mulAddRecFN_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFN_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFN_preMul_io_mulAddC),
    .io_toPostMul_highExpA(mulAddRecFN_preMul_io_toPostMul_highExpA),
    .io_toPostMul_isNaN_isQuietNaNA(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA),
    .io_toPostMul_highExpB(mulAddRecFN_preMul_io_toPostMul_highExpB),
    .io_toPostMul_isNaN_isQuietNaNB(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB),
    .io_toPostMul_signProd(mulAddRecFN_preMul_io_toPostMul_signProd),
    .io_toPostMul_isZeroProd(mulAddRecFN_preMul_io_toPostMul_isZeroProd),
    .io_toPostMul_opSignC(mulAddRecFN_preMul_io_toPostMul_opSignC),
    .io_toPostMul_highExpC(mulAddRecFN_preMul_io_toPostMul_highExpC),
    .io_toPostMul_isNaN_isQuietNaNC(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC),
    .io_toPostMul_isCDominant(mulAddRecFN_preMul_io_toPostMul_isCDominant),
    .io_toPostMul_CAlignDist_0(mulAddRecFN_preMul_io_toPostMul_CAlignDist_0),
    .io_toPostMul_CAlignDist(mulAddRecFN_preMul_io_toPostMul_CAlignDist),
    .io_toPostMul_bit0AlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC),
    .io_toPostMul_highAlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC),
    .io_toPostMul_sExpSum(mulAddRecFN_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_roundingMode(mulAddRecFN_preMul_io_toPostMul_roundingMode)
  );
  MulAddRecFN_postMul mulAddRecFN_postMul (
    .clk(mulAddRecFN_postMul_clk),
    .reset(mulAddRecFN_postMul_reset),
    .io_fromPreMul_highExpA(mulAddRecFN_postMul_io_fromPreMul_highExpA),
    .io_fromPreMul_isNaN_isQuietNaNA(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA),
    .io_fromPreMul_highExpB(mulAddRecFN_postMul_io_fromPreMul_highExpB),
    .io_fromPreMul_isNaN_isQuietNaNB(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB),
    .io_fromPreMul_signProd(mulAddRecFN_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isZeroProd(mulAddRecFN_postMul_io_fromPreMul_isZeroProd),
    .io_fromPreMul_opSignC(mulAddRecFN_postMul_io_fromPreMul_opSignC),
    .io_fromPreMul_highExpC(mulAddRecFN_postMul_io_fromPreMul_highExpC),
    .io_fromPreMul_isNaN_isQuietNaNC(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC),
    .io_fromPreMul_isCDominant(mulAddRecFN_postMul_io_fromPreMul_isCDominant),
    .io_fromPreMul_CAlignDist_0(mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0),
    .io_fromPreMul_CAlignDist(mulAddRecFN_postMul_io_fromPreMul_CAlignDist),
    .io_fromPreMul_bit0AlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC),
    .io_fromPreMul_highAlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC),
    .io_fromPreMul_sExpSum(mulAddRecFN_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_roundingMode(mulAddRecFN_postMul_io_fromPreMul_roundingMode),
    .io_mulAddResult(mulAddRecFN_postMul_io_mulAddResult),
    .io_out(mulAddRecFN_postMul_io_out),
    .io_exceptionFlags(mulAddRecFN_postMul_io_exceptionFlags)
  );
  assign io_out = mulAddRecFN_postMul_io_out;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign mulAddRecFN_preMul_clk = clk;
  assign mulAddRecFN_preMul_reset = reset;
  assign mulAddRecFN_preMul_io_op = io_op;
  assign mulAddRecFN_preMul_io_a = io_a;
  assign mulAddRecFN_preMul_io_b = io_b;
  assign mulAddRecFN_preMul_io_c = io_c;
  assign mulAddRecFN_preMul_io_roundingMode = io_roundingMode;
  assign mulAddRecFN_postMul_clk = clk;
  assign mulAddRecFN_postMul_reset = reset;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpA = mulAddRecFN_preMul_io_toPostMul_highExpA;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpB = mulAddRecFN_preMul_io_toPostMul_highExpB;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  assign mulAddRecFN_postMul_io_fromPreMul_signProd = mulAddRecFN_preMul_io_toPostMul_signProd;
  assign mulAddRecFN_postMul_io_fromPreMul_isZeroProd = mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  assign mulAddRecFN_postMul_io_fromPreMul_opSignC = mulAddRecFN_preMul_io_toPostMul_opSignC;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpC = mulAddRecFN_preMul_io_toPostMul_highExpC;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  assign mulAddRecFN_postMul_io_fromPreMul_isCDominant = mulAddRecFN_preMul_io_toPostMul_isCDominant;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0 = mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist = mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  assign mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_sExpSum = mulAddRecFN_preMul_io_toPostMul_sExpSum;
  assign mulAddRecFN_postMul_io_fromPreMul_roundingMode = mulAddRecFN_preMul_io_toPostMul_roundingMode;
  assign mulAddRecFN_postMul_io_mulAddResult = T_11;
  assign T_7 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign T_9 = {1'h0,mulAddRecFN_preMul_io_mulAddC};
  assign GEN_0 = {{1'd0}, T_7};
  assign T_10 = GEN_0 + T_9;
  assign T_11 = T_10[48:0];
endmodule
module FPUFMAPipe(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [32:0] GEN_26;
  wire [32:0] zero;
  reg  valid;
  reg [31:0] GEN_28;
  reg [4:0] in_cmd;
  reg [31:0] GEN_29;
  reg  in_ldst;
  reg [31:0] GEN_30;
  reg  in_wen;
  reg [31:0] GEN_31;
  reg  in_ren1;
  reg [31:0] GEN_32;
  reg  in_ren2;
  reg [31:0] GEN_33;
  reg  in_ren3;
  reg [31:0] GEN_34;
  reg  in_swap12;
  reg [31:0] GEN_35;
  reg  in_swap23;
  reg [31:0] GEN_36;
  reg  in_single;
  reg [31:0] GEN_37;
  reg  in_fromint;
  reg [31:0] GEN_38;
  reg  in_toint;
  reg [31:0] GEN_39;
  reg  in_fastpipe;
  reg [31:0] GEN_40;
  reg  in_fma;
  reg [31:0] GEN_41;
  reg  in_div;
  reg [31:0] GEN_42;
  reg  in_sqrt;
  reg [31:0] GEN_43;
  reg  in_round;
  reg [31:0] GEN_44;
  reg  in_wflags;
  reg [31:0] GEN_45;
  reg [2:0] in_rm;
  reg [31:0] GEN_46;
  reg [1:0] in_typ;
  reg [31:0] GEN_47;
  reg [64:0] in_in1;
  reg [95:0] GEN_48;
  reg [64:0] in_in2;
  reg [95:0] GEN_49;
  reg [64:0] in_in3;
  reg [95:0] GEN_50;
  wire  T_179;
  wire  T_180;
  wire  T_181;
  wire  T_182;
  wire [1:0] T_183;
  wire [64:0] GEN_0;
  wire  T_186;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  fma_clk;
  wire  fma_reset;
  wire [1:0] fma_io_op;
  wire [32:0] fma_io_a;
  wire [32:0] fma_io_b;
  wire [32:0] fma_io_c;
  wire [1:0] fma_io_roundingMode;
  wire [32:0] fma_io_out;
  wire [4:0] fma_io_exceptionFlags;
  wire [64:0] res_data;
  wire [4:0] res_exc;
  wire [31:0] GEN_27;
  wire [31:0] T_193;
  wire [64:0] T_194;
  reg  T_197;
  reg [31:0] GEN_51;
  reg [64:0] T_198_data;
  reg [95:0] GEN_52;
  reg [4:0] T_198_exc;
  reg [31:0] GEN_53;
  wire [64:0] GEN_24;
  wire [4:0] GEN_25;
  wire  T_209_valid;
  wire [64:0] T_209_bits_data;
  wire [4:0] T_209_bits_exc;
  MulAddRecFN fma (
    .clk(fma_clk),
    .reset(fma_reset),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags)
  );
  assign io_out_valid = T_209_valid;
  assign io_out_bits_data = T_209_bits_data;
  assign io_out_bits_exc = T_209_bits_exc;
  assign T_131 = io_in_bits_in1[32];
  assign T_132 = io_in_bits_in2[32];
  assign T_133 = T_131 ^ T_132;
  assign GEN_26 = {{32'd0}, T_133};
  assign zero = GEN_26 << 32;
  assign T_179 = io_in_bits_cmd[1];
  assign T_180 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T_181 = T_179 & T_180;
  assign T_182 = io_in_bits_cmd[0];
  assign T_183 = {T_181,T_182};
  assign GEN_0 = io_in_bits_swap23 ? {{33'd0}, 32'h80000000} : io_in_bits_in2;
  assign T_186 = T_180 == 1'h0;
  assign GEN_1 = T_186 ? {{32'd0}, zero} : io_in_bits_in3;
  assign GEN_2 = io_in_valid ? {{3'd0}, T_183} : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_0 : in_in2;
  assign GEN_23 = io_in_valid ? GEN_1 : in_in3;
  assign fma_clk = clk;
  assign fma_reset = reset;
  assign fma_io_op = in_cmd[1:0];
  assign fma_io_a = in_in1[32:0];
  assign fma_io_b = in_in2[32:0];
  assign fma_io_c = in_in3[32:0];
  assign fma_io_roundingMode = in_rm[1:0];
  assign res_data = T_194;
  assign res_exc = fma_io_exceptionFlags;
  assign GEN_27 = $signed(32'hffffffff);
  assign T_193 = $unsigned(GEN_27);
  assign T_194 = {T_193,fma_io_out};
  assign GEN_24 = valid ? res_data : T_198_data;
  assign GEN_25 = valid ? res_exc : T_198_exc;
  assign T_209_valid = T_197;
  assign T_209_bits_data = T_198_data;
  assign T_209_bits_exc = T_198_exc;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_28 = {1{$random}};
  valid = GEN_28[0:0];
  GEN_29 = {1{$random}};
  in_cmd = GEN_29[4:0];
  GEN_30 = {1{$random}};
  in_ldst = GEN_30[0:0];
  GEN_31 = {1{$random}};
  in_wen = GEN_31[0:0];
  GEN_32 = {1{$random}};
  in_ren1 = GEN_32[0:0];
  GEN_33 = {1{$random}};
  in_ren2 = GEN_33[0:0];
  GEN_34 = {1{$random}};
  in_ren3 = GEN_34[0:0];
  GEN_35 = {1{$random}};
  in_swap12 = GEN_35[0:0];
  GEN_36 = {1{$random}};
  in_swap23 = GEN_36[0:0];
  GEN_37 = {1{$random}};
  in_single = GEN_37[0:0];
  GEN_38 = {1{$random}};
  in_fromint = GEN_38[0:0];
  GEN_39 = {1{$random}};
  in_toint = GEN_39[0:0];
  GEN_40 = {1{$random}};
  in_fastpipe = GEN_40[0:0];
  GEN_41 = {1{$random}};
  in_fma = GEN_41[0:0];
  GEN_42 = {1{$random}};
  in_div = GEN_42[0:0];
  GEN_43 = {1{$random}};
  in_sqrt = GEN_43[0:0];
  GEN_44 = {1{$random}};
  in_round = GEN_44[0:0];
  GEN_45 = {1{$random}};
  in_wflags = GEN_45[0:0];
  GEN_46 = {1{$random}};
  in_rm = GEN_46[2:0];
  GEN_47 = {1{$random}};
  in_typ = GEN_47[1:0];
  GEN_48 = {3{$random}};
  in_in1 = GEN_48[64:0];
  GEN_49 = {3{$random}};
  in_in2 = GEN_49[64:0];
  GEN_50 = {3{$random}};
  in_in3 = GEN_50[64:0];
  GEN_51 = {1{$random}};
  T_197 = GEN_51[0:0];
  GEN_52 = {3{$random}};
  T_198_data = GEN_52[64:0];
  GEN_53 = {1{$random}};
  T_198_exc = GEN_53[4:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      in_cmd <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      in_ldst <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      in_wen <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      in_ren1 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      in_ren2 <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      in_ren3 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      in_swap12 <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      in_swap23 <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      in_single <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      in_fromint <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      in_toint <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      in_fastpipe <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      in_fma <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      in_div <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      in_sqrt <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      in_round <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      in_wflags <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      in_rm <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      in_typ <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      in_in1 <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      in_in2 <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      in_in3 <= GEN_23;
    end
    if(reset) begin
      T_197 <= 1'h0;
    end else begin
      T_197 <= valid;
    end
    if(1'h0) begin
    end else begin
      T_198_data <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      T_198_exc <= GEN_25;
    end
  end
endmodule
module MulAddRecFN_preMul_92(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [1:0] io_roundingMode,
  output [52:0] io_mulAddA,
  output [52:0] io_mulAddB,
  output [105:0] io_mulAddC,
  output [2:0] io_toPostMul_highExpA,
  output  io_toPostMul_isNaN_isQuietNaNA,
  output [2:0] io_toPostMul_highExpB,
  output  io_toPostMul_isNaN_isQuietNaNB,
  output  io_toPostMul_signProd,
  output  io_toPostMul_isZeroProd,
  output  io_toPostMul_opSignC,
  output [2:0] io_toPostMul_highExpC,
  output  io_toPostMul_isNaN_isQuietNaNC,
  output  io_toPostMul_isCDominant,
  output  io_toPostMul_CAlignDist_0,
  output [7:0] io_toPostMul_CAlignDist,
  output  io_toPostMul_bit0AlignedNegSigC,
  output [54:0] io_toPostMul_highAlignedNegSigC,
  output [13:0] io_toPostMul_sExpSum,
  output [1:0] io_toPostMul_roundingMode
);
  wire  signA;
  wire [11:0] expA;
  wire [51:0] fractA;
  wire [2:0] T_42;
  wire [2:0] GEN_0;
  wire  isZeroA;
  wire  T_45;
  wire [52:0] sigA;
  wire  signB;
  wire [11:0] expB;
  wire [51:0] fractB;
  wire [2:0] T_46;
  wire  isZeroB;
  wire  T_49;
  wire [52:0] sigB;
  wire  T_50;
  wire  T_51;
  wire  opSignC;
  wire [11:0] expC;
  wire [51:0] fractC;
  wire [2:0] T_52;
  wire  isZeroC;
  wire  T_55;
  wire [52:0] sigC;
  wire  T_56;
  wire  T_57;
  wire  signProd;
  wire  isZeroProd;
  wire  T_58;
  wire  T_60;
  wire [2:0] GEN_3;
  wire [3:0] T_62;
  wire [2:0] T_63;
  wire [10:0] T_64;
  wire [13:0] T_65;
  wire [13:0] GEN_4;
  wire [14:0] T_66;
  wire [13:0] T_67;
  wire [13:0] GEN_5;
  wire [14:0] T_69;
  wire [13:0] sExpAlignedProd;
  wire  doSubMags;
  wire [13:0] GEN_6;
  wire [14:0] T_70;
  wire [13:0] sNatCAlignDist;
  wire  T_71;
  wire  CAlignDist_floor;
  wire [12:0] T_72;
  wire [12:0] GEN_7;
  wire  T_74;
  wire  CAlignDist_0;
  wire [12:0] GEN_8;
  wire  T_79;
  wire  T_80;
  wire  isCDominant;
  wire [12:0] GEN_9;
  wire  T_84;
  wire [7:0] T_85;
  wire [7:0] T_87;
  wire [7:0] CAlignDist;
  wire [13:0] sExpSum;
  wire [256:0] GEN_10;
  wire [256:0] T_89;
  wire [52:0] T_90;
  wire [31:0] T_91;
  wire [15:0] T_96;
  wire [31:0] GEN_11;
  wire [31:0] T_97;
  wire [15:0] T_98;
  wire [31:0] GEN_12;
  wire [31:0] T_99;
  wire [31:0] T_101;
  wire [31:0] T_102;
  wire [23:0] T_106;
  wire [31:0] GEN_13;
  wire [31:0] T_107;
  wire [23:0] T_108;
  wire [31:0] GEN_14;
  wire [31:0] T_109;
  wire [31:0] T_111;
  wire [31:0] T_112;
  wire [27:0] T_116;
  wire [31:0] GEN_15;
  wire [31:0] T_117;
  wire [27:0] T_118;
  wire [31:0] GEN_16;
  wire [31:0] T_119;
  wire [31:0] T_121;
  wire [31:0] T_122;
  wire [29:0] T_126;
  wire [31:0] GEN_17;
  wire [31:0] T_127;
  wire [29:0] T_128;
  wire [31:0] GEN_18;
  wire [31:0] T_129;
  wire [31:0] T_131;
  wire [31:0] T_132;
  wire [30:0] T_136;
  wire [31:0] GEN_19;
  wire [31:0] T_137;
  wire [30:0] T_138;
  wire [31:0] GEN_20;
  wire [31:0] T_139;
  wire [31:0] T_141;
  wire [31:0] T_142;
  wire [20:0] T_143;
  wire [15:0] T_144;
  wire [7:0] T_149;
  wire [15:0] GEN_21;
  wire [15:0] T_150;
  wire [7:0] T_151;
  wire [15:0] GEN_22;
  wire [15:0] T_152;
  wire [15:0] T_154;
  wire [15:0] T_155;
  wire [11:0] T_159;
  wire [15:0] GEN_23;
  wire [15:0] T_160;
  wire [11:0] T_161;
  wire [15:0] GEN_24;
  wire [15:0] T_162;
  wire [15:0] T_164;
  wire [15:0] T_165;
  wire [13:0] T_169;
  wire [15:0] GEN_25;
  wire [15:0] T_170;
  wire [13:0] T_171;
  wire [15:0] GEN_26;
  wire [15:0] T_172;
  wire [15:0] T_174;
  wire [15:0] T_175;
  wire [14:0] T_179;
  wire [15:0] GEN_27;
  wire [15:0] T_180;
  wire [14:0] T_181;
  wire [15:0] GEN_28;
  wire [15:0] T_182;
  wire [15:0] T_184;
  wire [15:0] T_185;
  wire [4:0] T_186;
  wire [3:0] T_187;
  wire [1:0] T_188;
  wire  T_189;
  wire  T_190;
  wire [1:0] T_191;
  wire [1:0] T_192;
  wire  T_193;
  wire  T_194;
  wire [1:0] T_195;
  wire [3:0] T_196;
  wire  T_197;
  wire [4:0] T_198;
  wire [20:0] T_199;
  wire [52:0] CExtraMask;
  wire [52:0] T_200;
  wire [52:0] negSigC;
  wire [107:0] GEN_29;
  wire [108:0] T_202;
  wire [107:0] T_203;
  wire [53:0] T_204;
  wire [161:0] T_205;
  wire [161:0] T_206;
  wire [161:0] T_207;
  wire [52:0] T_208;
  wire [52:0] GEN_30;
  wire  T_210;
  wire  T_211;
  wire [161:0] T_212;
  wire [162:0] T_213;
  wire [161:0] alignedNegSigC;
  wire [105:0] T_214;
  wire  T_216;
  wire  T_218;
  wire  T_220;
  wire  T_221;
  wire [54:0] T_222;
  assign io_mulAddA = sigA;
  assign io_mulAddB = sigB;
  assign io_mulAddC = T_214;
  assign io_toPostMul_highExpA = T_42;
  assign io_toPostMul_isNaN_isQuietNaNA = T_216;
  assign io_toPostMul_highExpB = T_46;
  assign io_toPostMul_isNaN_isQuietNaNB = T_218;
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroProd = isZeroProd;
  assign io_toPostMul_opSignC = opSignC;
  assign io_toPostMul_highExpC = T_52;
  assign io_toPostMul_isNaN_isQuietNaNC = T_220;
  assign io_toPostMul_isCDominant = isCDominant;
  assign io_toPostMul_CAlignDist_0 = CAlignDist_0;
  assign io_toPostMul_CAlignDist = CAlignDist;
  assign io_toPostMul_bit0AlignedNegSigC = T_221;
  assign io_toPostMul_highAlignedNegSigC = T_222;
  assign io_toPostMul_sExpSum = sExpSum;
  assign io_toPostMul_roundingMode = io_roundingMode;
  assign signA = io_a[64];
  assign expA = io_a[63:52];
  assign fractA = io_a[51:0];
  assign T_42 = expA[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZeroA = T_42 == GEN_0;
  assign T_45 = isZeroA == 1'h0;
  assign sigA = {T_45,fractA};
  assign signB = io_b[64];
  assign expB = io_b[63:52];
  assign fractB = io_b[51:0];
  assign T_46 = expB[11:9];
  assign isZeroB = T_46 == GEN_0;
  assign T_49 = isZeroB == 1'h0;
  assign sigB = {T_49,fractB};
  assign T_50 = io_c[64];
  assign T_51 = io_op[0];
  assign opSignC = T_50 ^ T_51;
  assign expC = io_c[63:52];
  assign fractC = io_c[51:0];
  assign T_52 = expC[11:9];
  assign isZeroC = T_52 == GEN_0;
  assign T_55 = isZeroC == 1'h0;
  assign sigC = {T_55,fractC};
  assign T_56 = signA ^ signB;
  assign T_57 = io_op[1];
  assign signProd = T_56 ^ T_57;
  assign isZeroProd = isZeroA | isZeroB;
  assign T_58 = expB[11];
  assign T_60 = T_58 == 1'h0;
  assign GEN_3 = {{2'd0}, T_60};
  assign T_62 = 3'h0 - GEN_3;
  assign T_63 = T_62[2:0];
  assign T_64 = expB[10:0];
  assign T_65 = {T_63,T_64};
  assign GEN_4 = {{2'd0}, expA};
  assign T_66 = GEN_4 + T_65;
  assign T_67 = T_66[13:0];
  assign GEN_5 = {{8'd0}, 6'h38};
  assign T_69 = T_67 + GEN_5;
  assign sExpAlignedProd = T_69[13:0];
  assign doSubMags = signProd ^ opSignC;
  assign GEN_6 = {{2'd0}, expC};
  assign T_70 = sExpAlignedProd - GEN_6;
  assign sNatCAlignDist = T_70[13:0];
  assign T_71 = sNatCAlignDist[13];
  assign CAlignDist_floor = isZeroProd | T_71;
  assign T_72 = sNatCAlignDist[12:0];
  assign GEN_7 = {{12'd0}, 1'h0};
  assign T_74 = T_72 == GEN_7;
  assign CAlignDist_0 = CAlignDist_floor | T_74;
  assign GEN_8 = {{7'd0}, 6'h36};
  assign T_79 = T_72 < GEN_8;
  assign T_80 = CAlignDist_floor | T_79;
  assign isCDominant = T_55 & T_80;
  assign GEN_9 = {{5'd0}, 8'ha1};
  assign T_84 = T_72 < GEN_9;
  assign T_85 = sNatCAlignDist[7:0];
  assign T_87 = T_84 ? T_85 : 8'ha1;
  assign CAlignDist = CAlignDist_floor ? {{7'd0}, 1'h0} : T_87;
  assign sExpSum = CAlignDist_floor ? {{2'd0}, expC} : sExpAlignedProd;
  assign GEN_10 = $signed(257'h10000000000000000000000000000000000000000000000000000000000000000);
  assign T_89 = $signed(GEN_10) >>> CAlignDist;
  assign T_90 = T_89[147:95];
  assign T_91 = T_90[31:0];
  assign T_96 = T_91[31:16];
  assign GEN_11 = {{16'd0}, T_96};
  assign T_97 = GEN_11 & 32'hffff;
  assign T_98 = T_91[15:0];
  assign GEN_12 = {{16'd0}, T_98};
  assign T_99 = GEN_12 << 16;
  assign T_101 = T_99 & 32'hffff0000;
  assign T_102 = T_97 | T_101;
  assign T_106 = T_102[31:8];
  assign GEN_13 = {{8'd0}, T_106};
  assign T_107 = GEN_13 & 32'hff00ff;
  assign T_108 = T_102[23:0];
  assign GEN_14 = {{8'd0}, T_108};
  assign T_109 = GEN_14 << 8;
  assign T_111 = T_109 & 32'hff00ff00;
  assign T_112 = T_107 | T_111;
  assign T_116 = T_112[31:4];
  assign GEN_15 = {{4'd0}, T_116};
  assign T_117 = GEN_15 & 32'hf0f0f0f;
  assign T_118 = T_112[27:0];
  assign GEN_16 = {{4'd0}, T_118};
  assign T_119 = GEN_16 << 4;
  assign T_121 = T_119 & 32'hf0f0f0f0;
  assign T_122 = T_117 | T_121;
  assign T_126 = T_122[31:2];
  assign GEN_17 = {{2'd0}, T_126};
  assign T_127 = GEN_17 & 32'h33333333;
  assign T_128 = T_122[29:0];
  assign GEN_18 = {{2'd0}, T_128};
  assign T_129 = GEN_18 << 2;
  assign T_131 = T_129 & 32'hcccccccc;
  assign T_132 = T_127 | T_131;
  assign T_136 = T_132[31:1];
  assign GEN_19 = {{1'd0}, T_136};
  assign T_137 = GEN_19 & 32'h55555555;
  assign T_138 = T_132[30:0];
  assign GEN_20 = {{1'd0}, T_138};
  assign T_139 = GEN_20 << 1;
  assign T_141 = T_139 & 32'haaaaaaaa;
  assign T_142 = T_137 | T_141;
  assign T_143 = T_90[52:32];
  assign T_144 = T_143[15:0];
  assign T_149 = T_144[15:8];
  assign GEN_21 = {{8'd0}, T_149};
  assign T_150 = GEN_21 & 16'hff;
  assign T_151 = T_144[7:0];
  assign GEN_22 = {{8'd0}, T_151};
  assign T_152 = GEN_22 << 8;
  assign T_154 = T_152 & 16'hff00;
  assign T_155 = T_150 | T_154;
  assign T_159 = T_155[15:4];
  assign GEN_23 = {{4'd0}, T_159};
  assign T_160 = GEN_23 & 16'hf0f;
  assign T_161 = T_155[11:0];
  assign GEN_24 = {{4'd0}, T_161};
  assign T_162 = GEN_24 << 4;
  assign T_164 = T_162 & 16'hf0f0;
  assign T_165 = T_160 | T_164;
  assign T_169 = T_165[15:2];
  assign GEN_25 = {{2'd0}, T_169};
  assign T_170 = GEN_25 & 16'h3333;
  assign T_171 = T_165[13:0];
  assign GEN_26 = {{2'd0}, T_171};
  assign T_172 = GEN_26 << 2;
  assign T_174 = T_172 & 16'hcccc;
  assign T_175 = T_170 | T_174;
  assign T_179 = T_175[15:1];
  assign GEN_27 = {{1'd0}, T_179};
  assign T_180 = GEN_27 & 16'h5555;
  assign T_181 = T_175[14:0];
  assign GEN_28 = {{1'd0}, T_181};
  assign T_182 = GEN_28 << 1;
  assign T_184 = T_182 & 16'haaaa;
  assign T_185 = T_180 | T_184;
  assign T_186 = T_143[20:16];
  assign T_187 = T_186[3:0];
  assign T_188 = T_187[1:0];
  assign T_189 = T_188[0];
  assign T_190 = T_188[1];
  assign T_191 = {T_189,T_190};
  assign T_192 = T_187[3:2];
  assign T_193 = T_192[0];
  assign T_194 = T_192[1];
  assign T_195 = {T_193,T_194};
  assign T_196 = {T_191,T_195};
  assign T_197 = T_186[4];
  assign T_198 = {T_196,T_197};
  assign T_199 = {T_185,T_198};
  assign CExtraMask = {T_142,T_199};
  assign T_200 = ~ sigC;
  assign negSigC = doSubMags ? T_200 : sigC;
  assign GEN_29 = {{107'd0}, doSubMags};
  assign T_202 = 108'h0 - GEN_29;
  assign T_203 = T_202[107:0];
  assign T_204 = {doSubMags,negSigC};
  assign T_205 = {T_204,T_203};
  assign T_206 = $signed(T_205);
  assign T_207 = $signed(T_206) >>> CAlignDist;
  assign T_208 = sigC & CExtraMask;
  assign GEN_30 = {{52'd0}, 1'h0};
  assign T_210 = T_208 != GEN_30;
  assign T_211 = T_210 ^ doSubMags;
  assign T_212 = $unsigned(T_207);
  assign T_213 = {T_212,T_211};
  assign alignedNegSigC = T_213[161:0];
  assign T_214 = alignedNegSigC[106:1];
  assign T_216 = fractA[51];
  assign T_218 = fractB[51];
  assign T_220 = fractC[51];
  assign T_221 = alignedNegSigC[0];
  assign T_222 = alignedNegSigC[161:107];
endmodule
module MulAddRecFN_postMul_93(
  input   clk,
  input   reset,
  input  [2:0] io_fromPreMul_highExpA,
  input   io_fromPreMul_isNaN_isQuietNaNA,
  input  [2:0] io_fromPreMul_highExpB,
  input   io_fromPreMul_isNaN_isQuietNaNB,
  input   io_fromPreMul_signProd,
  input   io_fromPreMul_isZeroProd,
  input   io_fromPreMul_opSignC,
  input  [2:0] io_fromPreMul_highExpC,
  input   io_fromPreMul_isNaN_isQuietNaNC,
  input   io_fromPreMul_isCDominant,
  input   io_fromPreMul_CAlignDist_0,
  input  [7:0] io_fromPreMul_CAlignDist,
  input   io_fromPreMul_bit0AlignedNegSigC,
  input  [54:0] io_fromPreMul_highAlignedNegSigC,
  input  [13:0] io_fromPreMul_sExpSum,
  input  [1:0] io_fromPreMul_roundingMode,
  input  [106:0] io_mulAddResult,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [2:0] GEN_0;
  wire  isZeroA;
  wire [1:0] T_38;
  wire  isSpecialA;
  wire  T_40;
  wire  T_42;
  wire  isInfA;
  wire  isNaNA;
  wire  T_45;
  wire  isSigNaNA;
  wire  isZeroB;
  wire [1:0] T_47;
  wire  isSpecialB;
  wire  T_49;
  wire  T_51;
  wire  isInfB;
  wire  isNaNB;
  wire  T_54;
  wire  isSigNaNB;
  wire  isZeroC;
  wire [1:0] T_56;
  wire  isSpecialC;
  wire  T_58;
  wire  T_60;
  wire  isInfC;
  wire  isNaNC;
  wire  T_63;
  wire  isSigNaNC;
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  doSubMags;
  wire  T_66;
  wire [54:0] GEN_3;
  wire [55:0] T_68;
  wire [54:0] T_69;
  wire [54:0] T_70;
  wire [105:0] T_71;
  wire [160:0] T_72;
  wire [161:0] sigSum;
  wire [107:0] T_74;
  wire [108:0] GEN_4;
  wire [108:0] T_77;
  wire [108:0] T_78;
  wire [107:0] T_80;
  wire  T_81;
  wire  T_83;
  wire  T_85;
  wire  T_87;
  wire  T_89;
  wire  T_91;
  wire  T_93;
  wire  T_95;
  wire  T_97;
  wire  T_99;
  wire  T_101;
  wire  T_103;
  wire  T_105;
  wire  T_107;
  wire  T_109;
  wire  T_111;
  wire  T_113;
  wire  T_115;
  wire  T_117;
  wire  T_119;
  wire  T_121;
  wire  T_123;
  wire  T_125;
  wire  T_127;
  wire  T_129;
  wire  T_131;
  wire  T_133;
  wire  T_135;
  wire  T_137;
  wire  T_139;
  wire  T_141;
  wire  T_143;
  wire  T_145;
  wire  T_147;
  wire  T_149;
  wire  T_151;
  wire  T_153;
  wire  T_155;
  wire  T_157;
  wire  T_159;
  wire  T_161;
  wire  T_163;
  wire  T_165;
  wire  T_167;
  wire  T_169;
  wire  T_171;
  wire  T_173;
  wire  T_175;
  wire  T_177;
  wire  T_179;
  wire  T_181;
  wire  T_183;
  wire  T_185;
  wire  T_187;
  wire  T_189;
  wire  T_191;
  wire  T_193;
  wire  T_195;
  wire  T_197;
  wire  T_199;
  wire  T_201;
  wire  T_203;
  wire  T_205;
  wire  T_207;
  wire  T_209;
  wire  T_211;
  wire  T_213;
  wire  T_215;
  wire  T_217;
  wire  T_219;
  wire  T_221;
  wire  T_223;
  wire  T_225;
  wire  T_227;
  wire  T_229;
  wire  T_231;
  wire  T_233;
  wire  T_235;
  wire  T_237;
  wire  T_239;
  wire  T_241;
  wire  T_243;
  wire  T_245;
  wire  T_247;
  wire  T_249;
  wire  T_251;
  wire  T_253;
  wire  T_255;
  wire  T_257;
  wire  T_259;
  wire  T_261;
  wire  T_263;
  wire  T_265;
  wire  T_267;
  wire  T_269;
  wire  T_271;
  wire  T_273;
  wire  T_275;
  wire  T_277;
  wire  T_279;
  wire  T_281;
  wire  T_283;
  wire  T_285;
  wire  T_287;
  wire  T_289;
  wire  T_291;
  wire  T_293;
  wire [1:0] T_295;
  wire [1:0] T_296;
  wire [2:0] T_297;
  wire [2:0] T_298;
  wire [2:0] T_299;
  wire [2:0] T_300;
  wire [3:0] T_301;
  wire [3:0] T_302;
  wire [3:0] T_303;
  wire [3:0] T_304;
  wire [3:0] T_305;
  wire [3:0] T_306;
  wire [3:0] T_307;
  wire [3:0] T_308;
  wire [4:0] T_309;
  wire [4:0] T_310;
  wire [4:0] T_311;
  wire [4:0] T_312;
  wire [4:0] T_313;
  wire [4:0] T_314;
  wire [4:0] T_315;
  wire [4:0] T_316;
  wire [4:0] T_317;
  wire [4:0] T_318;
  wire [4:0] T_319;
  wire [4:0] T_320;
  wire [4:0] T_321;
  wire [4:0] T_322;
  wire [4:0] T_323;
  wire [4:0] T_324;
  wire [5:0] T_325;
  wire [5:0] T_326;
  wire [5:0] T_327;
  wire [5:0] T_328;
  wire [5:0] T_329;
  wire [5:0] T_330;
  wire [5:0] T_331;
  wire [5:0] T_332;
  wire [5:0] T_333;
  wire [5:0] T_334;
  wire [5:0] T_335;
  wire [5:0] T_336;
  wire [5:0] T_337;
  wire [5:0] T_338;
  wire [5:0] T_339;
  wire [5:0] T_340;
  wire [5:0] T_341;
  wire [5:0] T_342;
  wire [5:0] T_343;
  wire [5:0] T_344;
  wire [5:0] T_345;
  wire [5:0] T_346;
  wire [5:0] T_347;
  wire [5:0] T_348;
  wire [5:0] T_349;
  wire [5:0] T_350;
  wire [5:0] T_351;
  wire [5:0] T_352;
  wire [5:0] T_353;
  wire [5:0] T_354;
  wire [5:0] T_355;
  wire [5:0] T_356;
  wire [6:0] T_357;
  wire [6:0] T_358;
  wire [6:0] T_359;
  wire [6:0] T_360;
  wire [6:0] T_361;
  wire [6:0] T_362;
  wire [6:0] T_363;
  wire [6:0] T_364;
  wire [6:0] T_365;
  wire [6:0] T_366;
  wire [6:0] T_367;
  wire [6:0] T_368;
  wire [6:0] T_369;
  wire [6:0] T_370;
  wire [6:0] T_371;
  wire [6:0] T_372;
  wire [6:0] T_373;
  wire [6:0] T_374;
  wire [6:0] T_375;
  wire [6:0] T_376;
  wire [6:0] T_377;
  wire [6:0] T_378;
  wire [6:0] T_379;
  wire [6:0] T_380;
  wire [6:0] T_381;
  wire [6:0] T_382;
  wire [6:0] T_383;
  wire [6:0] T_384;
  wire [6:0] T_385;
  wire [6:0] T_386;
  wire [6:0] T_387;
  wire [6:0] T_388;
  wire [6:0] T_389;
  wire [6:0] T_390;
  wire [6:0] T_391;
  wire [6:0] T_392;
  wire [6:0] T_393;
  wire [6:0] T_394;
  wire [6:0] T_395;
  wire [6:0] T_396;
  wire [6:0] T_397;
  wire [6:0] T_398;
  wire [6:0] T_399;
  wire [6:0] T_400;
  wire [7:0] GEN_6;
  wire [8:0] T_401;
  wire [7:0] estNormPos_dist;
  wire [31:0] T_402;
  wire [31:0] GEN_7;
  wire  T_404;
  wire [43:0] T_405;
  wire [43:0] GEN_8;
  wire  T_407;
  wire [1:0] firstReduceSigSum;
  wire [161:0] complSigSum;
  wire [31:0] T_408;
  wire  T_410;
  wire [43:0] T_411;
  wire  T_413;
  wire [1:0] firstReduceComplSigSum;
  wire  T_414;
  wire [7:0] GEN_11;
  wire [8:0] T_416;
  wire [7:0] T_417;
  wire [5:0] T_418;
  wire [7:0] CDom_estNormDist;
  wire  T_420;
  wire  T_421;
  wire  T_423;
  wire  T_424;
  wire [85:0] T_425;
  wire [1:0] GEN_12;
  wire  T_427;
  wire [86:0] T_428;
  wire [86:0] T_430;
  wire  T_434;
  wire [85:0] T_435;
  wire  T_436;
  wire [86:0] T_437;
  wire [86:0] T_439;
  wire [86:0] T_440;
  wire  T_444;
  wire [85:0] T_445;
  wire  T_447;
  wire [86:0] T_448;
  wire [86:0] T_450;
  wire [86:0] T_451;
  wire  T_453;
  wire [85:0] T_454;
  wire  T_455;
  wire [86:0] T_456;
  wire [86:0] T_458;
  wire [86:0] CDom_firstNormAbsSigSum;
  wire [64:0] T_459;
  wire  T_462;
  wire  T_464;
  wire [65:0] T_465;
  wire  T_467;
  wire  T_468;
  wire [85:0] GEN_14;
  wire [86:0] T_470;
  wire [85:0] T_471;
  wire [86:0] T_472;
  wire [86:0] T_473;
  wire [85:0] T_474;
  wire [10:0] T_475;
  wire [10:0] GEN_15;
  wire  T_477;
  wire [10:0] T_478;
  wire  T_480;
  wire  T_481;
  wire [86:0] T_482;
  wire  T_483;
  wire  T_484;
  wire [64:0] T_485;
  wire [21:0] GEN_17;
  wire [22:0] T_487;
  wire [21:0] T_488;
  wire [86:0] T_489;
  wire [86:0] T_490;
  wire [32:0] T_492;
  wire [53:0] GEN_18;
  wire [54:0] T_494;
  wire [53:0] T_495;
  wire [86:0] T_496;
  wire [86:0] T_497;
  wire [86:0] notCDom_pos_firstNormAbsSigSum;
  wire [63:0] T_498;
  wire [64:0] T_500;
  wire [1:0] T_503;
  wire [87:0] GEN_19;
  wire [87:0] T_504;
  wire [87:0] T_505;
  wire [86:0] T_506;
  wire  T_509;
  wire [87:0] T_510;
  wire [65:0] T_513;
  wire [87:0] GEN_21;
  wire [87:0] T_514;
  wire [87:0] T_515;
  wire [33:0] T_517;
  wire [87:0] GEN_22;
  wire [87:0] T_518;
  wire [87:0] T_519;
  wire [87:0] notCDom_neg_cFirstNormAbsSigSum;
  wire  notCDom_signSigSum;
  wire  T_521;
  wire  T_522;
  wire  doNegSignSum;
  wire [7:0] estNormDist;
  wire [87:0] T_524;
  wire [86:0] T_525;
  wire [87:0] cFirstNormAbsSigSum;
  wire  T_527;
  wire  T_529;
  wire  T_530;
  wire  doIncrSig;
  wire [4:0] estNormDist_5;
  wire [4:0] normTo2ShiftDist;
  wire [32:0] GEN_23;
  wire [32:0] T_532;
  wire [30:0] T_533;
  wire [15:0] T_534;
  wire [7:0] T_539;
  wire [15:0] GEN_24;
  wire [15:0] T_540;
  wire [7:0] T_541;
  wire [15:0] GEN_25;
  wire [15:0] T_542;
  wire [15:0] T_544;
  wire [15:0] T_545;
  wire [11:0] T_549;
  wire [15:0] GEN_26;
  wire [15:0] T_550;
  wire [11:0] T_551;
  wire [15:0] GEN_27;
  wire [15:0] T_552;
  wire [15:0] T_554;
  wire [15:0] T_555;
  wire [13:0] T_559;
  wire [15:0] GEN_28;
  wire [15:0] T_560;
  wire [13:0] T_561;
  wire [15:0] GEN_29;
  wire [15:0] T_562;
  wire [15:0] T_564;
  wire [15:0] T_565;
  wire [14:0] T_569;
  wire [15:0] GEN_30;
  wire [15:0] T_570;
  wire [14:0] T_571;
  wire [15:0] GEN_31;
  wire [15:0] T_572;
  wire [15:0] T_574;
  wire [15:0] T_575;
  wire [14:0] T_576;
  wire [7:0] T_577;
  wire [3:0] T_582;
  wire [7:0] GEN_32;
  wire [7:0] T_583;
  wire [3:0] T_584;
  wire [7:0] GEN_33;
  wire [7:0] T_585;
  wire [7:0] T_587;
  wire [7:0] T_588;
  wire [5:0] T_592;
  wire [7:0] GEN_34;
  wire [7:0] T_593;
  wire [5:0] T_594;
  wire [7:0] GEN_35;
  wire [7:0] T_595;
  wire [7:0] T_597;
  wire [7:0] T_598;
  wire [6:0] T_602;
  wire [7:0] GEN_36;
  wire [7:0] T_603;
  wire [6:0] T_604;
  wire [7:0] GEN_37;
  wire [7:0] T_605;
  wire [7:0] T_607;
  wire [7:0] T_608;
  wire [6:0] T_609;
  wire [3:0] T_610;
  wire [1:0] T_611;
  wire  T_612;
  wire  T_613;
  wire [1:0] T_614;
  wire [1:0] T_615;
  wire  T_616;
  wire  T_617;
  wire [1:0] T_618;
  wire [3:0] T_619;
  wire [2:0] T_620;
  wire [1:0] T_621;
  wire  T_622;
  wire  T_623;
  wire [1:0] T_624;
  wire  T_625;
  wire [2:0] T_626;
  wire [6:0] T_627;
  wire [14:0] T_628;
  wire [30:0] T_629;
  wire [31:0] absSigSumExtraMask;
  wire [86:0] T_631;
  wire [86:0] T_632;
  wire [31:0] T_633;
  wire [31:0] T_634;
  wire [31:0] T_635;
  wire  T_637;
  wire [31:0] T_639;
  wire  T_641;
  wire  T_642;
  wire [87:0] T_643;
  wire [56:0] sigX3;
  wire [1:0] T_644;
  wire  sigX3Shift1;
  wire [13:0] GEN_41;
  wire [14:0] T_646;
  wire [13:0] sExpX3;
  wire [2:0] T_647;
  wire  isZeroY;
  wire  T_649;
  wire  signY;
  wire [12:0] sExpX3_13;
  wire  T_650;
  wire [55:0] GEN_43;
  wire [56:0] T_652;
  wire [55:0] T_653;
  wire [12:0] T_654;
  wire [8192:0] GEN_44;
  wire [8192:0] T_656;
  wire [53:0] T_657;
  wire [31:0] T_658;
  wire [15:0] T_663;
  wire [31:0] GEN_45;
  wire [31:0] T_664;
  wire [15:0] T_665;
  wire [31:0] GEN_46;
  wire [31:0] T_666;
  wire [31:0] T_668;
  wire [31:0] T_669;
  wire [23:0] T_673;
  wire [31:0] GEN_47;
  wire [31:0] T_674;
  wire [23:0] T_675;
  wire [31:0] GEN_48;
  wire [31:0] T_676;
  wire [31:0] T_678;
  wire [31:0] T_679;
  wire [27:0] T_683;
  wire [31:0] GEN_49;
  wire [31:0] T_684;
  wire [27:0] T_685;
  wire [31:0] GEN_50;
  wire [31:0] T_686;
  wire [31:0] T_688;
  wire [31:0] T_689;
  wire [29:0] T_693;
  wire [31:0] GEN_51;
  wire [31:0] T_694;
  wire [29:0] T_695;
  wire [31:0] GEN_52;
  wire [31:0] T_696;
  wire [31:0] T_698;
  wire [31:0] T_699;
  wire [30:0] T_703;
  wire [31:0] GEN_53;
  wire [31:0] T_704;
  wire [30:0] T_705;
  wire [31:0] GEN_54;
  wire [31:0] T_706;
  wire [31:0] T_708;
  wire [31:0] T_709;
  wire [21:0] T_710;
  wire [15:0] T_711;
  wire [7:0] T_716;
  wire [15:0] GEN_55;
  wire [15:0] T_717;
  wire [7:0] T_718;
  wire [15:0] GEN_56;
  wire [15:0] T_719;
  wire [15:0] T_721;
  wire [15:0] T_722;
  wire [11:0] T_726;
  wire [15:0] GEN_57;
  wire [15:0] T_727;
  wire [11:0] T_728;
  wire [15:0] GEN_58;
  wire [15:0] T_729;
  wire [15:0] T_731;
  wire [15:0] T_732;
  wire [13:0] T_736;
  wire [15:0] GEN_59;
  wire [15:0] T_737;
  wire [13:0] T_738;
  wire [15:0] GEN_60;
  wire [15:0] T_739;
  wire [15:0] T_741;
  wire [15:0] T_742;
  wire [14:0] T_746;
  wire [15:0] GEN_61;
  wire [15:0] T_747;
  wire [14:0] T_748;
  wire [15:0] GEN_62;
  wire [15:0] T_749;
  wire [15:0] T_751;
  wire [15:0] T_752;
  wire [5:0] T_753;
  wire [3:0] T_754;
  wire [1:0] T_755;
  wire  T_756;
  wire  T_757;
  wire [1:0] T_758;
  wire [1:0] T_759;
  wire  T_760;
  wire  T_761;
  wire [1:0] T_762;
  wire [3:0] T_763;
  wire [1:0] T_764;
  wire  T_765;
  wire  T_766;
  wire [1:0] T_767;
  wire [5:0] T_768;
  wire [21:0] T_769;
  wire [53:0] T_770;
  wire  T_771;
  wire [53:0] GEN_63;
  wire [53:0] T_772;
  wire [55:0] T_774;
  wire [55:0] roundMask;
  wire [54:0] T_775;
  wire [54:0] T_776;
  wire [55:0] GEN_64;
  wire [55:0] roundPosMask;
  wire [56:0] GEN_65;
  wire [56:0] T_777;
  wire [56:0] GEN_66;
  wire  roundPosBit;
  wire [56:0] GEN_67;
  wire [56:0] T_780;
  wire  anyRoundExtra;
  wire [56:0] T_782;
  wire [56:0] T_784;
  wire  allRoundExtra;
  wire  anyRound;
  wire  allRound;
  wire  roundDirectUp;
  wire  T_787;
  wire  T_788;
  wire  T_789;
  wire  T_790;
  wire  T_793;
  wire  T_794;
  wire  T_795;
  wire  T_796;
  wire  T_797;
  wire  T_798;
  wire  T_799;
  wire  T_800;
  wire  T_801;
  wire  roundUp;
  wire  T_805;
  wire  T_806;
  wire  T_807;
  wire  T_808;
  wire  T_810;
  wire  T_811;
  wire  roundEven;
  wire  T_813;
  wire  roundInexact;
  wire [56:0] GEN_71;
  wire [56:0] T_814;
  wire [54:0] T_815;
  wire [55:0] T_817;
  wire [54:0] T_818;
  wire  T_820;
  wire  T_822;
  wire  T_823;
  wire [55:0] T_824;
  wire [56:0] GEN_73;
  wire [56:0] T_825;
  wire [54:0] T_826;
  wire [54:0] T_828;
  wire [54:0] T_830;
  wire [54:0] T_831;
  wire [54:0] T_834;
  wire [54:0] T_836;
  wire [54:0] sigY3;
  wire  T_837;
  wire [13:0] GEN_74;
  wire [14:0] T_839;
  wire [13:0] T_840;
  wire [13:0] T_842;
  wire  T_843;
  wire [13:0] T_845;
  wire [13:0] T_846;
  wire [1:0] T_847;
  wire  T_849;
  wire [14:0] T_851;
  wire [13:0] T_852;
  wire [13:0] T_854;
  wire [13:0] sExpY;
  wire [11:0] expY;
  wire [51:0] T_855;
  wire [51:0] T_856;
  wire [51:0] fractY;
  wire [2:0] T_857;
  wire [2:0] GEN_77;
  wire  overflowY;
  wire  T_860;
  wire  T_861;
  wire [11:0] GEN_78;
  wire  T_864;
  wire  T_865;
  wire  totalUnderflowY;
  wire [10:0] T_869;
  wire [12:0] GEN_79;
  wire  T_870;
  wire  T_871;
  wire  underflowY;
  wire  T_872;
  wire  T_874;
  wire  T_875;
  wire  roundMagUp;
  wire  overflowY_roundMagUp;
  wire  mulSpecial;
  wire  addSpecial;
  wire  notSpecial_addZeros;
  wire  T_877;
  wire  T_879;
  wire  commonCase;
  wire  T_880;
  wire  T_881;
  wire  T_882;
  wire  T_884;
  wire  T_886;
  wire  T_887;
  wire  T_888;
  wire  T_889;
  wire  T_890;
  wire  T_891;
  wire  notSigNaN_invalid;
  wire  T_892;
  wire  T_893;
  wire  invalid;
  wire  overflow;
  wire  underflow;
  wire  T_894;
  wire  inexact;
  wire  T_895;
  wire  notSpecial_isZeroOut;
  wire  T_896;
  wire  pegMinFiniteMagOut;
  wire  T_898;
  wire  pegMaxFiniteMagOut;
  wire  T_900;
  wire  T_901;
  wire  notNaN_isInfOut;
  wire  T_902;
  wire  T_903;
  wire  isNaNOut;
  wire  T_906;
  wire  T_908;
  wire  T_909;
  wire  T_910;
  wire  T_911;
  wire  T_913;
  wire  T_914;
  wire  T_915;
  wire  T_916;
  wire  T_919;
  wire  T_920;
  wire  T_921;
  wire  uncommonCaseSignOut;
  wire  T_923;
  wire  T_924;
  wire  T_925;
  wire  signOut;
  wire [11:0] T_928;
  wire [11:0] T_929;
  wire [11:0] T_930;
  wire [11:0] T_934;
  wire [11:0] T_935;
  wire [11:0] T_936;
  wire [11:0] T_939;
  wire [11:0] T_940;
  wire [11:0] T_941;
  wire [11:0] T_944;
  wire [11:0] T_945;
  wire [11:0] T_946;
  wire [11:0] T_949;
  wire [11:0] T_950;
  wire [11:0] T_953;
  wire [11:0] T_954;
  wire [11:0] T_957;
  wire [11:0] T_958;
  wire [11:0] T_961;
  wire [11:0] expOut;
  wire  T_962;
  wire  T_963;
  wire [51:0] T_967;
  wire [51:0] T_968;
  wire [51:0] GEN_80;
  wire [52:0] T_970;
  wire [51:0] T_971;
  wire [51:0] fractOut;
  wire [12:0] T_972;
  wire [64:0] T_973;
  wire [1:0] T_975;
  wire [1:0] T_976;
  wire [2:0] T_977;
  wire [4:0] T_978;
  assign io_out = T_973;
  assign io_exceptionFlags = T_978;
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZeroA = io_fromPreMul_highExpA == GEN_0;
  assign T_38 = io_fromPreMul_highExpA[2:1];
  assign isSpecialA = T_38 == 2'h3;
  assign T_40 = io_fromPreMul_highExpA[0];
  assign T_42 = T_40 == 1'h0;
  assign isInfA = isSpecialA & T_42;
  assign isNaNA = isSpecialA & T_40;
  assign T_45 = io_fromPreMul_isNaN_isQuietNaNA == 1'h0;
  assign isSigNaNA = isNaNA & T_45;
  assign isZeroB = io_fromPreMul_highExpB == GEN_0;
  assign T_47 = io_fromPreMul_highExpB[2:1];
  assign isSpecialB = T_47 == 2'h3;
  assign T_49 = io_fromPreMul_highExpB[0];
  assign T_51 = T_49 == 1'h0;
  assign isInfB = isSpecialB & T_51;
  assign isNaNB = isSpecialB & T_49;
  assign T_54 = io_fromPreMul_isNaN_isQuietNaNB == 1'h0;
  assign isSigNaNB = isNaNB & T_54;
  assign isZeroC = io_fromPreMul_highExpC == GEN_0;
  assign T_56 = io_fromPreMul_highExpC[2:1];
  assign isSpecialC = T_56 == 2'h3;
  assign T_58 = io_fromPreMul_highExpC[0];
  assign T_60 = T_58 == 1'h0;
  assign isInfC = isSpecialC & T_60;
  assign isNaNC = isSpecialC & T_58;
  assign T_63 = io_fromPreMul_isNaN_isQuietNaNC == 1'h0;
  assign isSigNaNC = isNaNC & T_63;
  assign roundingMode_nearest_even = io_fromPreMul_roundingMode == 2'h0;
  assign roundingMode_min = io_fromPreMul_roundingMode == 2'h2;
  assign roundingMode_max = io_fromPreMul_roundingMode == 2'h3;
  assign doSubMags = io_fromPreMul_signProd ^ io_fromPreMul_opSignC;
  assign T_66 = io_mulAddResult[106];
  assign GEN_3 = {{54'd0}, 1'h1};
  assign T_68 = io_fromPreMul_highAlignedNegSigC + GEN_3;
  assign T_69 = T_68[54:0];
  assign T_70 = T_66 ? T_69 : io_fromPreMul_highAlignedNegSigC;
  assign T_71 = io_mulAddResult[105:0];
  assign T_72 = {T_70,T_71};
  assign sigSum = {T_72,io_fromPreMul_bit0AlignedNegSigC};
  assign T_74 = sigSum[108:1];
  assign GEN_4 = {{1'd0}, T_74};
  assign T_77 = GEN_4 << 1;
  assign T_78 = GEN_4 ^ T_77;
  assign T_80 = T_78[107:0];
  assign T_81 = T_80[107];
  assign T_83 = T_80[106];
  assign T_85 = T_80[105];
  assign T_87 = T_80[104];
  assign T_89 = T_80[103];
  assign T_91 = T_80[102];
  assign T_93 = T_80[101];
  assign T_95 = T_80[100];
  assign T_97 = T_80[99];
  assign T_99 = T_80[98];
  assign T_101 = T_80[97];
  assign T_103 = T_80[96];
  assign T_105 = T_80[95];
  assign T_107 = T_80[94];
  assign T_109 = T_80[93];
  assign T_111 = T_80[92];
  assign T_113 = T_80[91];
  assign T_115 = T_80[90];
  assign T_117 = T_80[89];
  assign T_119 = T_80[88];
  assign T_121 = T_80[87];
  assign T_123 = T_80[86];
  assign T_125 = T_80[85];
  assign T_127 = T_80[84];
  assign T_129 = T_80[83];
  assign T_131 = T_80[82];
  assign T_133 = T_80[81];
  assign T_135 = T_80[80];
  assign T_137 = T_80[79];
  assign T_139 = T_80[78];
  assign T_141 = T_80[77];
  assign T_143 = T_80[76];
  assign T_145 = T_80[75];
  assign T_147 = T_80[74];
  assign T_149 = T_80[73];
  assign T_151 = T_80[72];
  assign T_153 = T_80[71];
  assign T_155 = T_80[70];
  assign T_157 = T_80[69];
  assign T_159 = T_80[68];
  assign T_161 = T_80[67];
  assign T_163 = T_80[66];
  assign T_165 = T_80[65];
  assign T_167 = T_80[64];
  assign T_169 = T_80[63];
  assign T_171 = T_80[62];
  assign T_173 = T_80[61];
  assign T_175 = T_80[60];
  assign T_177 = T_80[59];
  assign T_179 = T_80[58];
  assign T_181 = T_80[57];
  assign T_183 = T_80[56];
  assign T_185 = T_80[55];
  assign T_187 = T_80[54];
  assign T_189 = T_80[53];
  assign T_191 = T_80[52];
  assign T_193 = T_80[51];
  assign T_195 = T_80[50];
  assign T_197 = T_80[49];
  assign T_199 = T_80[48];
  assign T_201 = T_80[47];
  assign T_203 = T_80[46];
  assign T_205 = T_80[45];
  assign T_207 = T_80[44];
  assign T_209 = T_80[43];
  assign T_211 = T_80[42];
  assign T_213 = T_80[41];
  assign T_215 = T_80[40];
  assign T_217 = T_80[39];
  assign T_219 = T_80[38];
  assign T_221 = T_80[37];
  assign T_223 = T_80[36];
  assign T_225 = T_80[35];
  assign T_227 = T_80[34];
  assign T_229 = T_80[33];
  assign T_231 = T_80[32];
  assign T_233 = T_80[31];
  assign T_235 = T_80[30];
  assign T_237 = T_80[29];
  assign T_239 = T_80[28];
  assign T_241 = T_80[27];
  assign T_243 = T_80[26];
  assign T_245 = T_80[25];
  assign T_247 = T_80[24];
  assign T_249 = T_80[23];
  assign T_251 = T_80[22];
  assign T_253 = T_80[21];
  assign T_255 = T_80[20];
  assign T_257 = T_80[19];
  assign T_259 = T_80[18];
  assign T_261 = T_80[17];
  assign T_263 = T_80[16];
  assign T_265 = T_80[15];
  assign T_267 = T_80[14];
  assign T_269 = T_80[13];
  assign T_271 = T_80[12];
  assign T_273 = T_80[11];
  assign T_275 = T_80[10];
  assign T_277 = T_80[9];
  assign T_279 = T_80[8];
  assign T_281 = T_80[7];
  assign T_283 = T_80[6];
  assign T_285 = T_80[5];
  assign T_287 = T_80[4];
  assign T_289 = T_80[3];
  assign T_291 = T_80[2];
  assign T_293 = T_80[1];
  assign T_295 = T_291 ? 2'h2 : {{1'd0}, T_293};
  assign T_296 = T_289 ? 2'h3 : T_295;
  assign T_297 = T_287 ? 3'h4 : {{1'd0}, T_296};
  assign T_298 = T_285 ? 3'h5 : T_297;
  assign T_299 = T_283 ? 3'h6 : T_298;
  assign T_300 = T_281 ? 3'h7 : T_299;
  assign T_301 = T_279 ? 4'h8 : {{1'd0}, T_300};
  assign T_302 = T_277 ? 4'h9 : T_301;
  assign T_303 = T_275 ? 4'ha : T_302;
  assign T_304 = T_273 ? 4'hb : T_303;
  assign T_305 = T_271 ? 4'hc : T_304;
  assign T_306 = T_269 ? 4'hd : T_305;
  assign T_307 = T_267 ? 4'he : T_306;
  assign T_308 = T_265 ? 4'hf : T_307;
  assign T_309 = T_263 ? 5'h10 : {{1'd0}, T_308};
  assign T_310 = T_261 ? 5'h11 : T_309;
  assign T_311 = T_259 ? 5'h12 : T_310;
  assign T_312 = T_257 ? 5'h13 : T_311;
  assign T_313 = T_255 ? 5'h14 : T_312;
  assign T_314 = T_253 ? 5'h15 : T_313;
  assign T_315 = T_251 ? 5'h16 : T_314;
  assign T_316 = T_249 ? 5'h17 : T_315;
  assign T_317 = T_247 ? 5'h18 : T_316;
  assign T_318 = T_245 ? 5'h19 : T_317;
  assign T_319 = T_243 ? 5'h1a : T_318;
  assign T_320 = T_241 ? 5'h1b : T_319;
  assign T_321 = T_239 ? 5'h1c : T_320;
  assign T_322 = T_237 ? 5'h1d : T_321;
  assign T_323 = T_235 ? 5'h1e : T_322;
  assign T_324 = T_233 ? 5'h1f : T_323;
  assign T_325 = T_231 ? 6'h20 : {{1'd0}, T_324};
  assign T_326 = T_229 ? 6'h21 : T_325;
  assign T_327 = T_227 ? 6'h22 : T_326;
  assign T_328 = T_225 ? 6'h23 : T_327;
  assign T_329 = T_223 ? 6'h24 : T_328;
  assign T_330 = T_221 ? 6'h25 : T_329;
  assign T_331 = T_219 ? 6'h26 : T_330;
  assign T_332 = T_217 ? 6'h27 : T_331;
  assign T_333 = T_215 ? 6'h28 : T_332;
  assign T_334 = T_213 ? 6'h29 : T_333;
  assign T_335 = T_211 ? 6'h2a : T_334;
  assign T_336 = T_209 ? 6'h2b : T_335;
  assign T_337 = T_207 ? 6'h2c : T_336;
  assign T_338 = T_205 ? 6'h2d : T_337;
  assign T_339 = T_203 ? 6'h2e : T_338;
  assign T_340 = T_201 ? 6'h2f : T_339;
  assign T_341 = T_199 ? 6'h30 : T_340;
  assign T_342 = T_197 ? 6'h31 : T_341;
  assign T_343 = T_195 ? 6'h32 : T_342;
  assign T_344 = T_193 ? 6'h33 : T_343;
  assign T_345 = T_191 ? 6'h34 : T_344;
  assign T_346 = T_189 ? 6'h35 : T_345;
  assign T_347 = T_187 ? 6'h36 : T_346;
  assign T_348 = T_185 ? 6'h37 : T_347;
  assign T_349 = T_183 ? 6'h38 : T_348;
  assign T_350 = T_181 ? 6'h39 : T_349;
  assign T_351 = T_179 ? 6'h3a : T_350;
  assign T_352 = T_177 ? 6'h3b : T_351;
  assign T_353 = T_175 ? 6'h3c : T_352;
  assign T_354 = T_173 ? 6'h3d : T_353;
  assign T_355 = T_171 ? 6'h3e : T_354;
  assign T_356 = T_169 ? 6'h3f : T_355;
  assign T_357 = T_167 ? 7'h40 : {{1'd0}, T_356};
  assign T_358 = T_165 ? 7'h41 : T_357;
  assign T_359 = T_163 ? 7'h42 : T_358;
  assign T_360 = T_161 ? 7'h43 : T_359;
  assign T_361 = T_159 ? 7'h44 : T_360;
  assign T_362 = T_157 ? 7'h45 : T_361;
  assign T_363 = T_155 ? 7'h46 : T_362;
  assign T_364 = T_153 ? 7'h47 : T_363;
  assign T_365 = T_151 ? 7'h48 : T_364;
  assign T_366 = T_149 ? 7'h49 : T_365;
  assign T_367 = T_147 ? 7'h4a : T_366;
  assign T_368 = T_145 ? 7'h4b : T_367;
  assign T_369 = T_143 ? 7'h4c : T_368;
  assign T_370 = T_141 ? 7'h4d : T_369;
  assign T_371 = T_139 ? 7'h4e : T_370;
  assign T_372 = T_137 ? 7'h4f : T_371;
  assign T_373 = T_135 ? 7'h50 : T_372;
  assign T_374 = T_133 ? 7'h51 : T_373;
  assign T_375 = T_131 ? 7'h52 : T_374;
  assign T_376 = T_129 ? 7'h53 : T_375;
  assign T_377 = T_127 ? 7'h54 : T_376;
  assign T_378 = T_125 ? 7'h55 : T_377;
  assign T_379 = T_123 ? 7'h56 : T_378;
  assign T_380 = T_121 ? 7'h57 : T_379;
  assign T_381 = T_119 ? 7'h58 : T_380;
  assign T_382 = T_117 ? 7'h59 : T_381;
  assign T_383 = T_115 ? 7'h5a : T_382;
  assign T_384 = T_113 ? 7'h5b : T_383;
  assign T_385 = T_111 ? 7'h5c : T_384;
  assign T_386 = T_109 ? 7'h5d : T_385;
  assign T_387 = T_107 ? 7'h5e : T_386;
  assign T_388 = T_105 ? 7'h5f : T_387;
  assign T_389 = T_103 ? 7'h60 : T_388;
  assign T_390 = T_101 ? 7'h61 : T_389;
  assign T_391 = T_99 ? 7'h62 : T_390;
  assign T_392 = T_97 ? 7'h63 : T_391;
  assign T_393 = T_95 ? 7'h64 : T_392;
  assign T_394 = T_93 ? 7'h65 : T_393;
  assign T_395 = T_91 ? 7'h66 : T_394;
  assign T_396 = T_89 ? 7'h67 : T_395;
  assign T_397 = T_87 ? 7'h68 : T_396;
  assign T_398 = T_85 ? 7'h69 : T_397;
  assign T_399 = T_83 ? 7'h6a : T_398;
  assign T_400 = T_81 ? 7'h6b : T_399;
  assign GEN_6 = {{1'd0}, T_400};
  assign T_401 = 8'ha0 - GEN_6;
  assign estNormPos_dist = T_401[7:0];
  assign T_402 = sigSum[75:44];
  assign GEN_7 = {{31'd0}, 1'h0};
  assign T_404 = T_402 != GEN_7;
  assign T_405 = sigSum[43:0];
  assign GEN_8 = {{43'd0}, 1'h0};
  assign T_407 = T_405 != GEN_8;
  assign firstReduceSigSum = {T_404,T_407};
  assign complSigSum = ~ sigSum;
  assign T_408 = complSigSum[75:44];
  assign T_410 = T_408 != GEN_7;
  assign T_411 = complSigSum[43:0];
  assign T_413 = T_411 != GEN_8;
  assign firstReduceComplSigSum = {T_410,T_413};
  assign T_414 = io_fromPreMul_CAlignDist_0 | doSubMags;
  assign GEN_11 = {{7'd0}, 1'h1};
  assign T_416 = io_fromPreMul_CAlignDist - GEN_11;
  assign T_417 = T_416[7:0];
  assign T_418 = T_417[5:0];
  assign CDom_estNormDist = T_414 ? io_fromPreMul_CAlignDist : {{2'd0}, T_418};
  assign T_420 = doSubMags == 1'h0;
  assign T_421 = CDom_estNormDist[5];
  assign T_423 = T_421 == 1'h0;
  assign T_424 = T_420 & T_423;
  assign T_425 = sigSum[161:76];
  assign GEN_12 = {{1'd0}, 1'h0};
  assign T_427 = firstReduceSigSum != GEN_12;
  assign T_428 = {T_425,T_427};
  assign T_430 = T_424 ? T_428 : {{86'd0}, 1'h0};
  assign T_434 = T_420 & T_421;
  assign T_435 = sigSum[129:44];
  assign T_436 = firstReduceSigSum[0];
  assign T_437 = {T_435,T_436};
  assign T_439 = T_434 ? T_437 : {{86'd0}, 1'h0};
  assign T_440 = T_430 | T_439;
  assign T_444 = doSubMags & T_423;
  assign T_445 = complSigSum[161:76];
  assign T_447 = firstReduceComplSigSum != GEN_12;
  assign T_448 = {T_445,T_447};
  assign T_450 = T_444 ? T_448 : {{86'd0}, 1'h0};
  assign T_451 = T_440 | T_450;
  assign T_453 = doSubMags & T_421;
  assign T_454 = complSigSum[129:44];
  assign T_455 = firstReduceComplSigSum[0];
  assign T_456 = {T_454,T_455};
  assign T_458 = T_453 ? T_456 : {{86'd0}, 1'h0};
  assign CDom_firstNormAbsSigSum = T_451 | T_458;
  assign T_459 = sigSum[108:44];
  assign T_462 = T_455 == 1'h0;
  assign T_464 = doSubMags ? T_462 : T_436;
  assign T_465 = {T_459,T_464};
  assign T_467 = estNormPos_dist[4];
  assign T_468 = sigSum[1];
  assign GEN_14 = {{85'd0}, doSubMags};
  assign T_470 = 86'h0 - GEN_14;
  assign T_471 = T_470[85:0];
  assign T_472 = {T_468,T_471};
  assign T_473 = T_467 ? {{21'd0}, T_465} : T_472;
  assign T_474 = sigSum[97:12];
  assign T_475 = complSigSum[11:1];
  assign GEN_15 = {{10'd0}, 1'h0};
  assign T_477 = T_475 == GEN_15;
  assign T_478 = sigSum[11:1];
  assign T_480 = T_478 != GEN_15;
  assign T_481 = doSubMags ? T_477 : T_480;
  assign T_482 = {T_474,T_481};
  assign T_483 = estNormPos_dist[6];
  assign T_484 = estNormPos_dist[5];
  assign T_485 = sigSum[65:1];
  assign GEN_17 = {{21'd0}, doSubMags};
  assign T_487 = 22'h0 - GEN_17;
  assign T_488 = T_487[21:0];
  assign T_489 = {T_485,T_488};
  assign T_490 = T_484 ? T_489 : T_482;
  assign T_492 = sigSum[33:1];
  assign GEN_18 = {{53'd0}, doSubMags};
  assign T_494 = 54'h0 - GEN_18;
  assign T_495 = T_494[53:0];
  assign T_496 = {T_492,T_495};
  assign T_497 = T_484 ? T_473 : T_496;
  assign notCDom_pos_firstNormAbsSigSum = T_483 ? T_490 : T_497;
  assign T_498 = complSigSum[107:44];
  assign T_500 = {T_498,T_455};
  assign T_503 = complSigSum[2:1];
  assign GEN_19 = {{86'd0}, T_503};
  assign T_504 = GEN_19 << 86;
  assign T_505 = T_467 ? {{23'd0}, T_500} : T_504;
  assign T_506 = complSigSum[98:12];
  assign T_509 = T_475 != GEN_15;
  assign T_510 = {T_506,T_509};
  assign T_513 = complSigSum[66:1];
  assign GEN_21 = {{22'd0}, T_513};
  assign T_514 = GEN_21 << 22;
  assign T_515 = T_484 ? T_514 : T_510;
  assign T_517 = complSigSum[34:1];
  assign GEN_22 = {{54'd0}, T_517};
  assign T_518 = GEN_22 << 54;
  assign T_519 = T_484 ? T_505 : T_518;
  assign notCDom_neg_cFirstNormAbsSigSum = T_483 ? T_515 : T_519;
  assign notCDom_signSigSum = sigSum[109];
  assign T_521 = isZeroC == 1'h0;
  assign T_522 = doSubMags & T_521;
  assign doNegSignSum = io_fromPreMul_isCDominant ? T_522 : notCDom_signSigSum;
  assign estNormDist = io_fromPreMul_isCDominant ? CDom_estNormDist : estNormPos_dist;
  assign T_524 = io_fromPreMul_isCDominant ? {{1'd0}, CDom_firstNormAbsSigSum} : notCDom_neg_cFirstNormAbsSigSum;
  assign T_525 = io_fromPreMul_isCDominant ? CDom_firstNormAbsSigSum : notCDom_pos_firstNormAbsSigSum;
  assign cFirstNormAbsSigSum = notCDom_signSigSum ? T_524 : {{1'd0}, T_525};
  assign T_527 = io_fromPreMul_isCDominant == 1'h0;
  assign T_529 = notCDom_signSigSum == 1'h0;
  assign T_530 = T_527 & T_529;
  assign doIncrSig = T_530 & doSubMags;
  assign estNormDist_5 = estNormDist[4:0];
  assign normTo2ShiftDist = ~ estNormDist_5;
  assign GEN_23 = $signed(33'h100000000);
  assign T_532 = $signed(GEN_23) >>> normTo2ShiftDist;
  assign T_533 = T_532[31:1];
  assign T_534 = T_533[15:0];
  assign T_539 = T_534[15:8];
  assign GEN_24 = {{8'd0}, T_539};
  assign T_540 = GEN_24 & 16'hff;
  assign T_541 = T_534[7:0];
  assign GEN_25 = {{8'd0}, T_541};
  assign T_542 = GEN_25 << 8;
  assign T_544 = T_542 & 16'hff00;
  assign T_545 = T_540 | T_544;
  assign T_549 = T_545[15:4];
  assign GEN_26 = {{4'd0}, T_549};
  assign T_550 = GEN_26 & 16'hf0f;
  assign T_551 = T_545[11:0];
  assign GEN_27 = {{4'd0}, T_551};
  assign T_552 = GEN_27 << 4;
  assign T_554 = T_552 & 16'hf0f0;
  assign T_555 = T_550 | T_554;
  assign T_559 = T_555[15:2];
  assign GEN_28 = {{2'd0}, T_559};
  assign T_560 = GEN_28 & 16'h3333;
  assign T_561 = T_555[13:0];
  assign GEN_29 = {{2'd0}, T_561};
  assign T_562 = GEN_29 << 2;
  assign T_564 = T_562 & 16'hcccc;
  assign T_565 = T_560 | T_564;
  assign T_569 = T_565[15:1];
  assign GEN_30 = {{1'd0}, T_569};
  assign T_570 = GEN_30 & 16'h5555;
  assign T_571 = T_565[14:0];
  assign GEN_31 = {{1'd0}, T_571};
  assign T_572 = GEN_31 << 1;
  assign T_574 = T_572 & 16'haaaa;
  assign T_575 = T_570 | T_574;
  assign T_576 = T_533[30:16];
  assign T_577 = T_576[7:0];
  assign T_582 = T_577[7:4];
  assign GEN_32 = {{4'd0}, T_582};
  assign T_583 = GEN_32 & 8'hf;
  assign T_584 = T_577[3:0];
  assign GEN_33 = {{4'd0}, T_584};
  assign T_585 = GEN_33 << 4;
  assign T_587 = T_585 & 8'hf0;
  assign T_588 = T_583 | T_587;
  assign T_592 = T_588[7:2];
  assign GEN_34 = {{2'd0}, T_592};
  assign T_593 = GEN_34 & 8'h33;
  assign T_594 = T_588[5:0];
  assign GEN_35 = {{2'd0}, T_594};
  assign T_595 = GEN_35 << 2;
  assign T_597 = T_595 & 8'hcc;
  assign T_598 = T_593 | T_597;
  assign T_602 = T_598[7:1];
  assign GEN_36 = {{1'd0}, T_602};
  assign T_603 = GEN_36 & 8'h55;
  assign T_604 = T_598[6:0];
  assign GEN_37 = {{1'd0}, T_604};
  assign T_605 = GEN_37 << 1;
  assign T_607 = T_605 & 8'haa;
  assign T_608 = T_603 | T_607;
  assign T_609 = T_576[14:8];
  assign T_610 = T_609[3:0];
  assign T_611 = T_610[1:0];
  assign T_612 = T_611[0];
  assign T_613 = T_611[1];
  assign T_614 = {T_612,T_613};
  assign T_615 = T_610[3:2];
  assign T_616 = T_615[0];
  assign T_617 = T_615[1];
  assign T_618 = {T_616,T_617};
  assign T_619 = {T_614,T_618};
  assign T_620 = T_609[6:4];
  assign T_621 = T_620[1:0];
  assign T_622 = T_621[0];
  assign T_623 = T_621[1];
  assign T_624 = {T_622,T_623};
  assign T_625 = T_620[2];
  assign T_626 = {T_624,T_625};
  assign T_627 = {T_619,T_626};
  assign T_628 = {T_608,T_627};
  assign T_629 = {T_575,T_628};
  assign absSigSumExtraMask = {T_629,1'h1};
  assign T_631 = cFirstNormAbsSigSum[87:1];
  assign T_632 = T_631 >> normTo2ShiftDist;
  assign T_633 = cFirstNormAbsSigSum[31:0];
  assign T_634 = ~ T_633;
  assign T_635 = T_634 & absSigSumExtraMask;
  assign T_637 = T_635 == GEN_7;
  assign T_639 = T_633 & absSigSumExtraMask;
  assign T_641 = T_639 != GEN_7;
  assign T_642 = doIncrSig ? T_637 : T_641;
  assign T_643 = {T_632,T_642};
  assign sigX3 = T_643[56:0];
  assign T_644 = sigX3[56:55];
  assign sigX3Shift1 = T_644 == GEN_12;
  assign GEN_41 = {{6'd0}, estNormDist};
  assign T_646 = io_fromPreMul_sExpSum - GEN_41;
  assign sExpX3 = T_646[13:0];
  assign T_647 = sigX3[56:54];
  assign isZeroY = T_647 == GEN_0;
  assign T_649 = io_fromPreMul_signProd ^ doNegSignSum;
  assign signY = isZeroY ? roundingMode_min : T_649;
  assign sExpX3_13 = sExpX3[12:0];
  assign T_650 = sExpX3[13];
  assign GEN_43 = {{55'd0}, T_650};
  assign T_652 = 56'h0 - GEN_43;
  assign T_653 = T_652[55:0];
  assign T_654 = ~ sExpX3_13;
  assign GEN_44 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign T_656 = $signed(GEN_44) >>> T_654;
  assign T_657 = T_656[1027:974];
  assign T_658 = T_657[31:0];
  assign T_663 = T_658[31:16];
  assign GEN_45 = {{16'd0}, T_663};
  assign T_664 = GEN_45 & 32'hffff;
  assign T_665 = T_658[15:0];
  assign GEN_46 = {{16'd0}, T_665};
  assign T_666 = GEN_46 << 16;
  assign T_668 = T_666 & 32'hffff0000;
  assign T_669 = T_664 | T_668;
  assign T_673 = T_669[31:8];
  assign GEN_47 = {{8'd0}, T_673};
  assign T_674 = GEN_47 & 32'hff00ff;
  assign T_675 = T_669[23:0];
  assign GEN_48 = {{8'd0}, T_675};
  assign T_676 = GEN_48 << 8;
  assign T_678 = T_676 & 32'hff00ff00;
  assign T_679 = T_674 | T_678;
  assign T_683 = T_679[31:4];
  assign GEN_49 = {{4'd0}, T_683};
  assign T_684 = GEN_49 & 32'hf0f0f0f;
  assign T_685 = T_679[27:0];
  assign GEN_50 = {{4'd0}, T_685};
  assign T_686 = GEN_50 << 4;
  assign T_688 = T_686 & 32'hf0f0f0f0;
  assign T_689 = T_684 | T_688;
  assign T_693 = T_689[31:2];
  assign GEN_51 = {{2'd0}, T_693};
  assign T_694 = GEN_51 & 32'h33333333;
  assign T_695 = T_689[29:0];
  assign GEN_52 = {{2'd0}, T_695};
  assign T_696 = GEN_52 << 2;
  assign T_698 = T_696 & 32'hcccccccc;
  assign T_699 = T_694 | T_698;
  assign T_703 = T_699[31:1];
  assign GEN_53 = {{1'd0}, T_703};
  assign T_704 = GEN_53 & 32'h55555555;
  assign T_705 = T_699[30:0];
  assign GEN_54 = {{1'd0}, T_705};
  assign T_706 = GEN_54 << 1;
  assign T_708 = T_706 & 32'haaaaaaaa;
  assign T_709 = T_704 | T_708;
  assign T_710 = T_657[53:32];
  assign T_711 = T_710[15:0];
  assign T_716 = T_711[15:8];
  assign GEN_55 = {{8'd0}, T_716};
  assign T_717 = GEN_55 & 16'hff;
  assign T_718 = T_711[7:0];
  assign GEN_56 = {{8'd0}, T_718};
  assign T_719 = GEN_56 << 8;
  assign T_721 = T_719 & 16'hff00;
  assign T_722 = T_717 | T_721;
  assign T_726 = T_722[15:4];
  assign GEN_57 = {{4'd0}, T_726};
  assign T_727 = GEN_57 & 16'hf0f;
  assign T_728 = T_722[11:0];
  assign GEN_58 = {{4'd0}, T_728};
  assign T_729 = GEN_58 << 4;
  assign T_731 = T_729 & 16'hf0f0;
  assign T_732 = T_727 | T_731;
  assign T_736 = T_732[15:2];
  assign GEN_59 = {{2'd0}, T_736};
  assign T_737 = GEN_59 & 16'h3333;
  assign T_738 = T_732[13:0];
  assign GEN_60 = {{2'd0}, T_738};
  assign T_739 = GEN_60 << 2;
  assign T_741 = T_739 & 16'hcccc;
  assign T_742 = T_737 | T_741;
  assign T_746 = T_742[15:1];
  assign GEN_61 = {{1'd0}, T_746};
  assign T_747 = GEN_61 & 16'h5555;
  assign T_748 = T_742[14:0];
  assign GEN_62 = {{1'd0}, T_748};
  assign T_749 = GEN_62 << 1;
  assign T_751 = T_749 & 16'haaaa;
  assign T_752 = T_747 | T_751;
  assign T_753 = T_710[21:16];
  assign T_754 = T_753[3:0];
  assign T_755 = T_754[1:0];
  assign T_756 = T_755[0];
  assign T_757 = T_755[1];
  assign T_758 = {T_756,T_757};
  assign T_759 = T_754[3:2];
  assign T_760 = T_759[0];
  assign T_761 = T_759[1];
  assign T_762 = {T_760,T_761};
  assign T_763 = {T_758,T_762};
  assign T_764 = T_753[5:4];
  assign T_765 = T_764[0];
  assign T_766 = T_764[1];
  assign T_767 = {T_765,T_766};
  assign T_768 = {T_763,T_767};
  assign T_769 = {T_752,T_768};
  assign T_770 = {T_709,T_769};
  assign T_771 = sigX3[55];
  assign GEN_63 = {{53'd0}, T_771};
  assign T_772 = T_770 | GEN_63;
  assign T_774 = {T_772,2'h3};
  assign roundMask = T_653 | T_774;
  assign T_775 = roundMask[55:1];
  assign T_776 = ~ T_775;
  assign GEN_64 = {{1'd0}, T_776};
  assign roundPosMask = GEN_64 & roundMask;
  assign GEN_65 = {{1'd0}, roundPosMask};
  assign T_777 = sigX3 & GEN_65;
  assign GEN_66 = {{56'd0}, 1'h0};
  assign roundPosBit = T_777 != GEN_66;
  assign GEN_67 = {{2'd0}, T_775};
  assign T_780 = sigX3 & GEN_67;
  assign anyRoundExtra = T_780 != GEN_66;
  assign T_782 = ~ sigX3;
  assign T_784 = T_782 & GEN_67;
  assign allRoundExtra = T_784 == GEN_66;
  assign anyRound = roundPosBit | anyRoundExtra;
  assign allRound = roundPosBit & allRoundExtra;
  assign roundDirectUp = signY ? roundingMode_min : roundingMode_max;
  assign T_787 = doIncrSig == 1'h0;
  assign T_788 = T_787 & roundingMode_nearest_even;
  assign T_789 = T_788 & roundPosBit;
  assign T_790 = T_789 & anyRoundExtra;
  assign T_793 = T_787 & roundDirectUp;
  assign T_794 = T_793 & anyRound;
  assign T_795 = T_790 | T_794;
  assign T_796 = doIncrSig & allRound;
  assign T_797 = T_795 | T_796;
  assign T_798 = doIncrSig & roundingMode_nearest_even;
  assign T_799 = T_798 & roundPosBit;
  assign T_800 = T_797 | T_799;
  assign T_801 = doIncrSig & roundDirectUp;
  assign roundUp = T_800 | T_801;
  assign T_805 = roundPosBit == 1'h0;
  assign T_806 = roundingMode_nearest_even & T_805;
  assign T_807 = T_806 & allRoundExtra;
  assign T_808 = roundingMode_nearest_even & roundPosBit;
  assign T_810 = anyRoundExtra == 1'h0;
  assign T_811 = T_808 & T_810;
  assign roundEven = doIncrSig ? T_807 : T_811;
  assign T_813 = allRound == 1'h0;
  assign roundInexact = doIncrSig ? T_813 : anyRound;
  assign GEN_71 = {{1'd0}, roundMask};
  assign T_814 = sigX3 | GEN_71;
  assign T_815 = T_814[56:2];
  assign T_817 = T_815 + GEN_3;
  assign T_818 = T_817[54:0];
  assign T_820 = roundUp == 1'h0;
  assign T_822 = roundEven == 1'h0;
  assign T_823 = T_820 & T_822;
  assign T_824 = ~ roundMask;
  assign GEN_73 = {{1'd0}, T_824};
  assign T_825 = sigX3 & GEN_73;
  assign T_826 = T_825[56:2];
  assign T_828 = T_823 ? T_826 : {{54'd0}, 1'h0};
  assign T_830 = roundUp ? T_818 : {{54'd0}, 1'h0};
  assign T_831 = T_828 | T_830;
  assign T_834 = T_818 & T_776;
  assign T_836 = roundEven ? T_834 : {{54'd0}, 1'h0};
  assign sigY3 = T_831 | T_836;
  assign T_837 = sigY3[54];
  assign GEN_74 = {{13'd0}, 1'h1};
  assign T_839 = sExpX3 + GEN_74;
  assign T_840 = T_839[13:0];
  assign T_842 = T_837 ? T_840 : {{13'd0}, 1'h0};
  assign T_843 = sigY3[53];
  assign T_845 = T_843 ? sExpX3 : {{13'd0}, 1'h0};
  assign T_846 = T_842 | T_845;
  assign T_847 = sigY3[54:53];
  assign T_849 = T_847 == GEN_12;
  assign T_851 = sExpX3 - GEN_74;
  assign T_852 = T_851[13:0];
  assign T_854 = T_849 ? T_852 : {{13'd0}, 1'h0};
  assign sExpY = T_846 | T_854;
  assign expY = sExpY[11:0];
  assign T_855 = sigY3[51:0];
  assign T_856 = sigY3[52:1];
  assign fractY = sigX3Shift1 ? T_855 : T_856;
  assign T_857 = sExpY[12:10];
  assign GEN_77 = {{1'd0}, 2'h3};
  assign overflowY = T_857 == GEN_77;
  assign T_860 = isZeroY == 1'h0;
  assign T_861 = sExpY[12];
  assign GEN_78 = {{2'd0}, 10'h3ce};
  assign T_864 = expY < GEN_78;
  assign T_865 = T_861 | T_864;
  assign totalUnderflowY = T_860 & T_865;
  assign T_869 = sigX3Shift1 ? 11'h402 : 11'h401;
  assign GEN_79 = {{2'd0}, T_869};
  assign T_870 = sExpX3_13 <= GEN_79;
  assign T_871 = T_650 | T_870;
  assign underflowY = roundInexact & T_871;
  assign T_872 = roundingMode_min & signY;
  assign T_874 = signY == 1'h0;
  assign T_875 = roundingMode_max & T_874;
  assign roundMagUp = T_872 | T_875;
  assign overflowY_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign mulSpecial = isSpecialA | isSpecialB;
  assign addSpecial = mulSpecial | isSpecialC;
  assign notSpecial_addZeros = io_fromPreMul_isZeroProd & isZeroC;
  assign T_877 = addSpecial == 1'h0;
  assign T_879 = notSpecial_addZeros == 1'h0;
  assign commonCase = T_877 & T_879;
  assign T_880 = isInfA & isZeroB;
  assign T_881 = isZeroA & isInfB;
  assign T_882 = T_880 | T_881;
  assign T_884 = isNaNA == 1'h0;
  assign T_886 = isNaNB == 1'h0;
  assign T_887 = T_884 & T_886;
  assign T_888 = isInfA | isInfB;
  assign T_889 = T_887 & T_888;
  assign T_890 = T_889 & isInfC;
  assign T_891 = T_890 & doSubMags;
  assign notSigNaN_invalid = T_882 | T_891;
  assign T_892 = isSigNaNA | isSigNaNB;
  assign T_893 = T_892 | isSigNaNC;
  assign invalid = T_893 | notSigNaN_invalid;
  assign overflow = commonCase & overflowY;
  assign underflow = commonCase & underflowY;
  assign T_894 = commonCase & roundInexact;
  assign inexact = overflow | T_894;
  assign T_895 = notSpecial_addZeros | isZeroY;
  assign notSpecial_isZeroOut = T_895 | totalUnderflowY;
  assign T_896 = commonCase & totalUnderflowY;
  assign pegMinFiniteMagOut = T_896 & roundMagUp;
  assign T_898 = overflowY_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = overflow & T_898;
  assign T_900 = T_888 | isInfC;
  assign T_901 = overflow & overflowY_roundMagUp;
  assign notNaN_isInfOut = T_900 | T_901;
  assign T_902 = isNaNA | isNaNB;
  assign T_903 = T_902 | isNaNC;
  assign isNaNOut = T_903 | notSigNaN_invalid;
  assign T_906 = T_420 & io_fromPreMul_opSignC;
  assign T_908 = isSpecialC == 1'h0;
  assign T_909 = mulSpecial & T_908;
  assign T_910 = T_909 & io_fromPreMul_signProd;
  assign T_911 = T_906 | T_910;
  assign T_913 = mulSpecial == 1'h0;
  assign T_914 = T_913 & isSpecialC;
  assign T_915 = T_914 & io_fromPreMul_opSignC;
  assign T_916 = T_911 | T_915;
  assign T_919 = T_913 & notSpecial_addZeros;
  assign T_920 = T_919 & doSubMags;
  assign T_921 = T_920 & roundingMode_min;
  assign uncommonCaseSignOut = T_916 | T_921;
  assign T_923 = isNaNOut == 1'h0;
  assign T_924 = T_923 & uncommonCaseSignOut;
  assign T_925 = commonCase & signY;
  assign signOut = T_924 | T_925;
  assign T_928 = notSpecial_isZeroOut ? 12'he00 : 12'h0;
  assign T_929 = ~ T_928;
  assign T_930 = expY & T_929;
  assign T_934 = pegMinFiniteMagOut ? 12'hc31 : 12'h0;
  assign T_935 = ~ T_934;
  assign T_936 = T_930 & T_935;
  assign T_939 = pegMaxFiniteMagOut ? 12'h400 : 12'h0;
  assign T_940 = ~ T_939;
  assign T_941 = T_936 & T_940;
  assign T_944 = notNaN_isInfOut ? {{2'd0}, 10'h200} : 12'h0;
  assign T_945 = ~ T_944;
  assign T_946 = T_941 & T_945;
  assign T_949 = pegMinFiniteMagOut ? {{2'd0}, 10'h3ce} : 12'h0;
  assign T_950 = T_946 | T_949;
  assign T_953 = pegMaxFiniteMagOut ? 12'hbff : 12'h0;
  assign T_954 = T_950 | T_953;
  assign T_957 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign T_958 = T_954 | T_957;
  assign T_961 = isNaNOut ? 12'he00 : 12'h0;
  assign expOut = T_958 | T_961;
  assign T_962 = totalUnderflowY & roundMagUp;
  assign T_963 = T_962 | isNaNOut;
  assign T_967 = isNaNOut ? 52'h8000000000000 : {{51'd0}, 1'h0};
  assign T_968 = T_963 ? T_967 : fractY;
  assign GEN_80 = {{51'd0}, pegMaxFiniteMagOut};
  assign T_970 = 52'h0 - GEN_80;
  assign T_971 = T_970[51:0];
  assign fractOut = T_968 | T_971;
  assign T_972 = {signOut,expOut};
  assign T_973 = {T_972,fractOut};
  assign T_975 = {underflow,inexact};
  assign T_976 = {invalid,1'h0};
  assign T_977 = {T_976,overflow};
  assign T_978 = {T_977,T_975};
endmodule
module MulAddRecFN_91(
  input   clk,
  input   reset,
  input  [1:0] io_op,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [64:0] io_c,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  mulAddRecFN_preMul_clk;
  wire  mulAddRecFN_preMul_reset;
  wire [1:0] mulAddRecFN_preMul_io_op;
  wire [64:0] mulAddRecFN_preMul_io_a;
  wire [64:0] mulAddRecFN_preMul_io_b;
  wire [64:0] mulAddRecFN_preMul_io_c;
  wire [1:0] mulAddRecFN_preMul_io_roundingMode;
  wire [52:0] mulAddRecFN_preMul_io_mulAddA;
  wire [52:0] mulAddRecFN_preMul_io_mulAddB;
  wire [105:0] mulAddRecFN_preMul_io_mulAddC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpA;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpB;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_preMul_io_toPostMul_signProd;
  wire  mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  wire  mulAddRecFN_preMul_io_toPostMul_opSignC;
  wire [2:0] mulAddRecFN_preMul_io_toPostMul_highExpC;
  wire  mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_preMul_io_toPostMul_isCDominant;
  wire  mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  wire [7:0] mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  wire  mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  wire [54:0] mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  wire [13:0] mulAddRecFN_preMul_io_toPostMul_sExpSum;
  wire [1:0] mulAddRecFN_preMul_io_toPostMul_roundingMode;
  wire  mulAddRecFN_postMul_clk;
  wire  mulAddRecFN_postMul_reset;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpA;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpB;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB;
  wire  mulAddRecFN_postMul_io_fromPreMul_signProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_isZeroProd;
  wire  mulAddRecFN_postMul_io_fromPreMul_opSignC;
  wire [2:0] mulAddRecFN_postMul_io_fromPreMul_highExpC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC;
  wire  mulAddRecFN_postMul_io_fromPreMul_isCDominant;
  wire  mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0;
  wire [7:0] mulAddRecFN_postMul_io_fromPreMul_CAlignDist;
  wire  mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC;
  wire [54:0] mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC;
  wire [13:0] mulAddRecFN_postMul_io_fromPreMul_sExpSum;
  wire [1:0] mulAddRecFN_postMul_io_fromPreMul_roundingMode;
  wire [106:0] mulAddRecFN_postMul_io_mulAddResult;
  wire [64:0] mulAddRecFN_postMul_io_out;
  wire [4:0] mulAddRecFN_postMul_io_exceptionFlags;
  wire [105:0] T_7;
  wire [106:0] T_9;
  wire [106:0] GEN_0;
  wire [107:0] T_10;
  wire [106:0] T_11;
  MulAddRecFN_preMul_92 mulAddRecFN_preMul (
    .clk(mulAddRecFN_preMul_clk),
    .reset(mulAddRecFN_preMul_reset),
    .io_op(mulAddRecFN_preMul_io_op),
    .io_a(mulAddRecFN_preMul_io_a),
    .io_b(mulAddRecFN_preMul_io_b),
    .io_c(mulAddRecFN_preMul_io_c),
    .io_roundingMode(mulAddRecFN_preMul_io_roundingMode),
    .io_mulAddA(mulAddRecFN_preMul_io_mulAddA),
    .io_mulAddB(mulAddRecFN_preMul_io_mulAddB),
    .io_mulAddC(mulAddRecFN_preMul_io_mulAddC),
    .io_toPostMul_highExpA(mulAddRecFN_preMul_io_toPostMul_highExpA),
    .io_toPostMul_isNaN_isQuietNaNA(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA),
    .io_toPostMul_highExpB(mulAddRecFN_preMul_io_toPostMul_highExpB),
    .io_toPostMul_isNaN_isQuietNaNB(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB),
    .io_toPostMul_signProd(mulAddRecFN_preMul_io_toPostMul_signProd),
    .io_toPostMul_isZeroProd(mulAddRecFN_preMul_io_toPostMul_isZeroProd),
    .io_toPostMul_opSignC(mulAddRecFN_preMul_io_toPostMul_opSignC),
    .io_toPostMul_highExpC(mulAddRecFN_preMul_io_toPostMul_highExpC),
    .io_toPostMul_isNaN_isQuietNaNC(mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC),
    .io_toPostMul_isCDominant(mulAddRecFN_preMul_io_toPostMul_isCDominant),
    .io_toPostMul_CAlignDist_0(mulAddRecFN_preMul_io_toPostMul_CAlignDist_0),
    .io_toPostMul_CAlignDist(mulAddRecFN_preMul_io_toPostMul_CAlignDist),
    .io_toPostMul_bit0AlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC),
    .io_toPostMul_highAlignedNegSigC(mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC),
    .io_toPostMul_sExpSum(mulAddRecFN_preMul_io_toPostMul_sExpSum),
    .io_toPostMul_roundingMode(mulAddRecFN_preMul_io_toPostMul_roundingMode)
  );
  MulAddRecFN_postMul_93 mulAddRecFN_postMul (
    .clk(mulAddRecFN_postMul_clk),
    .reset(mulAddRecFN_postMul_reset),
    .io_fromPreMul_highExpA(mulAddRecFN_postMul_io_fromPreMul_highExpA),
    .io_fromPreMul_isNaN_isQuietNaNA(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA),
    .io_fromPreMul_highExpB(mulAddRecFN_postMul_io_fromPreMul_highExpB),
    .io_fromPreMul_isNaN_isQuietNaNB(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB),
    .io_fromPreMul_signProd(mulAddRecFN_postMul_io_fromPreMul_signProd),
    .io_fromPreMul_isZeroProd(mulAddRecFN_postMul_io_fromPreMul_isZeroProd),
    .io_fromPreMul_opSignC(mulAddRecFN_postMul_io_fromPreMul_opSignC),
    .io_fromPreMul_highExpC(mulAddRecFN_postMul_io_fromPreMul_highExpC),
    .io_fromPreMul_isNaN_isQuietNaNC(mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC),
    .io_fromPreMul_isCDominant(mulAddRecFN_postMul_io_fromPreMul_isCDominant),
    .io_fromPreMul_CAlignDist_0(mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0),
    .io_fromPreMul_CAlignDist(mulAddRecFN_postMul_io_fromPreMul_CAlignDist),
    .io_fromPreMul_bit0AlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC),
    .io_fromPreMul_highAlignedNegSigC(mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC),
    .io_fromPreMul_sExpSum(mulAddRecFN_postMul_io_fromPreMul_sExpSum),
    .io_fromPreMul_roundingMode(mulAddRecFN_postMul_io_fromPreMul_roundingMode),
    .io_mulAddResult(mulAddRecFN_postMul_io_mulAddResult),
    .io_out(mulAddRecFN_postMul_io_out),
    .io_exceptionFlags(mulAddRecFN_postMul_io_exceptionFlags)
  );
  assign io_out = mulAddRecFN_postMul_io_out;
  assign io_exceptionFlags = mulAddRecFN_postMul_io_exceptionFlags;
  assign mulAddRecFN_preMul_clk = clk;
  assign mulAddRecFN_preMul_reset = reset;
  assign mulAddRecFN_preMul_io_op = io_op;
  assign mulAddRecFN_preMul_io_a = io_a;
  assign mulAddRecFN_preMul_io_b = io_b;
  assign mulAddRecFN_preMul_io_c = io_c;
  assign mulAddRecFN_preMul_io_roundingMode = io_roundingMode;
  assign mulAddRecFN_postMul_clk = clk;
  assign mulAddRecFN_postMul_reset = reset;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpA = mulAddRecFN_preMul_io_toPostMul_highExpA;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNA = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNA;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpB = mulAddRecFN_preMul_io_toPostMul_highExpB;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNB = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNB;
  assign mulAddRecFN_postMul_io_fromPreMul_signProd = mulAddRecFN_preMul_io_toPostMul_signProd;
  assign mulAddRecFN_postMul_io_fromPreMul_isZeroProd = mulAddRecFN_preMul_io_toPostMul_isZeroProd;
  assign mulAddRecFN_postMul_io_fromPreMul_opSignC = mulAddRecFN_preMul_io_toPostMul_opSignC;
  assign mulAddRecFN_postMul_io_fromPreMul_highExpC = mulAddRecFN_preMul_io_toPostMul_highExpC;
  assign mulAddRecFN_postMul_io_fromPreMul_isNaN_isQuietNaNC = mulAddRecFN_preMul_io_toPostMul_isNaN_isQuietNaNC;
  assign mulAddRecFN_postMul_io_fromPreMul_isCDominant = mulAddRecFN_preMul_io_toPostMul_isCDominant;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist_0 = mulAddRecFN_preMul_io_toPostMul_CAlignDist_0;
  assign mulAddRecFN_postMul_io_fromPreMul_CAlignDist = mulAddRecFN_preMul_io_toPostMul_CAlignDist;
  assign mulAddRecFN_postMul_io_fromPreMul_bit0AlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_bit0AlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_highAlignedNegSigC = mulAddRecFN_preMul_io_toPostMul_highAlignedNegSigC;
  assign mulAddRecFN_postMul_io_fromPreMul_sExpSum = mulAddRecFN_preMul_io_toPostMul_sExpSum;
  assign mulAddRecFN_postMul_io_fromPreMul_roundingMode = mulAddRecFN_preMul_io_toPostMul_roundingMode;
  assign mulAddRecFN_postMul_io_mulAddResult = T_11;
  assign T_7 = mulAddRecFN_preMul_io_mulAddA * mulAddRecFN_preMul_io_mulAddB;
  assign T_9 = {1'h0,mulAddRecFN_preMul_io_mulAddC};
  assign GEN_0 = {{1'd0}, T_7};
  assign T_10 = GEN_0 + T_9;
  assign T_11 = T_10[106:0];
endmodule
module FPUFMAPipe_90(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  wire  T_131;
  wire  T_132;
  wire  T_133;
  wire [64:0] GEN_28;
  wire [64:0] zero;
  reg  valid;
  reg [31:0] GEN_30;
  reg [4:0] in_cmd;
  reg [31:0] GEN_31;
  reg  in_ldst;
  reg [31:0] GEN_32;
  reg  in_wen;
  reg [31:0] GEN_33;
  reg  in_ren1;
  reg [31:0] GEN_34;
  reg  in_ren2;
  reg [31:0] GEN_35;
  reg  in_ren3;
  reg [31:0] GEN_36;
  reg  in_swap12;
  reg [31:0] GEN_37;
  reg  in_swap23;
  reg [31:0] GEN_38;
  reg  in_single;
  reg [31:0] GEN_39;
  reg  in_fromint;
  reg [31:0] GEN_40;
  reg  in_toint;
  reg [31:0] GEN_41;
  reg  in_fastpipe;
  reg [31:0] GEN_42;
  reg  in_fma;
  reg [31:0] GEN_43;
  reg  in_div;
  reg [31:0] GEN_44;
  reg  in_sqrt;
  reg [31:0] GEN_45;
  reg  in_round;
  reg [31:0] GEN_46;
  reg  in_wflags;
  reg [31:0] GEN_47;
  reg [2:0] in_rm;
  reg [31:0] GEN_48;
  reg [1:0] in_typ;
  reg [31:0] GEN_49;
  reg [64:0] in_in1;
  reg [95:0] GEN_50;
  reg [64:0] in_in2;
  reg [95:0] GEN_51;
  reg [64:0] in_in3;
  reg [95:0] GEN_52;
  wire  T_179;
  wire  T_180;
  wire  T_181;
  wire  T_182;
  wire [1:0] T_183;
  wire [64:0] GEN_0;
  wire  T_186;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  fma_clk;
  wire  fma_reset;
  wire [1:0] fma_io_op;
  wire [64:0] fma_io_a;
  wire [64:0] fma_io_b;
  wire [64:0] fma_io_c;
  wire [1:0] fma_io_roundingMode;
  wire [64:0] fma_io_out;
  wire [4:0] fma_io_exceptionFlags;
  wire [64:0] res_data;
  wire [4:0] res_exc;
  wire [31:0] GEN_29;
  wire [31:0] T_193;
  wire [96:0] T_194;
  reg  T_197;
  reg [31:0] GEN_53;
  reg [64:0] T_198_data;
  reg [95:0] GEN_54;
  reg [4:0] T_198_exc;
  reg [31:0] GEN_55;
  wire [64:0] GEN_24;
  wire [4:0] GEN_25;
  reg  T_203;
  reg [31:0] GEN_56;
  reg [64:0] T_204_data;
  reg [95:0] GEN_57;
  reg [4:0] T_204_exc;
  reg [31:0] GEN_58;
  wire [64:0] GEN_26;
  wire [4:0] GEN_27;
  wire  T_215_valid;
  wire [64:0] T_215_bits_data;
  wire [4:0] T_215_bits_exc;
  MulAddRecFN_91 fma (
    .clk(fma_clk),
    .reset(fma_reset),
    .io_op(fma_io_op),
    .io_a(fma_io_a),
    .io_b(fma_io_b),
    .io_c(fma_io_c),
    .io_roundingMode(fma_io_roundingMode),
    .io_out(fma_io_out),
    .io_exceptionFlags(fma_io_exceptionFlags)
  );
  assign io_out_valid = T_215_valid;
  assign io_out_bits_data = T_215_bits_data;
  assign io_out_bits_exc = T_215_bits_exc;
  assign T_131 = io_in_bits_in1[64];
  assign T_132 = io_in_bits_in2[64];
  assign T_133 = T_131 ^ T_132;
  assign GEN_28 = {{64'd0}, T_133};
  assign zero = GEN_28 << 64;
  assign T_179 = io_in_bits_cmd[1];
  assign T_180 = io_in_bits_ren3 | io_in_bits_swap23;
  assign T_181 = T_179 & T_180;
  assign T_182 = io_in_bits_cmd[0];
  assign T_183 = {T_181,T_182};
  assign GEN_0 = io_in_bits_swap23 ? {{1'd0}, 64'h8000000000000000} : io_in_bits_in2;
  assign T_186 = T_180 == 1'h0;
  assign GEN_1 = T_186 ? zero : io_in_bits_in3;
  assign GEN_2 = io_in_valid ? {{3'd0}, T_183} : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? io_in_bits_in1 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_0 : in_in2;
  assign GEN_23 = io_in_valid ? GEN_1 : in_in3;
  assign fma_clk = clk;
  assign fma_reset = reset;
  assign fma_io_op = in_cmd[1:0];
  assign fma_io_a = in_in1;
  assign fma_io_b = in_in2;
  assign fma_io_c = in_in3;
  assign fma_io_roundingMode = in_rm[1:0];
  assign res_data = T_194[64:0];
  assign res_exc = fma_io_exceptionFlags;
  assign GEN_29 = $signed(32'hffffffff);
  assign T_193 = $unsigned(GEN_29);
  assign T_194 = {T_193,fma_io_out};
  assign GEN_24 = valid ? res_data : T_198_data;
  assign GEN_25 = valid ? res_exc : T_198_exc;
  assign GEN_26 = T_197 ? T_198_data : T_204_data;
  assign GEN_27 = T_197 ? T_198_exc : T_204_exc;
  assign T_215_valid = T_203;
  assign T_215_bits_data = T_204_data;
  assign T_215_bits_exc = T_204_exc;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_30 = {1{$random}};
  valid = GEN_30[0:0];
  GEN_31 = {1{$random}};
  in_cmd = GEN_31[4:0];
  GEN_32 = {1{$random}};
  in_ldst = GEN_32[0:0];
  GEN_33 = {1{$random}};
  in_wen = GEN_33[0:0];
  GEN_34 = {1{$random}};
  in_ren1 = GEN_34[0:0];
  GEN_35 = {1{$random}};
  in_ren2 = GEN_35[0:0];
  GEN_36 = {1{$random}};
  in_ren3 = GEN_36[0:0];
  GEN_37 = {1{$random}};
  in_swap12 = GEN_37[0:0];
  GEN_38 = {1{$random}};
  in_swap23 = GEN_38[0:0];
  GEN_39 = {1{$random}};
  in_single = GEN_39[0:0];
  GEN_40 = {1{$random}};
  in_fromint = GEN_40[0:0];
  GEN_41 = {1{$random}};
  in_toint = GEN_41[0:0];
  GEN_42 = {1{$random}};
  in_fastpipe = GEN_42[0:0];
  GEN_43 = {1{$random}};
  in_fma = GEN_43[0:0];
  GEN_44 = {1{$random}};
  in_div = GEN_44[0:0];
  GEN_45 = {1{$random}};
  in_sqrt = GEN_45[0:0];
  GEN_46 = {1{$random}};
  in_round = GEN_46[0:0];
  GEN_47 = {1{$random}};
  in_wflags = GEN_47[0:0];
  GEN_48 = {1{$random}};
  in_rm = GEN_48[2:0];
  GEN_49 = {1{$random}};
  in_typ = GEN_49[1:0];
  GEN_50 = {3{$random}};
  in_in1 = GEN_50[64:0];
  GEN_51 = {3{$random}};
  in_in2 = GEN_51[64:0];
  GEN_52 = {3{$random}};
  in_in3 = GEN_52[64:0];
  GEN_53 = {1{$random}};
  T_197 = GEN_53[0:0];
  GEN_54 = {3{$random}};
  T_198_data = GEN_54[64:0];
  GEN_55 = {1{$random}};
  T_198_exc = GEN_55[4:0];
  GEN_56 = {1{$random}};
  T_203 = GEN_56[0:0];
  GEN_57 = {3{$random}};
  T_204_data = GEN_57[64:0];
  GEN_58 = {1{$random}};
  T_204_exc = GEN_58[4:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      in_cmd <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      in_ldst <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      in_wen <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      in_ren1 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      in_ren2 <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      in_ren3 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      in_swap12 <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      in_swap23 <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      in_single <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      in_fromint <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      in_toint <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      in_fastpipe <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      in_fma <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      in_div <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      in_sqrt <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      in_round <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      in_wflags <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      in_rm <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      in_typ <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      in_in1 <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      in_in2 <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      in_in3 <= GEN_23;
    end
    if(reset) begin
      T_197 <= 1'h0;
    end else begin
      T_197 <= valid;
    end
    if(1'h0) begin
    end else begin
      T_198_data <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      T_198_exc <= GEN_25;
    end
    if(reset) begin
      T_203 <= 1'h0;
    end else begin
      T_203 <= T_197;
    end
    if(1'h0) begin
    end else begin
      T_204_data <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      T_204_exc <= GEN_27;
    end
  end
endmodule
module RecFNToRecFN(
  input   clk,
  input   reset,
  input  [32:0] io_in,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [8:0] T_4;
  wire [1:0] T_5;
  wire  T_7;
  wire  T_15_sign;
  wire  T_15_isNaN;
  wire  T_15_isInf;
  wire  T_15_isZero;
  wire [9:0] T_15_sExp;
  wire [26:0] T_15_sig;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire [2:0] T_29;
  wire [2:0] GEN_0;
  wire  T_31;
  wire [9:0] T_32;
  wire [22:0] T_34;
  wire [24:0] T_36;
  wire [26:0] T_37;
  wire [11:0] GEN_1;
  wire [11:0] GEN_2;
  wire [12:0] T_39;
  wire [11:0] T_40;
  wire [11:0] T_41;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [12:0] outRawFloat_sExp;
  wire [55:0] outRawFloat_sig;
  wire [55:0] GEN_3;
  wire [55:0] T_55;
  wire  T_56;
  wire  T_58;
  wire  invalidExc;
  wire  T_60;
  wire  T_61;
  wire [11:0] T_62;
  wire [11:0] T_65;
  wire [11:0] T_66;
  wire [11:0] T_67;
  wire  T_68;
  wire [11:0] T_71;
  wire [11:0] T_72;
  wire [11:0] T_73;
  wire [11:0] T_76;
  wire [11:0] T_77;
  wire [11:0] T_80;
  wire [11:0] T_81;
  wire [51:0] T_84;
  wire [51:0] T_85;
  wire [12:0] T_86;
  wire [64:0] T_87;
  wire [4:0] T_89;
  assign io_out = T_87;
  assign io_exceptionFlags = T_89;
  assign T_4 = io_in[31:23];
  assign T_5 = T_4[8:7];
  assign T_7 = T_5 == 2'h3;
  assign T_15_sign = T_22;
  assign T_15_isNaN = T_24;
  assign T_15_isInf = T_28;
  assign T_15_isZero = T_31;
  assign T_15_sExp = T_32;
  assign T_15_sig = T_37;
  assign T_22 = io_in[32];
  assign T_23 = T_4[6];
  assign T_24 = T_7 & T_23;
  assign T_27 = T_23 == 1'h0;
  assign T_28 = T_7 & T_27;
  assign T_29 = T_4[8:6];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_31 = T_29 == GEN_0;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_34 = io_in[22:0];
  assign T_36 = {2'h1,T_34};
  assign T_37 = {T_36,2'h0};
  assign GEN_1 = {{2{T_15_sExp[9]}},T_15_sExp};
  assign GEN_2 = $signed(12'h700);
  assign T_39 = $signed(GEN_1) + $signed(GEN_2);
  assign T_40 = T_39[11:0];
  assign T_41 = $signed(T_40);
  assign outRawFloat_sign = T_15_sign;
  assign outRawFloat_isNaN = T_15_isNaN;
  assign outRawFloat_isInf = T_15_isInf;
  assign outRawFloat_isZero = T_15_isZero;
  assign outRawFloat_sExp = {{1{T_41[11]}},T_41};
  assign outRawFloat_sig = T_55;
  assign GEN_3 = {{29'd0}, T_15_sig};
  assign T_55 = GEN_3 << 29;
  assign T_56 = outRawFloat_sig[53];
  assign T_58 = T_56 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_58;
  assign T_60 = outRawFloat_isNaN == 1'h0;
  assign T_61 = outRawFloat_sign & T_60;
  assign T_62 = outRawFloat_sExp[11:0];
  assign T_65 = outRawFloat_isZero ? 12'hc00 : {{11'd0}, 1'h0};
  assign T_66 = ~ T_65;
  assign T_67 = T_62 & T_66;
  assign T_68 = outRawFloat_isZero | outRawFloat_isInf;
  assign T_71 = T_68 ? 12'h200 : {{11'd0}, 1'h0};
  assign T_72 = ~ T_71;
  assign T_73 = T_67 & T_72;
  assign T_76 = outRawFloat_isInf ? 12'hc00 : {{11'd0}, 1'h0};
  assign T_77 = T_73 | T_76;
  assign T_80 = outRawFloat_isNaN ? 12'he00 : {{11'd0}, 1'h0};
  assign T_81 = T_77 | T_80;
  assign T_84 = outRawFloat_sig[53:2];
  assign T_85 = outRawFloat_isNaN ? 52'h8000000000000 : T_84;
  assign T_86 = {T_61,T_81};
  assign T_87 = {T_86,T_85};
  assign T_89 = {invalidExc,4'h0};
endmodule
module CompareRecFN(
  input   clk,
  input   reset,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input   io_signaling,
  output  io_lt,
  output  io_eq,
  output  io_gt,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_7;
  wire [1:0] T_8;
  wire  T_10;
  wire  rawA_sign;
  wire  rawA_isNaN;
  wire  rawA_isInf;
  wire  rawA_isZero;
  wire [12:0] rawA_sExp;
  wire [55:0] rawA_sig;
  wire  T_24;
  wire  T_25;
  wire  T_26;
  wire  T_29;
  wire  T_30;
  wire [2:0] T_31;
  wire [2:0] GEN_0;
  wire  T_33;
  wire [12:0] T_34;
  wire [51:0] T_36;
  wire [53:0] T_38;
  wire [55:0] T_39;
  wire [11:0] T_40;
  wire [1:0] T_41;
  wire  T_43;
  wire  rawB_sign;
  wire  rawB_isNaN;
  wire  rawB_isInf;
  wire  rawB_isZero;
  wire [12:0] rawB_sExp;
  wire [55:0] rawB_sig;
  wire  T_57;
  wire  T_58;
  wire  T_59;
  wire  T_62;
  wire  T_63;
  wire [2:0] T_64;
  wire  T_66;
  wire [12:0] T_67;
  wire [51:0] T_69;
  wire [53:0] T_71;
  wire [55:0] T_72;
  wire  T_74;
  wire  T_76;
  wire  ordered;
  wire  bothInfs;
  wire  bothZeros;
  wire  eqExps;
  wire  T_77;
  wire  T_78;
  wire  T_79;
  wire  common_ltMags;
  wire  T_80;
  wire  common_eqMags;
  wire  T_82;
  wire  T_84;
  wire  T_85;
  wire  T_87;
  wire  T_89;
  wire  T_90;
  wire  T_92;
  wire  T_93;
  wire  T_96;
  wire  T_97;
  wire  T_98;
  wire  T_99;
  wire  ordered_lt;
  wire  T_100;
  wire  T_101;
  wire  T_102;
  wire  ordered_eq;
  wire  T_103;
  wire  T_105;
  wire  T_106;
  wire  T_107;
  wire  T_109;
  wire  T_110;
  wire  T_111;
  wire  T_113;
  wire  T_114;
  wire  invalid;
  wire  T_115;
  wire  T_116;
  wire  T_118;
  wire  T_119;
  wire  T_121;
  wire  T_122;
  wire [4:0] T_124;
  assign io_lt = T_115;
  assign io_eq = T_116;
  assign io_gt = T_122;
  assign io_exceptionFlags = T_124;
  assign T_7 = io_a[63:52];
  assign T_8 = T_7[11:10];
  assign T_10 = T_8 == 2'h3;
  assign rawA_sign = T_24;
  assign rawA_isNaN = T_26;
  assign rawA_isInf = T_30;
  assign rawA_isZero = T_33;
  assign rawA_sExp = T_34;
  assign rawA_sig = T_39;
  assign T_24 = io_a[64];
  assign T_25 = T_7[9];
  assign T_26 = T_10 & T_25;
  assign T_29 = T_25 == 1'h0;
  assign T_30 = T_10 & T_29;
  assign T_31 = T_7[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_33 = T_31 == GEN_0;
  assign T_34 = {1'b0,$signed(T_7)};
  assign T_36 = io_a[51:0];
  assign T_38 = {2'h1,T_36};
  assign T_39 = {T_38,2'h0};
  assign T_40 = io_b[63:52];
  assign T_41 = T_40[11:10];
  assign T_43 = T_41 == 2'h3;
  assign rawB_sign = T_57;
  assign rawB_isNaN = T_59;
  assign rawB_isInf = T_63;
  assign rawB_isZero = T_66;
  assign rawB_sExp = T_67;
  assign rawB_sig = T_72;
  assign T_57 = io_b[64];
  assign T_58 = T_40[9];
  assign T_59 = T_43 & T_58;
  assign T_62 = T_58 == 1'h0;
  assign T_63 = T_43 & T_62;
  assign T_64 = T_40[11:9];
  assign T_66 = T_64 == GEN_0;
  assign T_67 = {1'b0,$signed(T_40)};
  assign T_69 = io_b[51:0];
  assign T_71 = {2'h1,T_69};
  assign T_72 = {T_71,2'h0};
  assign T_74 = rawA_isNaN == 1'h0;
  assign T_76 = rawB_isNaN == 1'h0;
  assign ordered = T_74 & T_76;
  assign bothInfs = rawA_isInf & rawB_isInf;
  assign bothZeros = rawA_isZero & rawB_isZero;
  assign eqExps = $signed(rawA_sExp) == $signed(rawB_sExp);
  assign T_77 = $signed(rawA_sExp) < $signed(rawB_sExp);
  assign T_78 = rawA_sig < rawB_sig;
  assign T_79 = eqExps & T_78;
  assign common_ltMags = T_77 | T_79;
  assign T_80 = rawA_sig == rawB_sig;
  assign common_eqMags = eqExps & T_80;
  assign T_82 = bothZeros == 1'h0;
  assign T_84 = rawB_sign == 1'h0;
  assign T_85 = rawA_sign & T_84;
  assign T_87 = bothInfs == 1'h0;
  assign T_89 = common_ltMags == 1'h0;
  assign T_90 = rawA_sign & T_89;
  assign T_92 = common_eqMags == 1'h0;
  assign T_93 = T_90 & T_92;
  assign T_96 = T_84 & common_ltMags;
  assign T_97 = T_93 | T_96;
  assign T_98 = T_87 & T_97;
  assign T_99 = T_85 | T_98;
  assign ordered_lt = T_82 & T_99;
  assign T_100 = rawA_sign == rawB_sign;
  assign T_101 = bothInfs | common_eqMags;
  assign T_102 = T_100 & T_101;
  assign ordered_eq = bothZeros | T_102;
  assign T_103 = rawA_sig[53];
  assign T_105 = T_103 == 1'h0;
  assign T_106 = rawA_isNaN & T_105;
  assign T_107 = rawB_sig[53];
  assign T_109 = T_107 == 1'h0;
  assign T_110 = rawB_isNaN & T_109;
  assign T_111 = T_106 | T_110;
  assign T_113 = ordered == 1'h0;
  assign T_114 = io_signaling & T_113;
  assign invalid = T_111 | T_114;
  assign T_115 = ordered & ordered_lt;
  assign T_116 = ordered & ordered_eq;
  assign T_118 = ordered_lt == 1'h0;
  assign T_119 = ordered & T_118;
  assign T_121 = ordered_eq == 1'h0;
  assign T_122 = T_119 & T_121;
  assign T_124 = {invalid,4'h0};
endmodule
module RecFNToIN(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  input   io_signedOut,
  output [63:0] io_out,
  output [2:0] io_intExceptionFlags
);
  wire  sign;
  wire [11:0] exp;
  wire [51:0] fract;
  wire [2:0] T_5;
  wire [2:0] GEN_0;
  wire  isZero;
  wire [1:0] T_7;
  wire  isSpecial;
  wire  T_9;
  wire  isNaN;
  wire  notSpecial_magGeOne;
  wire [52:0] T_10;
  wire [5:0] T_11;
  wire [5:0] T_13;
  wire [115:0] GEN_1;
  wire [115:0] shiftedSig;
  wire [63:0] unroundedInt;
  wire [1:0] T_14;
  wire [50:0] T_15;
  wire [50:0] GEN_2;
  wire  T_17;
  wire [2:0] roundBits;
  wire [1:0] T_18;
  wire [1:0] GEN_3;
  wire  T_20;
  wire  T_22;
  wire  roundInexact;
  wire [1:0] T_23;
  wire [1:0] T_24;
  wire  T_26;
  wire [1:0] T_28;
  wire  T_30;
  wire  T_31;
  wire [10:0] T_32;
  wire [10:0] T_33;
  wire [10:0] GEN_6;
  wire  T_35;
  wire  T_40;
  wire  roundIncr_nearestEven;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire  T_45;
  wire  T_46;
  wire  T_47;
  wire  T_49;
  wire  T_50;
  wire  T_51;
  wire  roundIncr;
  wire [63:0] T_52;
  wire [63:0] complUnroundedInt;
  wire  T_53;
  wire [63:0] GEN_8;
  wire [64:0] T_55;
  wire [63:0] T_56;
  wire [63:0] roundedInt;
  wire [61:0] T_57;
  wire [61:0] T_58;
  wire [61:0] GEN_9;
  wire  T_60;
  wire  roundCarryBut2;
  wire [10:0] GEN_10;
  wire  T_62;
  wire [10:0] GEN_11;
  wire  T_64;
  wire [62:0] T_67;
  wire [62:0] GEN_12;
  wire  T_69;
  wire  T_70;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire [10:0] GEN_13;
  wire  T_77;
  wire  T_78;
  wire  T_79;
  wire  T_80;
  wire  overflow_signed;
  wire  T_84;
  wire  T_87;
  wire  T_88;
  wire  T_89;
  wire  T_90;
  wire  T_91;
  wire  overflow_unsigned;
  wire  overflow;
  wire  T_93;
  wire  excSign;
  wire  T_94;
  wire [63:0] T_98;
  wire  T_100;
  wire  T_101;
  wire [62:0] T_104;
  wire [63:0] GEN_16;
  wire [63:0] T_105;
  wire  T_107;
  wire  T_110;
  wire [63:0] T_113;
  wire [63:0] excValue;
  wire  T_115;
  wire  T_116;
  wire  T_118;
  wire  inexact;
  wire  T_119;
  wire [63:0] T_120;
  wire [1:0] T_121;
  wire [2:0] T_122;
  assign io_out = T_120;
  assign io_intExceptionFlags = T_122;
  assign sign = io_in[64];
  assign exp = io_in[63:52];
  assign fract = io_in[51:0];
  assign T_5 = exp[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZero = T_5 == GEN_0;
  assign T_7 = exp[11:10];
  assign isSpecial = T_7 == 2'h3;
  assign T_9 = exp[9];
  assign isNaN = isSpecial & T_9;
  assign notSpecial_magGeOne = exp[11];
  assign T_10 = {notSpecial_magGeOne,fract};
  assign T_11 = exp[5:0];
  assign T_13 = notSpecial_magGeOne ? T_11 : {{5'd0}, 1'h0};
  assign GEN_1 = {{63'd0}, T_10};
  assign shiftedSig = GEN_1 << T_13;
  assign unroundedInt = shiftedSig[115:52];
  assign T_14 = shiftedSig[52:51];
  assign T_15 = shiftedSig[50:0];
  assign GEN_2 = {{50'd0}, 1'h0};
  assign T_17 = T_15 != GEN_2;
  assign roundBits = {T_14,T_17};
  assign T_18 = roundBits[1:0];
  assign GEN_3 = {{1'd0}, 1'h0};
  assign T_20 = T_18 != GEN_3;
  assign T_22 = isZero == 1'h0;
  assign roundInexact = notSpecial_magGeOne ? T_20 : T_22;
  assign T_23 = roundBits[2:1];
  assign T_24 = ~ T_23;
  assign T_26 = T_24 == GEN_3;
  assign T_28 = ~ T_18;
  assign T_30 = T_28 == GEN_3;
  assign T_31 = T_26 | T_30;
  assign T_32 = exp[10:0];
  assign T_33 = ~ T_32;
  assign GEN_6 = {{10'd0}, 1'h0};
  assign T_35 = T_33 == GEN_6;
  assign T_40 = T_35 ? T_20 : 1'h0;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T_31 : T_40;
  assign T_41 = io_roundingMode == 2'h0;
  assign T_42 = T_41 & roundIncr_nearestEven;
  assign T_43 = io_roundingMode == 2'h2;
  assign T_44 = sign & roundInexact;
  assign T_45 = T_43 & T_44;
  assign T_46 = T_42 | T_45;
  assign T_47 = io_roundingMode == 2'h3;
  assign T_49 = sign == 1'h0;
  assign T_50 = T_49 & roundInexact;
  assign T_51 = T_47 & T_50;
  assign roundIncr = T_46 | T_51;
  assign T_52 = ~ unroundedInt;
  assign complUnroundedInt = sign ? T_52 : unroundedInt;
  assign T_53 = roundIncr ^ sign;
  assign GEN_8 = {{63'd0}, 1'h1};
  assign T_55 = complUnroundedInt + GEN_8;
  assign T_56 = T_55[63:0];
  assign roundedInt = T_53 ? T_56 : complUnroundedInt;
  assign T_57 = unroundedInt[61:0];
  assign T_58 = ~ T_57;
  assign GEN_9 = {{61'd0}, 1'h0};
  assign T_60 = T_58 == GEN_9;
  assign roundCarryBut2 = T_60 & roundIncr;
  assign GEN_10 = {{4'd0}, 7'h40};
  assign T_62 = T_32 >= GEN_10;
  assign GEN_11 = {{5'd0}, 6'h3f};
  assign T_64 = T_32 == GEN_11;
  assign T_67 = unroundedInt[62:0];
  assign GEN_12 = {{62'd0}, 1'h0};
  assign T_69 = T_67 != GEN_12;
  assign T_70 = T_49 | T_69;
  assign T_71 = T_70 | roundIncr;
  assign T_72 = T_64 & T_71;
  assign T_73 = T_62 | T_72;
  assign GEN_13 = {{5'd0}, 6'h3e};
  assign T_77 = T_32 == GEN_13;
  assign T_78 = T_49 & T_77;
  assign T_79 = T_78 & roundCarryBut2;
  assign T_80 = T_73 | T_79;
  assign overflow_signed = notSpecial_magGeOne ? T_80 : 1'h0;
  assign T_84 = sign | T_62;
  assign T_87 = unroundedInt[62];
  assign T_88 = T_64 & T_87;
  assign T_89 = T_88 & roundCarryBut2;
  assign T_90 = T_84 | T_89;
  assign T_91 = sign & roundIncr;
  assign overflow_unsigned = notSpecial_magGeOne ? T_90 : T_91;
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign T_93 = isNaN == 1'h0;
  assign excSign = sign & T_93;
  assign T_94 = io_signedOut & excSign;
  assign T_98 = T_94 ? 64'h8000000000000000 : {{63'd0}, 1'h0};
  assign T_100 = excSign == 1'h0;
  assign T_101 = io_signedOut & T_100;
  assign T_104 = T_101 ? 63'h7fffffffffffffff : {{62'd0}, 1'h0};
  assign GEN_16 = {{1'd0}, T_104};
  assign T_105 = T_98 | GEN_16;
  assign T_107 = io_signedOut == 1'h0;
  assign T_110 = T_107 & T_100;
  assign T_113 = T_110 ? 64'hffffffffffffffff : {{63'd0}, 1'h0};
  assign excValue = T_105 | T_113;
  assign T_115 = isSpecial == 1'h0;
  assign T_116 = roundInexact & T_115;
  assign T_118 = overflow == 1'h0;
  assign inexact = T_116 & T_118;
  assign T_119 = isSpecial | overflow;
  assign T_120 = T_119 ? excValue : roundedInt;
  assign T_121 = {isSpecial,overflow};
  assign T_122 = {T_121,inexact};
endmodule
module RecFNToIN_95(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  input   io_signedOut,
  output [31:0] io_out,
  output [2:0] io_intExceptionFlags
);
  wire  sign;
  wire [11:0] exp;
  wire [51:0] fract;
  wire [2:0] T_5;
  wire [2:0] GEN_0;
  wire  isZero;
  wire [1:0] T_7;
  wire  isSpecial;
  wire  T_9;
  wire  isNaN;
  wire  notSpecial_magGeOne;
  wire [52:0] T_10;
  wire [4:0] T_11;
  wire [4:0] T_13;
  wire [83:0] GEN_1;
  wire [83:0] shiftedSig;
  wire [31:0] unroundedInt;
  wire [1:0] T_14;
  wire [50:0] T_15;
  wire [50:0] GEN_2;
  wire  T_17;
  wire [2:0] roundBits;
  wire [1:0] T_18;
  wire [1:0] GEN_3;
  wire  T_20;
  wire  T_22;
  wire  roundInexact;
  wire [1:0] T_23;
  wire [1:0] T_24;
  wire  T_26;
  wire [1:0] T_28;
  wire  T_30;
  wire  T_31;
  wire [10:0] T_32;
  wire [10:0] T_33;
  wire [10:0] GEN_6;
  wire  T_35;
  wire  T_40;
  wire  roundIncr_nearestEven;
  wire  T_41;
  wire  T_42;
  wire  T_43;
  wire  T_44;
  wire  T_45;
  wire  T_46;
  wire  T_47;
  wire  T_49;
  wire  T_50;
  wire  T_51;
  wire  roundIncr;
  wire [31:0] T_52;
  wire [31:0] complUnroundedInt;
  wire  T_53;
  wire [31:0] GEN_8;
  wire [32:0] T_55;
  wire [31:0] T_56;
  wire [31:0] roundedInt;
  wire [29:0] T_57;
  wire [29:0] T_58;
  wire [29:0] GEN_9;
  wire  T_60;
  wire  roundCarryBut2;
  wire [10:0] GEN_10;
  wire  T_62;
  wire [10:0] GEN_11;
  wire  T_64;
  wire [30:0] T_67;
  wire [30:0] GEN_12;
  wire  T_69;
  wire  T_70;
  wire  T_71;
  wire  T_72;
  wire  T_73;
  wire [10:0] GEN_13;
  wire  T_77;
  wire  T_78;
  wire  T_79;
  wire  T_80;
  wire  overflow_signed;
  wire  T_84;
  wire  T_87;
  wire  T_88;
  wire  T_89;
  wire  T_90;
  wire  T_91;
  wire  overflow_unsigned;
  wire  overflow;
  wire  T_93;
  wire  excSign;
  wire  T_94;
  wire [31:0] T_98;
  wire  T_100;
  wire  T_101;
  wire [30:0] T_104;
  wire [31:0] GEN_16;
  wire [31:0] T_105;
  wire  T_107;
  wire  T_110;
  wire [31:0] T_113;
  wire [31:0] excValue;
  wire  T_115;
  wire  T_116;
  wire  T_118;
  wire  inexact;
  wire  T_119;
  wire [31:0] T_120;
  wire [1:0] T_121;
  wire [2:0] T_122;
  assign io_out = T_120;
  assign io_intExceptionFlags = T_122;
  assign sign = io_in[64];
  assign exp = io_in[63:52];
  assign fract = io_in[51:0];
  assign T_5 = exp[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign isZero = T_5 == GEN_0;
  assign T_7 = exp[11:10];
  assign isSpecial = T_7 == 2'h3;
  assign T_9 = exp[9];
  assign isNaN = isSpecial & T_9;
  assign notSpecial_magGeOne = exp[11];
  assign T_10 = {notSpecial_magGeOne,fract};
  assign T_11 = exp[4:0];
  assign T_13 = notSpecial_magGeOne ? T_11 : {{4'd0}, 1'h0};
  assign GEN_1 = {{31'd0}, T_10};
  assign shiftedSig = GEN_1 << T_13;
  assign unroundedInt = shiftedSig[83:52];
  assign T_14 = shiftedSig[52:51];
  assign T_15 = shiftedSig[50:0];
  assign GEN_2 = {{50'd0}, 1'h0};
  assign T_17 = T_15 != GEN_2;
  assign roundBits = {T_14,T_17};
  assign T_18 = roundBits[1:0];
  assign GEN_3 = {{1'd0}, 1'h0};
  assign T_20 = T_18 != GEN_3;
  assign T_22 = isZero == 1'h0;
  assign roundInexact = notSpecial_magGeOne ? T_20 : T_22;
  assign T_23 = roundBits[2:1];
  assign T_24 = ~ T_23;
  assign T_26 = T_24 == GEN_3;
  assign T_28 = ~ T_18;
  assign T_30 = T_28 == GEN_3;
  assign T_31 = T_26 | T_30;
  assign T_32 = exp[10:0];
  assign T_33 = ~ T_32;
  assign GEN_6 = {{10'd0}, 1'h0};
  assign T_35 = T_33 == GEN_6;
  assign T_40 = T_35 ? T_20 : 1'h0;
  assign roundIncr_nearestEven = notSpecial_magGeOne ? T_31 : T_40;
  assign T_41 = io_roundingMode == 2'h0;
  assign T_42 = T_41 & roundIncr_nearestEven;
  assign T_43 = io_roundingMode == 2'h2;
  assign T_44 = sign & roundInexact;
  assign T_45 = T_43 & T_44;
  assign T_46 = T_42 | T_45;
  assign T_47 = io_roundingMode == 2'h3;
  assign T_49 = sign == 1'h0;
  assign T_50 = T_49 & roundInexact;
  assign T_51 = T_47 & T_50;
  assign roundIncr = T_46 | T_51;
  assign T_52 = ~ unroundedInt;
  assign complUnroundedInt = sign ? T_52 : unroundedInt;
  assign T_53 = roundIncr ^ sign;
  assign GEN_8 = {{31'd0}, 1'h1};
  assign T_55 = complUnroundedInt + GEN_8;
  assign T_56 = T_55[31:0];
  assign roundedInt = T_53 ? T_56 : complUnroundedInt;
  assign T_57 = unroundedInt[29:0];
  assign T_58 = ~ T_57;
  assign GEN_9 = {{29'd0}, 1'h0};
  assign T_60 = T_58 == GEN_9;
  assign roundCarryBut2 = T_60 & roundIncr;
  assign GEN_10 = {{5'd0}, 6'h20};
  assign T_62 = T_32 >= GEN_10;
  assign GEN_11 = {{6'd0}, 5'h1f};
  assign T_64 = T_32 == GEN_11;
  assign T_67 = unroundedInt[30:0];
  assign GEN_12 = {{30'd0}, 1'h0};
  assign T_69 = T_67 != GEN_12;
  assign T_70 = T_49 | T_69;
  assign T_71 = T_70 | roundIncr;
  assign T_72 = T_64 & T_71;
  assign T_73 = T_62 | T_72;
  assign GEN_13 = {{6'd0}, 5'h1e};
  assign T_77 = T_32 == GEN_13;
  assign T_78 = T_49 & T_77;
  assign T_79 = T_78 & roundCarryBut2;
  assign T_80 = T_73 | T_79;
  assign overflow_signed = notSpecial_magGeOne ? T_80 : 1'h0;
  assign T_84 = sign | T_62;
  assign T_87 = unroundedInt[30];
  assign T_88 = T_64 & T_87;
  assign T_89 = T_88 & roundCarryBut2;
  assign T_90 = T_84 | T_89;
  assign T_91 = sign & roundIncr;
  assign overflow_unsigned = notSpecial_magGeOne ? T_90 : T_91;
  assign overflow = io_signedOut ? overflow_signed : overflow_unsigned;
  assign T_93 = isNaN == 1'h0;
  assign excSign = sign & T_93;
  assign T_94 = io_signedOut & excSign;
  assign T_98 = T_94 ? 32'h80000000 : {{31'd0}, 1'h0};
  assign T_100 = excSign == 1'h0;
  assign T_101 = io_signedOut & T_100;
  assign T_104 = T_101 ? 31'h7fffffff : {{30'd0}, 1'h0};
  assign GEN_16 = {{1'd0}, T_104};
  assign T_105 = T_98 | GEN_16;
  assign T_107 = io_signedOut == 1'h0;
  assign T_110 = T_107 & T_100;
  assign T_113 = T_110 ? 32'hffffffff : {{31'd0}, 1'h0};
  assign excValue = T_105 | T_113;
  assign T_115 = isSpecial == 1'h0;
  assign T_116 = roundInexact & T_115;
  assign T_118 = overflow == 1'h0;
  assign inexact = T_116 & T_118;
  assign T_119 = isSpecial | overflow;
  assign T_120 = T_119 ? excValue : roundedInt;
  assign T_121 = {isSpecial,overflow};
  assign T_122 = {T_121,inexact};
endmodule
module FPToInt(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output [4:0] io_as_double_cmd,
  output  io_as_double_ldst,
  output  io_as_double_wen,
  output  io_as_double_ren1,
  output  io_as_double_ren2,
  output  io_as_double_ren3,
  output  io_as_double_swap12,
  output  io_as_double_swap23,
  output  io_as_double_single,
  output  io_as_double_fromint,
  output  io_as_double_toint,
  output  io_as_double_fastpipe,
  output  io_as_double_fma,
  output  io_as_double_div,
  output  io_as_double_sqrt,
  output  io_as_double_round,
  output  io_as_double_wflags,
  output [2:0] io_as_double_rm,
  output [1:0] io_as_double_typ,
  output [64:0] io_as_double_in1,
  output [64:0] io_as_double_in2,
  output [64:0] io_as_double_in3,
  output  io_out_valid,
  output  io_out_bits_lt,
  output [63:0] io_out_bits_store,
  output [63:0] io_out_bits_toint,
  output [4:0] io_out_bits_exc
);
  reg [4:0] in_cmd;
  reg [31:0] GEN_29;
  reg  in_ldst;
  reg [31:0] GEN_33;
  reg  in_wen;
  reg [31:0] GEN_37;
  reg  in_ren1;
  reg [31:0] GEN_38;
  reg  in_ren2;
  reg [31:0] GEN_39;
  reg  in_ren3;
  reg [31:0] GEN_43;
  reg  in_swap12;
  reg [31:0] GEN_44;
  reg  in_swap23;
  reg [31:0] GEN_45;
  reg  in_single;
  reg [31:0] GEN_46;
  reg  in_fromint;
  reg [31:0] GEN_48;
  reg  in_toint;
  reg [31:0] GEN_49;
  reg  in_fastpipe;
  reg [31:0] GEN_50;
  reg  in_fma;
  reg [31:0] GEN_51;
  reg  in_div;
  reg [31:0] GEN_52;
  reg  in_sqrt;
  reg [31:0] GEN_53;
  reg  in_round;
  reg [31:0] GEN_54;
  reg  in_wflags;
  reg [31:0] GEN_56;
  reg [2:0] in_rm;
  reg [31:0] GEN_57;
  reg [1:0] in_typ;
  reg [31:0] GEN_59;
  reg [64:0] in_in1;
  reg [95:0] GEN_62;
  reg [64:0] in_in2;
  reg [95:0] GEN_63;
  reg [64:0] in_in3;
  reg [95:0] GEN_64;
  reg  valid;
  reg [31:0] GEN_65;
  wire  RecFNToRecFN_227_clk;
  wire  RecFNToRecFN_227_reset;
  wire [32:0] RecFNToRecFN_227_io_in;
  wire [1:0] RecFNToRecFN_227_io_roundingMode;
  wire [64:0] RecFNToRecFN_227_io_out;
  wire [4:0] RecFNToRecFN_227_io_exceptionFlags;
  wire  RecFNToRecFN_94_229_clk;
  wire  RecFNToRecFN_94_229_reset;
  wire [32:0] RecFNToRecFN_94_229_io_in;
  wire [1:0] RecFNToRecFN_94_229_io_roundingMode;
  wire [64:0] RecFNToRecFN_94_229_io_out;
  wire [4:0] RecFNToRecFN_94_229_io_exceptionFlags;
  wire  T_232;
  wire  T_233;
  wire [4:0] GEN_28;
  wire [4:0] T_236;
  wire  T_237;
  wire  T_239;
  wire  T_240;
  wire [64:0] GEN_0;
  wire [64:0] GEN_1;
  wire [4:0] GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire [2:0] GEN_19;
  wire [1:0] GEN_20;
  wire [64:0] GEN_21;
  wire [64:0] GEN_22;
  wire [64:0] GEN_23;
  wire  T_241;
  wire [8:0] T_242;
  wire [22:0] T_243;
  wire [6:0] T_244;
  wire [6:0] GEN_30;
  wire  T_246;
  wire [2:0] T_247;
  wire [2:0] GEN_31;
  wire  T_249;
  wire [1:0] T_250;
  wire [1:0] GEN_32;
  wire  T_252;
  wire  T_253;
  wire  T_254;
  wire  T_259;
  wire  T_260;
  wire  T_263;
  wire  T_264;
  wire  T_267;
  wire  T_268;
  wire  T_269;
  wire [4:0] T_271;
  wire [4:0] GEN_34;
  wire [5:0] T_272;
  wire [4:0] T_273;
  wire [23:0] T_275;
  wire [23:0] T_276;
  wire [22:0] T_277;
  wire [7:0] T_278;
  wire [8:0] T_280;
  wire [7:0] T_281;
  wire [7:0] GEN_35;
  wire [8:0] T_283;
  wire [7:0] T_284;
  wire [7:0] T_285;
  wire  T_286;
  wire [22:0] T_288;
  wire [22:0] T_289;
  wire [8:0] T_290;
  wire [31:0] unrec_s;
  wire  T_291;
  wire [11:0] T_292;
  wire [51:0] T_293;
  wire [9:0] T_294;
  wire [9:0] GEN_36;
  wire  T_296;
  wire [2:0] T_297;
  wire  T_299;
  wire [1:0] T_300;
  wire  T_302;
  wire  T_303;
  wire  T_304;
  wire  T_309;
  wire  T_310;
  wire  T_313;
  wire  T_314;
  wire  T_317;
  wire  T_318;
  wire  T_319;
  wire [5:0] T_321;
  wire [5:0] GEN_40;
  wire [6:0] T_322;
  wire [5:0] T_323;
  wire [52:0] T_325;
  wire [52:0] T_326;
  wire [51:0] T_327;
  wire [10:0] T_328;
  wire [11:0] T_330;
  wire [10:0] T_331;
  wire [10:0] GEN_41;
  wire [11:0] T_333;
  wire [10:0] T_334;
  wire [10:0] T_335;
  wire  T_336;
  wire [51:0] T_338;
  wire [51:0] T_339;
  wire [11:0] T_340;
  wire [63:0] unrec_d;
  wire  T_341;
  wire [31:0] GEN_42;
  wire [32:0] T_343;
  wire [31:0] T_344;
  wire [63:0] T_345;
  wire [63:0] unrec_out;
  wire [1:0] T_350;
  wire  T_352;
  wire  T_359;
  wire  T_360;
  wire  T_361;
  wire  T_366;
  wire  T_368;
  wire  T_369;
  wire [2:0] GEN_47;
  wire  T_371;
  wire  T_374;
  wire  T_375;
  wire [2:0] T_376;
  wire  T_378;
  wire  T_379;
  wire  T_381;
  wire  T_382;
  wire  T_384;
  wire  T_386;
  wire  T_387;
  wire  T_390;
  wire  T_393;
  wire  T_396;
  wire  T_397;
  wire  T_398;
  wire  T_399;
  wire  T_400;
  wire [1:0] T_401;
  wire [1:0] T_402;
  wire [2:0] T_403;
  wire [4:0] T_404;
  wire [1:0] T_405;
  wire [1:0] T_406;
  wire [2:0] T_407;
  wire [4:0] T_408;
  wire [9:0] classify_s;
  wire [1:0] T_413;
  wire  T_415;
  wire  T_422;
  wire  T_423;
  wire  T_424;
  wire  T_429;
  wire  T_431;
  wire  T_432;
  wire  T_434;
  wire  T_437;
  wire  T_438;
  wire [2:0] T_439;
  wire  T_441;
  wire  T_442;
  wire  T_444;
  wire  T_445;
  wire  T_447;
  wire  T_449;
  wire  T_450;
  wire  T_453;
  wire  T_456;
  wire  T_459;
  wire  T_460;
  wire  T_461;
  wire  T_462;
  wire  T_463;
  wire [1:0] T_464;
  wire [1:0] T_465;
  wire [2:0] T_466;
  wire [4:0] T_467;
  wire [1:0] T_468;
  wire [1:0] T_469;
  wire [2:0] T_470;
  wire [4:0] T_471;
  wire [9:0] classify_d;
  wire [9:0] classify_out;
  wire  dcmp_clk;
  wire  dcmp_reset;
  wire [64:0] dcmp_io_a;
  wire [64:0] dcmp_io_b;
  wire  dcmp_io_signaling;
  wire  dcmp_io_lt;
  wire  dcmp_io_eq;
  wire  dcmp_io_gt;
  wire [4:0] dcmp_io_exceptionFlags;
  wire [2:0] T_473;
  wire [1:0] T_474;
  wire [2:0] GEN_55;
  wire [2:0] T_475;
  wire  dcmp_out;
  wire  d2l_clk;
  wire  d2l_reset;
  wire [64:0] d2l_io_in;
  wire [1:0] d2l_io_roundingMode;
  wire  d2l_io_signedOut;
  wire [63:0] d2l_io_out;
  wire [2:0] d2l_io_intExceptionFlags;
  wire  d2w_clk;
  wire  d2w_reset;
  wire [64:0] d2w_io_in;
  wire [1:0] d2w_io_roundingMode;
  wire  d2w_io_signedOut;
  wire [31:0] d2w_io_out;
  wire [2:0] d2w_io_intExceptionFlags;
  wire  T_477;
  wire  T_478;
  wire  T_481;
  wire [63:0] T_482;
  wire [4:0] T_486;
  wire [4:0] GEN_58;
  wire  T_487;
  wire [63:0] GEN_24;
  wire [4:0] GEN_25;
  wire [4:0] GEN_60;
  wire  T_491;
  wire  T_492;
  wire [63:0] T_493;
  wire [31:0] T_494;
  wire [63:0] T_495;
  wire [63:0] T_496;
  wire [2:0] T_498;
  wire [1:0] T_499;
  wire [1:0] GEN_61;
  wire  T_501;
  wire  T_503;
  wire [3:0] T_504;
  wire [4:0] T_505;
  wire [63:0] GEN_26;
  wire [4:0] GEN_27;
  RecFNToRecFN RecFNToRecFN_227 (
    .clk(RecFNToRecFN_227_clk),
    .reset(RecFNToRecFN_227_reset),
    .io_in(RecFNToRecFN_227_io_in),
    .io_roundingMode(RecFNToRecFN_227_io_roundingMode),
    .io_out(RecFNToRecFN_227_io_out),
    .io_exceptionFlags(RecFNToRecFN_227_io_exceptionFlags)
  );
  RecFNToRecFN RecFNToRecFN_94_229 (
    .clk(RecFNToRecFN_94_229_clk),
    .reset(RecFNToRecFN_94_229_reset),
    .io_in(RecFNToRecFN_94_229_io_in),
    .io_roundingMode(RecFNToRecFN_94_229_io_roundingMode),
    .io_out(RecFNToRecFN_94_229_io_out),
    .io_exceptionFlags(RecFNToRecFN_94_229_io_exceptionFlags)
  );
  CompareRecFN dcmp (
    .clk(dcmp_clk),
    .reset(dcmp_reset),
    .io_a(dcmp_io_a),
    .io_b(dcmp_io_b),
    .io_signaling(dcmp_io_signaling),
    .io_lt(dcmp_io_lt),
    .io_eq(dcmp_io_eq),
    .io_gt(dcmp_io_gt),
    .io_exceptionFlags(dcmp_io_exceptionFlags)
  );
  RecFNToIN d2l (
    .clk(d2l_clk),
    .reset(d2l_reset),
    .io_in(d2l_io_in),
    .io_roundingMode(d2l_io_roundingMode),
    .io_signedOut(d2l_io_signedOut),
    .io_out(d2l_io_out),
    .io_intExceptionFlags(d2l_io_intExceptionFlags)
  );
  RecFNToIN_95 d2w (
    .clk(d2w_clk),
    .reset(d2w_reset),
    .io_in(d2w_io_in),
    .io_roundingMode(d2w_io_roundingMode),
    .io_signedOut(d2w_io_signedOut),
    .io_out(d2w_io_out),
    .io_intExceptionFlags(d2w_io_intExceptionFlags)
  );
  assign io_as_double_cmd = in_cmd;
  assign io_as_double_ldst = in_ldst;
  assign io_as_double_wen = in_wen;
  assign io_as_double_ren1 = in_ren1;
  assign io_as_double_ren2 = in_ren2;
  assign io_as_double_ren3 = in_ren3;
  assign io_as_double_swap12 = in_swap12;
  assign io_as_double_swap23 = in_swap23;
  assign io_as_double_single = in_single;
  assign io_as_double_fromint = in_fromint;
  assign io_as_double_toint = in_toint;
  assign io_as_double_fastpipe = in_fastpipe;
  assign io_as_double_fma = in_fma;
  assign io_as_double_div = in_div;
  assign io_as_double_sqrt = in_sqrt;
  assign io_as_double_round = in_round;
  assign io_as_double_wflags = in_wflags;
  assign io_as_double_rm = in_rm;
  assign io_as_double_typ = in_typ;
  assign io_as_double_in1 = in_in1;
  assign io_as_double_in2 = in_in2;
  assign io_as_double_in3 = in_in3;
  assign io_out_valid = valid;
  assign io_out_bits_lt = dcmp_io_lt;
  assign io_out_bits_store = unrec_out;
  assign io_out_bits_toint = GEN_26;
  assign io_out_bits_exc = GEN_27;
  assign RecFNToRecFN_227_clk = clk;
  assign RecFNToRecFN_227_reset = reset;
  assign RecFNToRecFN_227_io_in = io_in_bits_in1[32:0];
  assign RecFNToRecFN_227_io_roundingMode = {{1'd0}, 1'h0};
  assign RecFNToRecFN_94_229_clk = clk;
  assign RecFNToRecFN_94_229_reset = reset;
  assign RecFNToRecFN_94_229_io_in = io_in_bits_in2[32:0];
  assign RecFNToRecFN_94_229_io_roundingMode = {{1'd0}, 1'h0};
  assign T_232 = io_in_bits_ldst == 1'h0;
  assign T_233 = io_in_bits_single & T_232;
  assign GEN_28 = {{1'd0}, 4'hc};
  assign T_236 = io_in_bits_cmd & GEN_28;
  assign T_237 = GEN_28 == T_236;
  assign T_239 = T_237 == 1'h0;
  assign T_240 = T_233 & T_239;
  assign GEN_0 = T_240 ? RecFNToRecFN_227_io_out : io_in_bits_in1;
  assign GEN_1 = T_240 ? RecFNToRecFN_94_229_io_out : io_in_bits_in2;
  assign GEN_2 = io_in_valid ? io_in_bits_cmd : in_cmd;
  assign GEN_3 = io_in_valid ? io_in_bits_ldst : in_ldst;
  assign GEN_4 = io_in_valid ? io_in_bits_wen : in_wen;
  assign GEN_5 = io_in_valid ? io_in_bits_ren1 : in_ren1;
  assign GEN_6 = io_in_valid ? io_in_bits_ren2 : in_ren2;
  assign GEN_7 = io_in_valid ? io_in_bits_ren3 : in_ren3;
  assign GEN_8 = io_in_valid ? io_in_bits_swap12 : in_swap12;
  assign GEN_9 = io_in_valid ? io_in_bits_swap23 : in_swap23;
  assign GEN_10 = io_in_valid ? io_in_bits_single : in_single;
  assign GEN_11 = io_in_valid ? io_in_bits_fromint : in_fromint;
  assign GEN_12 = io_in_valid ? io_in_bits_toint : in_toint;
  assign GEN_13 = io_in_valid ? io_in_bits_fastpipe : in_fastpipe;
  assign GEN_14 = io_in_valid ? io_in_bits_fma : in_fma;
  assign GEN_15 = io_in_valid ? io_in_bits_div : in_div;
  assign GEN_16 = io_in_valid ? io_in_bits_sqrt : in_sqrt;
  assign GEN_17 = io_in_valid ? io_in_bits_round : in_round;
  assign GEN_18 = io_in_valid ? io_in_bits_wflags : in_wflags;
  assign GEN_19 = io_in_valid ? io_in_bits_rm : in_rm;
  assign GEN_20 = io_in_valid ? io_in_bits_typ : in_typ;
  assign GEN_21 = io_in_valid ? GEN_0 : in_in1;
  assign GEN_22 = io_in_valid ? GEN_1 : in_in2;
  assign GEN_23 = io_in_valid ? io_in_bits_in3 : in_in3;
  assign T_241 = in_in1[32];
  assign T_242 = in_in1[31:23];
  assign T_243 = in_in1[22:0];
  assign T_244 = T_242[6:0];
  assign GEN_30 = {{5'd0}, 2'h2};
  assign T_246 = T_244 < GEN_30;
  assign T_247 = T_242[8:6];
  assign GEN_31 = {{2'd0}, 1'h1};
  assign T_249 = T_247 == GEN_31;
  assign T_250 = T_242[8:7];
  assign GEN_32 = {{1'd0}, 1'h1};
  assign T_252 = T_250 == GEN_32;
  assign T_253 = T_252 & T_246;
  assign T_254 = T_249 | T_253;
  assign T_259 = T_246 == 1'h0;
  assign T_260 = T_252 & T_259;
  assign T_263 = T_250 == 2'h2;
  assign T_264 = T_260 | T_263;
  assign T_267 = T_250 == 2'h3;
  assign T_268 = T_242[6];
  assign T_269 = T_267 & T_268;
  assign T_271 = T_242[4:0];
  assign GEN_34 = {{3'd0}, 2'h2};
  assign T_272 = GEN_34 - T_271;
  assign T_273 = T_272[4:0];
  assign T_275 = {1'h1,T_243};
  assign T_276 = T_275 >> T_273;
  assign T_277 = T_276[22:0];
  assign T_278 = T_242[7:0];
  assign T_280 = T_278 - 8'h81;
  assign T_281 = T_280[7:0];
  assign GEN_35 = {{7'd0}, T_267};
  assign T_283 = 8'h0 - GEN_35;
  assign T_284 = T_283[7:0];
  assign T_285 = T_264 ? T_281 : T_284;
  assign T_286 = T_264 | T_269;
  assign T_288 = T_254 ? T_277 : {{22'd0}, 1'h0};
  assign T_289 = T_286 ? T_243 : T_288;
  assign T_290 = {T_241,T_285};
  assign unrec_s = {T_290,T_289};
  assign T_291 = in_in1[64];
  assign T_292 = in_in1[63:52];
  assign T_293 = in_in1[51:0];
  assign T_294 = T_292[9:0];
  assign GEN_36 = {{8'd0}, 2'h2};
  assign T_296 = T_294 < GEN_36;
  assign T_297 = T_292[11:9];
  assign T_299 = T_297 == GEN_31;
  assign T_300 = T_292[11:10];
  assign T_302 = T_300 == GEN_32;
  assign T_303 = T_302 & T_296;
  assign T_304 = T_299 | T_303;
  assign T_309 = T_296 == 1'h0;
  assign T_310 = T_302 & T_309;
  assign T_313 = T_300 == 2'h2;
  assign T_314 = T_310 | T_313;
  assign T_317 = T_300 == 2'h3;
  assign T_318 = T_292[9];
  assign T_319 = T_317 & T_318;
  assign T_321 = T_292[5:0];
  assign GEN_40 = {{4'd0}, 2'h2};
  assign T_322 = GEN_40 - T_321;
  assign T_323 = T_322[5:0];
  assign T_325 = {1'h1,T_293};
  assign T_326 = T_325 >> T_323;
  assign T_327 = T_326[51:0];
  assign T_328 = T_292[10:0];
  assign T_330 = T_328 - 11'h401;
  assign T_331 = T_330[10:0];
  assign GEN_41 = {{10'd0}, T_317};
  assign T_333 = 11'h0 - GEN_41;
  assign T_334 = T_333[10:0];
  assign T_335 = T_314 ? T_331 : T_334;
  assign T_336 = T_314 | T_319;
  assign T_338 = T_304 ? T_327 : {{51'd0}, 1'h0};
  assign T_339 = T_336 ? T_293 : T_338;
  assign T_340 = {T_291,T_335};
  assign unrec_d = {T_340,T_339};
  assign T_341 = unrec_s[31];
  assign GEN_42 = {{31'd0}, T_341};
  assign T_343 = 32'h0 - GEN_42;
  assign T_344 = T_343[31:0];
  assign T_345 = {T_344,unrec_s};
  assign unrec_out = in_single ? T_345 : unrec_d;
  assign T_350 = T_247[2:1];
  assign T_352 = T_350 == 2'h3;
  assign T_359 = T_350 == GEN_32;
  assign T_360 = T_359 & T_246;
  assign T_361 = T_249 | T_360;
  assign T_366 = T_359 & T_259;
  assign T_368 = T_350 == 2'h2;
  assign T_369 = T_366 | T_368;
  assign GEN_47 = {{2'd0}, 1'h0};
  assign T_371 = T_247 == GEN_47;
  assign T_374 = T_268 == 1'h0;
  assign T_375 = T_352 & T_374;
  assign T_376 = ~ T_247;
  assign T_378 = T_376 == GEN_47;
  assign T_379 = T_243[22];
  assign T_381 = T_379 == 1'h0;
  assign T_382 = T_378 & T_381;
  assign T_384 = T_378 & T_379;
  assign T_386 = T_241 == 1'h0;
  assign T_387 = T_375 & T_386;
  assign T_390 = T_369 & T_386;
  assign T_393 = T_361 & T_386;
  assign T_396 = T_371 & T_386;
  assign T_397 = T_371 & T_241;
  assign T_398 = T_361 & T_241;
  assign T_399 = T_369 & T_241;
  assign T_400 = T_375 & T_241;
  assign T_401 = {T_399,T_400};
  assign T_402 = {T_396,T_397};
  assign T_403 = {T_402,T_398};
  assign T_404 = {T_403,T_401};
  assign T_405 = {T_390,T_393};
  assign T_406 = {T_384,T_382};
  assign T_407 = {T_406,T_387};
  assign T_408 = {T_407,T_405};
  assign classify_s = {T_408,T_404};
  assign T_413 = T_297[2:1];
  assign T_415 = T_413 == 2'h3;
  assign T_422 = T_413 == GEN_32;
  assign T_423 = T_422 & T_296;
  assign T_424 = T_299 | T_423;
  assign T_429 = T_422 & T_309;
  assign T_431 = T_413 == 2'h2;
  assign T_432 = T_429 | T_431;
  assign T_434 = T_297 == GEN_47;
  assign T_437 = T_318 == 1'h0;
  assign T_438 = T_415 & T_437;
  assign T_439 = ~ T_297;
  assign T_441 = T_439 == GEN_47;
  assign T_442 = T_293[51];
  assign T_444 = T_442 == 1'h0;
  assign T_445 = T_441 & T_444;
  assign T_447 = T_441 & T_442;
  assign T_449 = T_291 == 1'h0;
  assign T_450 = T_438 & T_449;
  assign T_453 = T_432 & T_449;
  assign T_456 = T_424 & T_449;
  assign T_459 = T_434 & T_449;
  assign T_460 = T_434 & T_291;
  assign T_461 = T_424 & T_291;
  assign T_462 = T_432 & T_291;
  assign T_463 = T_438 & T_291;
  assign T_464 = {T_462,T_463};
  assign T_465 = {T_459,T_460};
  assign T_466 = {T_465,T_461};
  assign T_467 = {T_466,T_464};
  assign T_468 = {T_453,T_456};
  assign T_469 = {T_447,T_445};
  assign T_470 = {T_469,T_450};
  assign T_471 = {T_470,T_468};
  assign classify_d = {T_471,T_467};
  assign classify_out = in_single ? classify_s : classify_d;
  assign dcmp_clk = clk;
  assign dcmp_reset = reset;
  assign dcmp_io_a = in_in1;
  assign dcmp_io_b = in_in2;
  assign dcmp_io_signaling = 1'h1;
  assign T_473 = ~ in_rm;
  assign T_474 = {dcmp_io_lt,dcmp_io_eq};
  assign GEN_55 = {{1'd0}, T_474};
  assign T_475 = T_473 & GEN_55;
  assign dcmp_out = T_475 != GEN_47;
  assign d2l_clk = clk;
  assign d2l_reset = reset;
  assign d2l_io_in = in_in1;
  assign d2l_io_roundingMode = in_rm[1:0];
  assign d2l_io_signedOut = T_478;
  assign d2w_clk = clk;
  assign d2w_reset = reset;
  assign d2w_io_in = in_in1;
  assign d2w_io_roundingMode = in_rm[1:0];
  assign d2w_io_signedOut = T_478;
  assign T_477 = in_typ[0];
  assign T_478 = ~ T_477;
  assign T_481 = in_rm[0];
  assign T_482 = T_481 ? {{54'd0}, classify_out} : unrec_out;
  assign T_486 = in_cmd & GEN_28;
  assign GEN_58 = {{2'd0}, 3'h4};
  assign T_487 = GEN_58 == T_486;
  assign GEN_24 = T_487 ? {{63'd0}, dcmp_out} : T_482;
  assign GEN_25 = T_487 ? dcmp_io_exceptionFlags : {{4'd0}, 1'h0};
  assign GEN_60 = {{1'd0}, 4'h8};
  assign T_491 = GEN_60 == T_486;
  assign T_492 = in_typ[1];
  assign T_493 = $signed(d2l_io_out);
  assign T_494 = $signed(d2w_io_out);
  assign T_495 = T_492 ? $signed(T_493) : $signed({{32{T_494[31]}},T_494});
  assign T_496 = $unsigned(T_495);
  assign T_498 = T_492 ? d2l_io_intExceptionFlags : d2w_io_intExceptionFlags;
  assign T_499 = T_498[2:1];
  assign GEN_61 = {{1'd0}, 1'h0};
  assign T_501 = T_499 != GEN_61;
  assign T_503 = T_498[0];
  assign T_504 = {T_501,3'h0};
  assign T_505 = {T_504,T_503};
  assign GEN_26 = T_491 ? T_496 : GEN_24;
  assign GEN_27 = T_491 ? T_505 : GEN_25;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_29 = {1{$random}};
  in_cmd = GEN_29[4:0];
  GEN_33 = {1{$random}};
  in_ldst = GEN_33[0:0];
  GEN_37 = {1{$random}};
  in_wen = GEN_37[0:0];
  GEN_38 = {1{$random}};
  in_ren1 = GEN_38[0:0];
  GEN_39 = {1{$random}};
  in_ren2 = GEN_39[0:0];
  GEN_43 = {1{$random}};
  in_ren3 = GEN_43[0:0];
  GEN_44 = {1{$random}};
  in_swap12 = GEN_44[0:0];
  GEN_45 = {1{$random}};
  in_swap23 = GEN_45[0:0];
  GEN_46 = {1{$random}};
  in_single = GEN_46[0:0];
  GEN_48 = {1{$random}};
  in_fromint = GEN_48[0:0];
  GEN_49 = {1{$random}};
  in_toint = GEN_49[0:0];
  GEN_50 = {1{$random}};
  in_fastpipe = GEN_50[0:0];
  GEN_51 = {1{$random}};
  in_fma = GEN_51[0:0];
  GEN_52 = {1{$random}};
  in_div = GEN_52[0:0];
  GEN_53 = {1{$random}};
  in_sqrt = GEN_53[0:0];
  GEN_54 = {1{$random}};
  in_round = GEN_54[0:0];
  GEN_56 = {1{$random}};
  in_wflags = GEN_56[0:0];
  GEN_57 = {1{$random}};
  in_rm = GEN_57[2:0];
  GEN_59 = {1{$random}};
  in_typ = GEN_59[1:0];
  GEN_62 = {3{$random}};
  in_in1 = GEN_62[64:0];
  GEN_63 = {3{$random}};
  in_in2 = GEN_63[64:0];
  GEN_64 = {3{$random}};
  in_in3 = GEN_64[64:0];
  GEN_65 = {1{$random}};
  valid = GEN_65[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      in_cmd <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      in_ldst <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      in_wen <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      in_ren1 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      in_ren2 <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      in_ren3 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      in_swap12 <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      in_swap23 <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      in_single <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      in_fromint <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      in_toint <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      in_fastpipe <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      in_fma <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      in_div <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      in_sqrt <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      in_round <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      in_wflags <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      in_rm <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      in_typ <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      in_in1 <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      in_in2 <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      in_in3 <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      valid <= io_in_valid;
    end
  end
endmodule
module INToRecFN(
  input   clk,
  input   reset,
  input   io_signedIn,
  input  [63:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  T_5;
  wire  sign;
  wire [63:0] GEN_0;
  wire [64:0] T_7;
  wire [63:0] T_8;
  wire [63:0] absIn;
  wire  T_10;
  wire  T_12;
  wire  T_14;
  wire  T_16;
  wire  T_18;
  wire  T_20;
  wire  T_22;
  wire  T_24;
  wire  T_26;
  wire  T_28;
  wire  T_30;
  wire  T_32;
  wire  T_34;
  wire  T_36;
  wire  T_38;
  wire  T_40;
  wire  T_42;
  wire  T_44;
  wire  T_46;
  wire  T_48;
  wire  T_50;
  wire  T_52;
  wire  T_54;
  wire  T_56;
  wire  T_58;
  wire  T_60;
  wire  T_62;
  wire  T_64;
  wire  T_66;
  wire  T_68;
  wire  T_70;
  wire  T_72;
  wire  T_74;
  wire  T_76;
  wire  T_78;
  wire  T_80;
  wire  T_82;
  wire  T_84;
  wire  T_86;
  wire  T_88;
  wire  T_90;
  wire  T_92;
  wire  T_94;
  wire  T_96;
  wire  T_98;
  wire  T_100;
  wire  T_102;
  wire  T_104;
  wire  T_106;
  wire  T_108;
  wire  T_110;
  wire  T_112;
  wire  T_114;
  wire  T_116;
  wire  T_118;
  wire  T_120;
  wire  T_122;
  wire  T_124;
  wire  T_126;
  wire  T_128;
  wire  T_130;
  wire  T_132;
  wire  T_134;
  wire [1:0] T_136;
  wire [1:0] T_137;
  wire [2:0] T_138;
  wire [2:0] T_139;
  wire [2:0] T_140;
  wire [2:0] T_141;
  wire [3:0] T_142;
  wire [3:0] T_143;
  wire [3:0] T_144;
  wire [3:0] T_145;
  wire [3:0] T_146;
  wire [3:0] T_147;
  wire [3:0] T_148;
  wire [3:0] T_149;
  wire [4:0] T_150;
  wire [4:0] T_151;
  wire [4:0] T_152;
  wire [4:0] T_153;
  wire [4:0] T_154;
  wire [4:0] T_155;
  wire [4:0] T_156;
  wire [4:0] T_157;
  wire [4:0] T_158;
  wire [4:0] T_159;
  wire [4:0] T_160;
  wire [4:0] T_161;
  wire [4:0] T_162;
  wire [4:0] T_163;
  wire [4:0] T_164;
  wire [4:0] T_165;
  wire [5:0] T_166;
  wire [5:0] T_167;
  wire [5:0] T_168;
  wire [5:0] T_169;
  wire [5:0] T_170;
  wire [5:0] T_171;
  wire [5:0] T_172;
  wire [5:0] T_173;
  wire [5:0] T_174;
  wire [5:0] T_175;
  wire [5:0] T_176;
  wire [5:0] T_177;
  wire [5:0] T_178;
  wire [5:0] T_179;
  wire [5:0] T_180;
  wire [5:0] T_181;
  wire [5:0] T_182;
  wire [5:0] T_183;
  wire [5:0] T_184;
  wire [5:0] T_185;
  wire [5:0] T_186;
  wire [5:0] T_187;
  wire [5:0] T_188;
  wire [5:0] T_189;
  wire [5:0] T_190;
  wire [5:0] T_191;
  wire [5:0] T_192;
  wire [5:0] T_193;
  wire [5:0] T_194;
  wire [5:0] T_195;
  wire [5:0] T_196;
  wire [5:0] T_197;
  wire [5:0] normCount;
  wire [126:0] GEN_1;
  wire [126:0] T_198;
  wire [63:0] normAbsIn;
  wire [1:0] T_200;
  wire [38:0] T_201;
  wire [38:0] GEN_2;
  wire  T_203;
  wire [2:0] roundBits;
  wire [1:0] T_204;
  wire [1:0] GEN_3;
  wire  roundInexact;
  wire  T_206;
  wire [1:0] T_207;
  wire [1:0] T_208;
  wire  T_210;
  wire [1:0] T_212;
  wire  T_214;
  wire  T_215;
  wire  T_217;
  wire  T_218;
  wire  T_219;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire  T_225;
  wire  T_226;
  wire  T_228;
  wire  round;
  wire [23:0] T_230;
  wire [24:0] unroundedNorm;
  wire [24:0] GEN_6;
  wire [25:0] T_233;
  wire [24:0] T_234;
  wire [24:0] roundedNorm;
  wire [5:0] T_235;
  wire [6:0] unroundedExp;
  wire [7:0] T_238;
  wire  T_239;
  wire [7:0] GEN_7;
  wire [8:0] T_240;
  wire [7:0] roundedExp;
  wire  T_241;
  wire [8:0] expOut;
  wire [22:0] T_245;
  wire [9:0] T_246;
  wire [32:0] T_247;
  wire [1:0] T_250;
  wire [4:0] T_252;
  assign io_out = T_247;
  assign io_exceptionFlags = T_252;
  assign T_5 = io_in[63];
  assign sign = io_signedIn & T_5;
  assign GEN_0 = {{63'd0}, 1'h0};
  assign T_7 = GEN_0 - io_in;
  assign T_8 = T_7[63:0];
  assign absIn = sign ? T_8 : io_in;
  assign T_10 = absIn[63];
  assign T_12 = absIn[62];
  assign T_14 = absIn[61];
  assign T_16 = absIn[60];
  assign T_18 = absIn[59];
  assign T_20 = absIn[58];
  assign T_22 = absIn[57];
  assign T_24 = absIn[56];
  assign T_26 = absIn[55];
  assign T_28 = absIn[54];
  assign T_30 = absIn[53];
  assign T_32 = absIn[52];
  assign T_34 = absIn[51];
  assign T_36 = absIn[50];
  assign T_38 = absIn[49];
  assign T_40 = absIn[48];
  assign T_42 = absIn[47];
  assign T_44 = absIn[46];
  assign T_46 = absIn[45];
  assign T_48 = absIn[44];
  assign T_50 = absIn[43];
  assign T_52 = absIn[42];
  assign T_54 = absIn[41];
  assign T_56 = absIn[40];
  assign T_58 = absIn[39];
  assign T_60 = absIn[38];
  assign T_62 = absIn[37];
  assign T_64 = absIn[36];
  assign T_66 = absIn[35];
  assign T_68 = absIn[34];
  assign T_70 = absIn[33];
  assign T_72 = absIn[32];
  assign T_74 = absIn[31];
  assign T_76 = absIn[30];
  assign T_78 = absIn[29];
  assign T_80 = absIn[28];
  assign T_82 = absIn[27];
  assign T_84 = absIn[26];
  assign T_86 = absIn[25];
  assign T_88 = absIn[24];
  assign T_90 = absIn[23];
  assign T_92 = absIn[22];
  assign T_94 = absIn[21];
  assign T_96 = absIn[20];
  assign T_98 = absIn[19];
  assign T_100 = absIn[18];
  assign T_102 = absIn[17];
  assign T_104 = absIn[16];
  assign T_106 = absIn[15];
  assign T_108 = absIn[14];
  assign T_110 = absIn[13];
  assign T_112 = absIn[12];
  assign T_114 = absIn[11];
  assign T_116 = absIn[10];
  assign T_118 = absIn[9];
  assign T_120 = absIn[8];
  assign T_122 = absIn[7];
  assign T_124 = absIn[6];
  assign T_126 = absIn[5];
  assign T_128 = absIn[4];
  assign T_130 = absIn[3];
  assign T_132 = absIn[2];
  assign T_134 = absIn[1];
  assign T_136 = T_132 ? 2'h2 : {{1'd0}, T_134};
  assign T_137 = T_130 ? 2'h3 : T_136;
  assign T_138 = T_128 ? 3'h4 : {{1'd0}, T_137};
  assign T_139 = T_126 ? 3'h5 : T_138;
  assign T_140 = T_124 ? 3'h6 : T_139;
  assign T_141 = T_122 ? 3'h7 : T_140;
  assign T_142 = T_120 ? 4'h8 : {{1'd0}, T_141};
  assign T_143 = T_118 ? 4'h9 : T_142;
  assign T_144 = T_116 ? 4'ha : T_143;
  assign T_145 = T_114 ? 4'hb : T_144;
  assign T_146 = T_112 ? 4'hc : T_145;
  assign T_147 = T_110 ? 4'hd : T_146;
  assign T_148 = T_108 ? 4'he : T_147;
  assign T_149 = T_106 ? 4'hf : T_148;
  assign T_150 = T_104 ? 5'h10 : {{1'd0}, T_149};
  assign T_151 = T_102 ? 5'h11 : T_150;
  assign T_152 = T_100 ? 5'h12 : T_151;
  assign T_153 = T_98 ? 5'h13 : T_152;
  assign T_154 = T_96 ? 5'h14 : T_153;
  assign T_155 = T_94 ? 5'h15 : T_154;
  assign T_156 = T_92 ? 5'h16 : T_155;
  assign T_157 = T_90 ? 5'h17 : T_156;
  assign T_158 = T_88 ? 5'h18 : T_157;
  assign T_159 = T_86 ? 5'h19 : T_158;
  assign T_160 = T_84 ? 5'h1a : T_159;
  assign T_161 = T_82 ? 5'h1b : T_160;
  assign T_162 = T_80 ? 5'h1c : T_161;
  assign T_163 = T_78 ? 5'h1d : T_162;
  assign T_164 = T_76 ? 5'h1e : T_163;
  assign T_165 = T_74 ? 5'h1f : T_164;
  assign T_166 = T_72 ? 6'h20 : {{1'd0}, T_165};
  assign T_167 = T_70 ? 6'h21 : T_166;
  assign T_168 = T_68 ? 6'h22 : T_167;
  assign T_169 = T_66 ? 6'h23 : T_168;
  assign T_170 = T_64 ? 6'h24 : T_169;
  assign T_171 = T_62 ? 6'h25 : T_170;
  assign T_172 = T_60 ? 6'h26 : T_171;
  assign T_173 = T_58 ? 6'h27 : T_172;
  assign T_174 = T_56 ? 6'h28 : T_173;
  assign T_175 = T_54 ? 6'h29 : T_174;
  assign T_176 = T_52 ? 6'h2a : T_175;
  assign T_177 = T_50 ? 6'h2b : T_176;
  assign T_178 = T_48 ? 6'h2c : T_177;
  assign T_179 = T_46 ? 6'h2d : T_178;
  assign T_180 = T_44 ? 6'h2e : T_179;
  assign T_181 = T_42 ? 6'h2f : T_180;
  assign T_182 = T_40 ? 6'h30 : T_181;
  assign T_183 = T_38 ? 6'h31 : T_182;
  assign T_184 = T_36 ? 6'h32 : T_183;
  assign T_185 = T_34 ? 6'h33 : T_184;
  assign T_186 = T_32 ? 6'h34 : T_185;
  assign T_187 = T_30 ? 6'h35 : T_186;
  assign T_188 = T_28 ? 6'h36 : T_187;
  assign T_189 = T_26 ? 6'h37 : T_188;
  assign T_190 = T_24 ? 6'h38 : T_189;
  assign T_191 = T_22 ? 6'h39 : T_190;
  assign T_192 = T_20 ? 6'h3a : T_191;
  assign T_193 = T_18 ? 6'h3b : T_192;
  assign T_194 = T_16 ? 6'h3c : T_193;
  assign T_195 = T_14 ? 6'h3d : T_194;
  assign T_196 = T_12 ? 6'h3e : T_195;
  assign T_197 = T_10 ? 6'h3f : T_196;
  assign normCount = ~ T_197;
  assign GEN_1 = {{63'd0}, absIn};
  assign T_198 = GEN_1 << normCount;
  assign normAbsIn = T_198[63:0];
  assign T_200 = normAbsIn[40:39];
  assign T_201 = normAbsIn[38:0];
  assign GEN_2 = {{38'd0}, 1'h0};
  assign T_203 = T_201 != GEN_2;
  assign roundBits = {T_200,T_203};
  assign T_204 = roundBits[1:0];
  assign GEN_3 = {{1'd0}, 1'h0};
  assign roundInexact = T_204 != GEN_3;
  assign T_206 = io_roundingMode == 2'h0;
  assign T_207 = roundBits[2:1];
  assign T_208 = ~ T_207;
  assign T_210 = T_208 == GEN_3;
  assign T_212 = ~ T_204;
  assign T_214 = T_212 == GEN_3;
  assign T_215 = T_210 | T_214;
  assign T_217 = T_206 ? T_215 : 1'h0;
  assign T_218 = io_roundingMode == 2'h2;
  assign T_219 = sign & roundInexact;
  assign T_221 = T_218 ? T_219 : 1'h0;
  assign T_222 = T_217 | T_221;
  assign T_223 = io_roundingMode == 2'h3;
  assign T_225 = sign == 1'h0;
  assign T_226 = T_225 & roundInexact;
  assign T_228 = T_223 ? T_226 : 1'h0;
  assign round = T_222 | T_228;
  assign T_230 = normAbsIn[63:40];
  assign unroundedNorm = {1'h0,T_230};
  assign GEN_6 = {{24'd0}, 1'h1};
  assign T_233 = unroundedNorm + GEN_6;
  assign T_234 = T_233[24:0];
  assign roundedNorm = round ? T_234 : unroundedNorm;
  assign T_235 = ~ normCount;
  assign unroundedExp = {1'h0,T_235};
  assign T_238 = {1'h0,unroundedExp};
  assign T_239 = roundedNorm[24];
  assign GEN_7 = {{7'd0}, T_239};
  assign T_240 = T_238 + GEN_7;
  assign roundedExp = T_240[7:0];
  assign T_241 = normAbsIn[63];
  assign expOut = {T_241,roundedExp};
  assign T_245 = roundedNorm[22:0];
  assign T_246 = {sign,expOut};
  assign T_247 = {T_246,T_245};
  assign T_250 = {1'h0,roundInexact};
  assign T_252 = {3'h0,T_250};
endmodule
module INToRecFN_96(
  input   clk,
  input   reset,
  input   io_signedIn,
  input  [63:0] io_in,
  input  [1:0] io_roundingMode,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  T_5;
  wire  sign;
  wire [63:0] GEN_0;
  wire [64:0] T_7;
  wire [63:0] T_8;
  wire [63:0] absIn;
  wire  T_10;
  wire  T_12;
  wire  T_14;
  wire  T_16;
  wire  T_18;
  wire  T_20;
  wire  T_22;
  wire  T_24;
  wire  T_26;
  wire  T_28;
  wire  T_30;
  wire  T_32;
  wire  T_34;
  wire  T_36;
  wire  T_38;
  wire  T_40;
  wire  T_42;
  wire  T_44;
  wire  T_46;
  wire  T_48;
  wire  T_50;
  wire  T_52;
  wire  T_54;
  wire  T_56;
  wire  T_58;
  wire  T_60;
  wire  T_62;
  wire  T_64;
  wire  T_66;
  wire  T_68;
  wire  T_70;
  wire  T_72;
  wire  T_74;
  wire  T_76;
  wire  T_78;
  wire  T_80;
  wire  T_82;
  wire  T_84;
  wire  T_86;
  wire  T_88;
  wire  T_90;
  wire  T_92;
  wire  T_94;
  wire  T_96;
  wire  T_98;
  wire  T_100;
  wire  T_102;
  wire  T_104;
  wire  T_106;
  wire  T_108;
  wire  T_110;
  wire  T_112;
  wire  T_114;
  wire  T_116;
  wire  T_118;
  wire  T_120;
  wire  T_122;
  wire  T_124;
  wire  T_126;
  wire  T_128;
  wire  T_130;
  wire  T_132;
  wire  T_134;
  wire [1:0] T_136;
  wire [1:0] T_137;
  wire [2:0] T_138;
  wire [2:0] T_139;
  wire [2:0] T_140;
  wire [2:0] T_141;
  wire [3:0] T_142;
  wire [3:0] T_143;
  wire [3:0] T_144;
  wire [3:0] T_145;
  wire [3:0] T_146;
  wire [3:0] T_147;
  wire [3:0] T_148;
  wire [3:0] T_149;
  wire [4:0] T_150;
  wire [4:0] T_151;
  wire [4:0] T_152;
  wire [4:0] T_153;
  wire [4:0] T_154;
  wire [4:0] T_155;
  wire [4:0] T_156;
  wire [4:0] T_157;
  wire [4:0] T_158;
  wire [4:0] T_159;
  wire [4:0] T_160;
  wire [4:0] T_161;
  wire [4:0] T_162;
  wire [4:0] T_163;
  wire [4:0] T_164;
  wire [4:0] T_165;
  wire [5:0] T_166;
  wire [5:0] T_167;
  wire [5:0] T_168;
  wire [5:0] T_169;
  wire [5:0] T_170;
  wire [5:0] T_171;
  wire [5:0] T_172;
  wire [5:0] T_173;
  wire [5:0] T_174;
  wire [5:0] T_175;
  wire [5:0] T_176;
  wire [5:0] T_177;
  wire [5:0] T_178;
  wire [5:0] T_179;
  wire [5:0] T_180;
  wire [5:0] T_181;
  wire [5:0] T_182;
  wire [5:0] T_183;
  wire [5:0] T_184;
  wire [5:0] T_185;
  wire [5:0] T_186;
  wire [5:0] T_187;
  wire [5:0] T_188;
  wire [5:0] T_189;
  wire [5:0] T_190;
  wire [5:0] T_191;
  wire [5:0] T_192;
  wire [5:0] T_193;
  wire [5:0] T_194;
  wire [5:0] T_195;
  wire [5:0] T_196;
  wire [5:0] T_197;
  wire [5:0] normCount;
  wire [126:0] GEN_1;
  wire [126:0] T_198;
  wire [63:0] normAbsIn;
  wire [1:0] T_200;
  wire [9:0] T_201;
  wire [9:0] GEN_2;
  wire  T_203;
  wire [2:0] roundBits;
  wire [1:0] T_204;
  wire [1:0] GEN_3;
  wire  roundInexact;
  wire  T_206;
  wire [1:0] T_207;
  wire [1:0] T_208;
  wire  T_210;
  wire [1:0] T_212;
  wire  T_214;
  wire  T_215;
  wire  T_217;
  wire  T_218;
  wire  T_219;
  wire  T_221;
  wire  T_222;
  wire  T_223;
  wire  T_225;
  wire  T_226;
  wire  T_228;
  wire  round;
  wire [52:0] T_230;
  wire [53:0] unroundedNorm;
  wire [53:0] GEN_6;
  wire [54:0] T_233;
  wire [53:0] T_234;
  wire [53:0] roundedNorm;
  wire [5:0] T_235;
  wire [9:0] unroundedExp;
  wire [10:0] T_238;
  wire  T_239;
  wire [10:0] GEN_7;
  wire [11:0] T_240;
  wire [10:0] roundedExp;
  wire  T_241;
  wire [11:0] expOut;
  wire [51:0] T_245;
  wire [12:0] T_246;
  wire [64:0] T_247;
  wire [1:0] T_250;
  wire [4:0] T_252;
  assign io_out = T_247;
  assign io_exceptionFlags = T_252;
  assign T_5 = io_in[63];
  assign sign = io_signedIn & T_5;
  assign GEN_0 = {{63'd0}, 1'h0};
  assign T_7 = GEN_0 - io_in;
  assign T_8 = T_7[63:0];
  assign absIn = sign ? T_8 : io_in;
  assign T_10 = absIn[63];
  assign T_12 = absIn[62];
  assign T_14 = absIn[61];
  assign T_16 = absIn[60];
  assign T_18 = absIn[59];
  assign T_20 = absIn[58];
  assign T_22 = absIn[57];
  assign T_24 = absIn[56];
  assign T_26 = absIn[55];
  assign T_28 = absIn[54];
  assign T_30 = absIn[53];
  assign T_32 = absIn[52];
  assign T_34 = absIn[51];
  assign T_36 = absIn[50];
  assign T_38 = absIn[49];
  assign T_40 = absIn[48];
  assign T_42 = absIn[47];
  assign T_44 = absIn[46];
  assign T_46 = absIn[45];
  assign T_48 = absIn[44];
  assign T_50 = absIn[43];
  assign T_52 = absIn[42];
  assign T_54 = absIn[41];
  assign T_56 = absIn[40];
  assign T_58 = absIn[39];
  assign T_60 = absIn[38];
  assign T_62 = absIn[37];
  assign T_64 = absIn[36];
  assign T_66 = absIn[35];
  assign T_68 = absIn[34];
  assign T_70 = absIn[33];
  assign T_72 = absIn[32];
  assign T_74 = absIn[31];
  assign T_76 = absIn[30];
  assign T_78 = absIn[29];
  assign T_80 = absIn[28];
  assign T_82 = absIn[27];
  assign T_84 = absIn[26];
  assign T_86 = absIn[25];
  assign T_88 = absIn[24];
  assign T_90 = absIn[23];
  assign T_92 = absIn[22];
  assign T_94 = absIn[21];
  assign T_96 = absIn[20];
  assign T_98 = absIn[19];
  assign T_100 = absIn[18];
  assign T_102 = absIn[17];
  assign T_104 = absIn[16];
  assign T_106 = absIn[15];
  assign T_108 = absIn[14];
  assign T_110 = absIn[13];
  assign T_112 = absIn[12];
  assign T_114 = absIn[11];
  assign T_116 = absIn[10];
  assign T_118 = absIn[9];
  assign T_120 = absIn[8];
  assign T_122 = absIn[7];
  assign T_124 = absIn[6];
  assign T_126 = absIn[5];
  assign T_128 = absIn[4];
  assign T_130 = absIn[3];
  assign T_132 = absIn[2];
  assign T_134 = absIn[1];
  assign T_136 = T_132 ? 2'h2 : {{1'd0}, T_134};
  assign T_137 = T_130 ? 2'h3 : T_136;
  assign T_138 = T_128 ? 3'h4 : {{1'd0}, T_137};
  assign T_139 = T_126 ? 3'h5 : T_138;
  assign T_140 = T_124 ? 3'h6 : T_139;
  assign T_141 = T_122 ? 3'h7 : T_140;
  assign T_142 = T_120 ? 4'h8 : {{1'd0}, T_141};
  assign T_143 = T_118 ? 4'h9 : T_142;
  assign T_144 = T_116 ? 4'ha : T_143;
  assign T_145 = T_114 ? 4'hb : T_144;
  assign T_146 = T_112 ? 4'hc : T_145;
  assign T_147 = T_110 ? 4'hd : T_146;
  assign T_148 = T_108 ? 4'he : T_147;
  assign T_149 = T_106 ? 4'hf : T_148;
  assign T_150 = T_104 ? 5'h10 : {{1'd0}, T_149};
  assign T_151 = T_102 ? 5'h11 : T_150;
  assign T_152 = T_100 ? 5'h12 : T_151;
  assign T_153 = T_98 ? 5'h13 : T_152;
  assign T_154 = T_96 ? 5'h14 : T_153;
  assign T_155 = T_94 ? 5'h15 : T_154;
  assign T_156 = T_92 ? 5'h16 : T_155;
  assign T_157 = T_90 ? 5'h17 : T_156;
  assign T_158 = T_88 ? 5'h18 : T_157;
  assign T_159 = T_86 ? 5'h19 : T_158;
  assign T_160 = T_84 ? 5'h1a : T_159;
  assign T_161 = T_82 ? 5'h1b : T_160;
  assign T_162 = T_80 ? 5'h1c : T_161;
  assign T_163 = T_78 ? 5'h1d : T_162;
  assign T_164 = T_76 ? 5'h1e : T_163;
  assign T_165 = T_74 ? 5'h1f : T_164;
  assign T_166 = T_72 ? 6'h20 : {{1'd0}, T_165};
  assign T_167 = T_70 ? 6'h21 : T_166;
  assign T_168 = T_68 ? 6'h22 : T_167;
  assign T_169 = T_66 ? 6'h23 : T_168;
  assign T_170 = T_64 ? 6'h24 : T_169;
  assign T_171 = T_62 ? 6'h25 : T_170;
  assign T_172 = T_60 ? 6'h26 : T_171;
  assign T_173 = T_58 ? 6'h27 : T_172;
  assign T_174 = T_56 ? 6'h28 : T_173;
  assign T_175 = T_54 ? 6'h29 : T_174;
  assign T_176 = T_52 ? 6'h2a : T_175;
  assign T_177 = T_50 ? 6'h2b : T_176;
  assign T_178 = T_48 ? 6'h2c : T_177;
  assign T_179 = T_46 ? 6'h2d : T_178;
  assign T_180 = T_44 ? 6'h2e : T_179;
  assign T_181 = T_42 ? 6'h2f : T_180;
  assign T_182 = T_40 ? 6'h30 : T_181;
  assign T_183 = T_38 ? 6'h31 : T_182;
  assign T_184 = T_36 ? 6'h32 : T_183;
  assign T_185 = T_34 ? 6'h33 : T_184;
  assign T_186 = T_32 ? 6'h34 : T_185;
  assign T_187 = T_30 ? 6'h35 : T_186;
  assign T_188 = T_28 ? 6'h36 : T_187;
  assign T_189 = T_26 ? 6'h37 : T_188;
  assign T_190 = T_24 ? 6'h38 : T_189;
  assign T_191 = T_22 ? 6'h39 : T_190;
  assign T_192 = T_20 ? 6'h3a : T_191;
  assign T_193 = T_18 ? 6'h3b : T_192;
  assign T_194 = T_16 ? 6'h3c : T_193;
  assign T_195 = T_14 ? 6'h3d : T_194;
  assign T_196 = T_12 ? 6'h3e : T_195;
  assign T_197 = T_10 ? 6'h3f : T_196;
  assign normCount = ~ T_197;
  assign GEN_1 = {{63'd0}, absIn};
  assign T_198 = GEN_1 << normCount;
  assign normAbsIn = T_198[63:0];
  assign T_200 = normAbsIn[11:10];
  assign T_201 = normAbsIn[9:0];
  assign GEN_2 = {{9'd0}, 1'h0};
  assign T_203 = T_201 != GEN_2;
  assign roundBits = {T_200,T_203};
  assign T_204 = roundBits[1:0];
  assign GEN_3 = {{1'd0}, 1'h0};
  assign roundInexact = T_204 != GEN_3;
  assign T_206 = io_roundingMode == 2'h0;
  assign T_207 = roundBits[2:1];
  assign T_208 = ~ T_207;
  assign T_210 = T_208 == GEN_3;
  assign T_212 = ~ T_204;
  assign T_214 = T_212 == GEN_3;
  assign T_215 = T_210 | T_214;
  assign T_217 = T_206 ? T_215 : 1'h0;
  assign T_218 = io_roundingMode == 2'h2;
  assign T_219 = sign & roundInexact;
  assign T_221 = T_218 ? T_219 : 1'h0;
  assign T_222 = T_217 | T_221;
  assign T_223 = io_roundingMode == 2'h3;
  assign T_225 = sign == 1'h0;
  assign T_226 = T_225 & roundInexact;
  assign T_228 = T_223 ? T_226 : 1'h0;
  assign round = T_222 | T_228;
  assign T_230 = normAbsIn[63:11];
  assign unroundedNorm = {1'h0,T_230};
  assign GEN_6 = {{53'd0}, 1'h1};
  assign T_233 = unroundedNorm + GEN_6;
  assign T_234 = T_233[53:0];
  assign roundedNorm = round ? T_234 : unroundedNorm;
  assign T_235 = ~ normCount;
  assign unroundedExp = {4'h0,T_235};
  assign T_238 = {1'h0,unroundedExp};
  assign T_239 = roundedNorm[53];
  assign GEN_7 = {{10'd0}, T_239};
  assign T_240 = T_238 + GEN_7;
  assign roundedExp = T_240[10:0];
  assign T_241 = normAbsIn[63];
  assign expOut = {T_241,roundedExp};
  assign T_245 = roundedNorm[51:0];
  assign T_246 = {sign,expOut};
  assign T_247 = {T_246,T_245};
  assign T_250 = {1'h0,roundInexact};
  assign T_252 = {3'h0,T_250};
endmodule
module IntToFP(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc
);
  reg  T_132;
  reg [31:0] GEN_60;
  reg [4:0] T_133_cmd;
  reg [31:0] GEN_61;
  reg  T_133_ldst;
  reg [31:0] GEN_62;
  reg  T_133_wen;
  reg [31:0] GEN_63;
  reg  T_133_ren1;
  reg [31:0] GEN_64;
  reg  T_133_ren2;
  reg [31:0] GEN_65;
  reg  T_133_ren3;
  reg [31:0] GEN_66;
  reg  T_133_swap12;
  reg [31:0] GEN_67;
  reg  T_133_swap23;
  reg [31:0] GEN_68;
  reg  T_133_single;
  reg [31:0] GEN_69;
  reg  T_133_fromint;
  reg [31:0] GEN_70;
  reg  T_133_toint;
  reg [31:0] GEN_71;
  reg  T_133_fastpipe;
  reg [31:0] GEN_72;
  reg  T_133_fma;
  reg [31:0] GEN_73;
  reg  T_133_div;
  reg [31:0] GEN_74;
  reg  T_133_sqrt;
  reg [31:0] GEN_75;
  reg  T_133_round;
  reg [31:0] GEN_76;
  reg  T_133_wflags;
  reg [31:0] GEN_77;
  reg [2:0] T_133_rm;
  reg [31:0] GEN_78;
  reg [1:0] T_133_typ;
  reg [31:0] GEN_79;
  reg [64:0] T_133_in1;
  reg [95:0] GEN_80;
  reg [64:0] T_133_in2;
  reg [95:0] GEN_81;
  reg [64:0] T_133_in3;
  reg [95:0] GEN_82;
  wire [4:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire [64:0] GEN_19;
  wire [64:0] GEN_20;
  wire [64:0] GEN_21;
  wire  in_valid;
  wire [4:0] in_bits_cmd;
  wire  in_bits_ldst;
  wire  in_bits_wen;
  wire  in_bits_ren1;
  wire  in_bits_ren2;
  wire  in_bits_ren3;
  wire  in_bits_swap12;
  wire  in_bits_swap23;
  wire  in_bits_single;
  wire  in_bits_fromint;
  wire  in_bits_toint;
  wire  in_bits_fastpipe;
  wire  in_bits_fma;
  wire  in_bits_div;
  wire  in_bits_sqrt;
  wire  in_bits_round;
  wire  in_bits_wflags;
  wire [2:0] in_bits_rm;
  wire [1:0] in_bits_typ;
  wire [64:0] in_bits_in1;
  wire [64:0] in_bits_in2;
  wire [64:0] in_bits_in3;
  wire [64:0] mux_data;
  wire [4:0] mux_exc;
  wire  T_257;
  wire [10:0] T_258;
  wire [51:0] T_259;
  wire [10:0] GEN_33;
  wire  T_261;
  wire [51:0] GEN_34;
  wire  T_263;
  wire  T_264;
  wire [63:0] GEN_35;
  wire [63:0] T_265;
  wire  T_266;
  wire  T_268;
  wire  T_270;
  wire  T_272;
  wire  T_274;
  wire  T_276;
  wire  T_278;
  wire  T_280;
  wire  T_282;
  wire  T_284;
  wire  T_286;
  wire  T_288;
  wire  T_290;
  wire  T_292;
  wire  T_294;
  wire  T_296;
  wire  T_298;
  wire  T_300;
  wire  T_302;
  wire  T_304;
  wire  T_306;
  wire  T_308;
  wire  T_310;
  wire  T_312;
  wire  T_314;
  wire  T_316;
  wire  T_318;
  wire  T_320;
  wire  T_322;
  wire  T_324;
  wire  T_326;
  wire  T_328;
  wire  T_330;
  wire  T_332;
  wire  T_334;
  wire  T_336;
  wire  T_338;
  wire  T_340;
  wire  T_342;
  wire  T_344;
  wire  T_346;
  wire  T_348;
  wire  T_350;
  wire  T_352;
  wire  T_354;
  wire  T_356;
  wire  T_358;
  wire  T_360;
  wire  T_362;
  wire  T_364;
  wire  T_366;
  wire  T_368;
  wire  T_370;
  wire  T_372;
  wire  T_374;
  wire  T_376;
  wire  T_378;
  wire  T_380;
  wire  T_382;
  wire  T_384;
  wire  T_386;
  wire  T_388;
  wire  T_390;
  wire [1:0] T_392;
  wire [1:0] T_393;
  wire [2:0] T_394;
  wire [2:0] T_395;
  wire [2:0] T_396;
  wire [2:0] T_397;
  wire [3:0] T_398;
  wire [3:0] T_399;
  wire [3:0] T_400;
  wire [3:0] T_401;
  wire [3:0] T_402;
  wire [3:0] T_403;
  wire [3:0] T_404;
  wire [3:0] T_405;
  wire [4:0] T_406;
  wire [4:0] T_407;
  wire [4:0] T_408;
  wire [4:0] T_409;
  wire [4:0] T_410;
  wire [4:0] T_411;
  wire [4:0] T_412;
  wire [4:0] T_413;
  wire [4:0] T_414;
  wire [4:0] T_415;
  wire [4:0] T_416;
  wire [4:0] T_417;
  wire [4:0] T_418;
  wire [4:0] T_419;
  wire [4:0] T_420;
  wire [4:0] T_421;
  wire [5:0] T_422;
  wire [5:0] T_423;
  wire [5:0] T_424;
  wire [5:0] T_425;
  wire [5:0] T_426;
  wire [5:0] T_427;
  wire [5:0] T_428;
  wire [5:0] T_429;
  wire [5:0] T_430;
  wire [5:0] T_431;
  wire [5:0] T_432;
  wire [5:0] T_433;
  wire [5:0] T_434;
  wire [5:0] T_435;
  wire [5:0] T_436;
  wire [5:0] T_437;
  wire [5:0] T_438;
  wire [5:0] T_439;
  wire [5:0] T_440;
  wire [5:0] T_441;
  wire [5:0] T_442;
  wire [5:0] T_443;
  wire [5:0] T_444;
  wire [5:0] T_445;
  wire [5:0] T_446;
  wire [5:0] T_447;
  wire [5:0] T_448;
  wire [5:0] T_449;
  wire [5:0] T_450;
  wire [5:0] T_451;
  wire [5:0] T_452;
  wire [5:0] T_453;
  wire [5:0] T_454;
  wire [114:0] GEN_36;
  wire [114:0] T_455;
  wire [50:0] T_456;
  wire [51:0] T_458;
  wire [11:0] GEN_37;
  wire [12:0] T_461;
  wire [11:0] T_462;
  wire [11:0] GEN_38;
  wire [11:0] T_463;
  wire [11:0] T_464;
  wire [1:0] T_468;
  wire [10:0] GEN_39;
  wire [10:0] T_469;
  wire [11:0] GEN_40;
  wire [12:0] T_470;
  wire [11:0] T_471;
  wire [1:0] T_472;
  wire  T_474;
  wire  T_476;
  wire  T_477;
  wire [2:0] GEN_41;
  wire [3:0] T_479;
  wire [2:0] T_480;
  wire [11:0] GEN_42;
  wire [11:0] T_481;
  wire [11:0] T_482;
  wire [11:0] T_483;
  wire [9:0] GEN_43;
  wire [9:0] T_484;
  wire [11:0] GEN_44;
  wire [11:0] T_485;
  wire [51:0] T_486;
  wire [12:0] T_487;
  wire [64:0] T_488;
  wire  T_490;
  wire [7:0] T_491;
  wire [22:0] T_492;
  wire [7:0] GEN_45;
  wire  T_494;
  wire [22:0] GEN_46;
  wire  T_496;
  wire  T_497;
  wire [31:0] GEN_47;
  wire [31:0] T_498;
  wire  T_499;
  wire  T_501;
  wire  T_503;
  wire  T_505;
  wire  T_507;
  wire  T_509;
  wire  T_511;
  wire  T_513;
  wire  T_515;
  wire  T_517;
  wire  T_519;
  wire  T_521;
  wire  T_523;
  wire  T_525;
  wire  T_527;
  wire  T_529;
  wire  T_531;
  wire  T_533;
  wire  T_535;
  wire  T_537;
  wire  T_539;
  wire  T_541;
  wire  T_543;
  wire  T_545;
  wire  T_547;
  wire  T_549;
  wire  T_551;
  wire  T_553;
  wire  T_555;
  wire  T_557;
  wire  T_559;
  wire [1:0] T_561;
  wire [1:0] T_562;
  wire [2:0] T_563;
  wire [2:0] T_564;
  wire [2:0] T_565;
  wire [2:0] T_566;
  wire [3:0] T_567;
  wire [3:0] T_568;
  wire [3:0] T_569;
  wire [3:0] T_570;
  wire [3:0] T_571;
  wire [3:0] T_572;
  wire [3:0] T_573;
  wire [3:0] T_574;
  wire [4:0] T_575;
  wire [4:0] T_576;
  wire [4:0] T_577;
  wire [4:0] T_578;
  wire [4:0] T_579;
  wire [4:0] T_580;
  wire [4:0] T_581;
  wire [4:0] T_582;
  wire [4:0] T_583;
  wire [4:0] T_584;
  wire [4:0] T_585;
  wire [4:0] T_586;
  wire [4:0] T_587;
  wire [4:0] T_588;
  wire [4:0] T_589;
  wire [4:0] T_590;
  wire [4:0] T_591;
  wire [53:0] GEN_48;
  wire [53:0] T_592;
  wire [21:0] T_593;
  wire [22:0] T_595;
  wire [8:0] GEN_49;
  wire [9:0] T_598;
  wire [8:0] T_599;
  wire [8:0] GEN_50;
  wire [8:0] T_600;
  wire [8:0] T_601;
  wire [1:0] T_605;
  wire [7:0] GEN_51;
  wire [7:0] T_606;
  wire [8:0] GEN_52;
  wire [9:0] T_607;
  wire [8:0] T_608;
  wire [1:0] T_609;
  wire  T_611;
  wire  T_613;
  wire  T_614;
  wire [2:0] GEN_53;
  wire [3:0] T_616;
  wire [2:0] T_617;
  wire [8:0] GEN_54;
  wire [8:0] T_618;
  wire [8:0] T_619;
  wire [8:0] T_620;
  wire [6:0] GEN_55;
  wire [6:0] T_621;
  wire [8:0] GEN_56;
  wire [8:0] T_622;
  wire [22:0] T_623;
  wire [9:0] T_624;
  wire [32:0] T_625;
  wire [31:0] GEN_57;
  wire [31:0] T_626;
  wire [64:0] T_627;
  wire [64:0] GEN_22;
  wire  T_628;
  wire [64:0] T_629;
  wire  T_630;
  wire [31:0] T_631;
  wire [32:0] T_632;
  wire [31:0] T_634;
  wire [32:0] T_635;
  wire [64:0] longValue;
  wire  l2s_clk;
  wire  l2s_reset;
  wire  l2s_io_signedIn;
  wire [63:0] l2s_io_in;
  wire [1:0] l2s_io_roundingMode;
  wire [32:0] l2s_io_out;
  wire [4:0] l2s_io_exceptionFlags;
  wire  T_637;
  wire [64:0] T_638;
  wire  l2d_clk;
  wire  l2d_reset;
  wire  l2d_io_signedIn;
  wire [63:0] l2d_io_in;
  wire [1:0] l2d_io_roundingMode;
  wire [64:0] l2d_io_out;
  wire [4:0] l2d_io_exceptionFlags;
  wire [4:0] GEN_58;
  wire [4:0] T_644;
  wire [4:0] GEN_59;
  wire  T_645;
  wire [64:0] T_648;
  wire [64:0] GEN_23;
  wire [4:0] GEN_24;
  wire  T_650;
  wire [64:0] GEN_25;
  wire [4:0] GEN_26;
  wire [64:0] GEN_27;
  wire [4:0] GEN_28;
  reg  T_653;
  reg [31:0] GEN_83;
  reg [64:0] T_654_data;
  reg [95:0] GEN_84;
  reg [4:0] T_654_exc;
  reg [31:0] GEN_85;
  wire [64:0] GEN_29;
  wire [4:0] GEN_30;
  reg  T_659;
  reg [31:0] GEN_86;
  reg [64:0] T_660_data;
  reg [95:0] GEN_87;
  reg [4:0] T_660_exc;
  reg [31:0] GEN_88;
  wire [64:0] GEN_31;
  wire [4:0] GEN_32;
  wire  T_671_valid;
  wire [64:0] T_671_bits_data;
  wire [4:0] T_671_bits_exc;
  INToRecFN l2s (
    .clk(l2s_clk),
    .reset(l2s_reset),
    .io_signedIn(l2s_io_signedIn),
    .io_in(l2s_io_in),
    .io_roundingMode(l2s_io_roundingMode),
    .io_out(l2s_io_out),
    .io_exceptionFlags(l2s_io_exceptionFlags)
  );
  INToRecFN_96 l2d (
    .clk(l2d_clk),
    .reset(l2d_reset),
    .io_signedIn(l2d_io_signedIn),
    .io_in(l2d_io_in),
    .io_roundingMode(l2d_io_roundingMode),
    .io_out(l2d_io_out),
    .io_exceptionFlags(l2d_io_exceptionFlags)
  );
  assign io_out_valid = T_671_valid;
  assign io_out_bits_data = T_671_bits_data;
  assign io_out_bits_exc = T_671_bits_exc;
  assign GEN_0 = io_in_valid ? io_in_bits_cmd : T_133_cmd;
  assign GEN_1 = io_in_valid ? io_in_bits_ldst : T_133_ldst;
  assign GEN_2 = io_in_valid ? io_in_bits_wen : T_133_wen;
  assign GEN_3 = io_in_valid ? io_in_bits_ren1 : T_133_ren1;
  assign GEN_4 = io_in_valid ? io_in_bits_ren2 : T_133_ren2;
  assign GEN_5 = io_in_valid ? io_in_bits_ren3 : T_133_ren3;
  assign GEN_6 = io_in_valid ? io_in_bits_swap12 : T_133_swap12;
  assign GEN_7 = io_in_valid ? io_in_bits_swap23 : T_133_swap23;
  assign GEN_8 = io_in_valid ? io_in_bits_single : T_133_single;
  assign GEN_9 = io_in_valid ? io_in_bits_fromint : T_133_fromint;
  assign GEN_10 = io_in_valid ? io_in_bits_toint : T_133_toint;
  assign GEN_11 = io_in_valid ? io_in_bits_fastpipe : T_133_fastpipe;
  assign GEN_12 = io_in_valid ? io_in_bits_fma : T_133_fma;
  assign GEN_13 = io_in_valid ? io_in_bits_div : T_133_div;
  assign GEN_14 = io_in_valid ? io_in_bits_sqrt : T_133_sqrt;
  assign GEN_15 = io_in_valid ? io_in_bits_round : T_133_round;
  assign GEN_16 = io_in_valid ? io_in_bits_wflags : T_133_wflags;
  assign GEN_17 = io_in_valid ? io_in_bits_rm : T_133_rm;
  assign GEN_18 = io_in_valid ? io_in_bits_typ : T_133_typ;
  assign GEN_19 = io_in_valid ? io_in_bits_in1 : T_133_in1;
  assign GEN_20 = io_in_valid ? io_in_bits_in2 : T_133_in2;
  assign GEN_21 = io_in_valid ? io_in_bits_in3 : T_133_in3;
  assign in_valid = T_132;
  assign in_bits_cmd = T_133_cmd;
  assign in_bits_ldst = T_133_ldst;
  assign in_bits_wen = T_133_wen;
  assign in_bits_ren1 = T_133_ren1;
  assign in_bits_ren2 = T_133_ren2;
  assign in_bits_ren3 = T_133_ren3;
  assign in_bits_swap12 = T_133_swap12;
  assign in_bits_swap23 = T_133_swap23;
  assign in_bits_single = T_133_single;
  assign in_bits_fromint = T_133_fromint;
  assign in_bits_toint = T_133_toint;
  assign in_bits_fastpipe = T_133_fastpipe;
  assign in_bits_fma = T_133_fma;
  assign in_bits_div = T_133_div;
  assign in_bits_sqrt = T_133_sqrt;
  assign in_bits_round = T_133_round;
  assign in_bits_wflags = T_133_wflags;
  assign in_bits_rm = T_133_rm;
  assign in_bits_typ = T_133_typ;
  assign in_bits_in1 = T_133_in1;
  assign in_bits_in2 = T_133_in2;
  assign in_bits_in3 = T_133_in3;
  assign mux_data = GEN_27;
  assign mux_exc = GEN_28;
  assign T_257 = in_bits_in1[63];
  assign T_258 = in_bits_in1[62:52];
  assign T_259 = in_bits_in1[51:0];
  assign GEN_33 = {{10'd0}, 1'h0};
  assign T_261 = T_258 == GEN_33;
  assign GEN_34 = {{51'd0}, 1'h0};
  assign T_263 = T_259 == GEN_34;
  assign T_264 = T_261 & T_263;
  assign GEN_35 = {{12'd0}, T_259};
  assign T_265 = GEN_35 << 12;
  assign T_266 = T_265[63];
  assign T_268 = T_265[62];
  assign T_270 = T_265[61];
  assign T_272 = T_265[60];
  assign T_274 = T_265[59];
  assign T_276 = T_265[58];
  assign T_278 = T_265[57];
  assign T_280 = T_265[56];
  assign T_282 = T_265[55];
  assign T_284 = T_265[54];
  assign T_286 = T_265[53];
  assign T_288 = T_265[52];
  assign T_290 = T_265[51];
  assign T_292 = T_265[50];
  assign T_294 = T_265[49];
  assign T_296 = T_265[48];
  assign T_298 = T_265[47];
  assign T_300 = T_265[46];
  assign T_302 = T_265[45];
  assign T_304 = T_265[44];
  assign T_306 = T_265[43];
  assign T_308 = T_265[42];
  assign T_310 = T_265[41];
  assign T_312 = T_265[40];
  assign T_314 = T_265[39];
  assign T_316 = T_265[38];
  assign T_318 = T_265[37];
  assign T_320 = T_265[36];
  assign T_322 = T_265[35];
  assign T_324 = T_265[34];
  assign T_326 = T_265[33];
  assign T_328 = T_265[32];
  assign T_330 = T_265[31];
  assign T_332 = T_265[30];
  assign T_334 = T_265[29];
  assign T_336 = T_265[28];
  assign T_338 = T_265[27];
  assign T_340 = T_265[26];
  assign T_342 = T_265[25];
  assign T_344 = T_265[24];
  assign T_346 = T_265[23];
  assign T_348 = T_265[22];
  assign T_350 = T_265[21];
  assign T_352 = T_265[20];
  assign T_354 = T_265[19];
  assign T_356 = T_265[18];
  assign T_358 = T_265[17];
  assign T_360 = T_265[16];
  assign T_362 = T_265[15];
  assign T_364 = T_265[14];
  assign T_366 = T_265[13];
  assign T_368 = T_265[12];
  assign T_370 = T_265[11];
  assign T_372 = T_265[10];
  assign T_374 = T_265[9];
  assign T_376 = T_265[8];
  assign T_378 = T_265[7];
  assign T_380 = T_265[6];
  assign T_382 = T_265[5];
  assign T_384 = T_265[4];
  assign T_386 = T_265[3];
  assign T_388 = T_265[2];
  assign T_390 = T_265[1];
  assign T_392 = T_388 ? 2'h2 : {{1'd0}, T_390};
  assign T_393 = T_386 ? 2'h3 : T_392;
  assign T_394 = T_384 ? 3'h4 : {{1'd0}, T_393};
  assign T_395 = T_382 ? 3'h5 : T_394;
  assign T_396 = T_380 ? 3'h6 : T_395;
  assign T_397 = T_378 ? 3'h7 : T_396;
  assign T_398 = T_376 ? 4'h8 : {{1'd0}, T_397};
  assign T_399 = T_374 ? 4'h9 : T_398;
  assign T_400 = T_372 ? 4'ha : T_399;
  assign T_401 = T_370 ? 4'hb : T_400;
  assign T_402 = T_368 ? 4'hc : T_401;
  assign T_403 = T_366 ? 4'hd : T_402;
  assign T_404 = T_364 ? 4'he : T_403;
  assign T_405 = T_362 ? 4'hf : T_404;
  assign T_406 = T_360 ? 5'h10 : {{1'd0}, T_405};
  assign T_407 = T_358 ? 5'h11 : T_406;
  assign T_408 = T_356 ? 5'h12 : T_407;
  assign T_409 = T_354 ? 5'h13 : T_408;
  assign T_410 = T_352 ? 5'h14 : T_409;
  assign T_411 = T_350 ? 5'h15 : T_410;
  assign T_412 = T_348 ? 5'h16 : T_411;
  assign T_413 = T_346 ? 5'h17 : T_412;
  assign T_414 = T_344 ? 5'h18 : T_413;
  assign T_415 = T_342 ? 5'h19 : T_414;
  assign T_416 = T_340 ? 5'h1a : T_415;
  assign T_417 = T_338 ? 5'h1b : T_416;
  assign T_418 = T_336 ? 5'h1c : T_417;
  assign T_419 = T_334 ? 5'h1d : T_418;
  assign T_420 = T_332 ? 5'h1e : T_419;
  assign T_421 = T_330 ? 5'h1f : T_420;
  assign T_422 = T_328 ? 6'h20 : {{1'd0}, T_421};
  assign T_423 = T_326 ? 6'h21 : T_422;
  assign T_424 = T_324 ? 6'h22 : T_423;
  assign T_425 = T_322 ? 6'h23 : T_424;
  assign T_426 = T_320 ? 6'h24 : T_425;
  assign T_427 = T_318 ? 6'h25 : T_426;
  assign T_428 = T_316 ? 6'h26 : T_427;
  assign T_429 = T_314 ? 6'h27 : T_428;
  assign T_430 = T_312 ? 6'h28 : T_429;
  assign T_431 = T_310 ? 6'h29 : T_430;
  assign T_432 = T_308 ? 6'h2a : T_431;
  assign T_433 = T_306 ? 6'h2b : T_432;
  assign T_434 = T_304 ? 6'h2c : T_433;
  assign T_435 = T_302 ? 6'h2d : T_434;
  assign T_436 = T_300 ? 6'h2e : T_435;
  assign T_437 = T_298 ? 6'h2f : T_436;
  assign T_438 = T_296 ? 6'h30 : T_437;
  assign T_439 = T_294 ? 6'h31 : T_438;
  assign T_440 = T_292 ? 6'h32 : T_439;
  assign T_441 = T_290 ? 6'h33 : T_440;
  assign T_442 = T_288 ? 6'h34 : T_441;
  assign T_443 = T_286 ? 6'h35 : T_442;
  assign T_444 = T_284 ? 6'h36 : T_443;
  assign T_445 = T_282 ? 6'h37 : T_444;
  assign T_446 = T_280 ? 6'h38 : T_445;
  assign T_447 = T_278 ? 6'h39 : T_446;
  assign T_448 = T_276 ? 6'h3a : T_447;
  assign T_449 = T_274 ? 6'h3b : T_448;
  assign T_450 = T_272 ? 6'h3c : T_449;
  assign T_451 = T_270 ? 6'h3d : T_450;
  assign T_452 = T_268 ? 6'h3e : T_451;
  assign T_453 = T_266 ? 6'h3f : T_452;
  assign T_454 = ~ T_453;
  assign GEN_36 = {{63'd0}, T_259};
  assign T_455 = GEN_36 << T_454;
  assign T_456 = T_455[50:0];
  assign T_458 = {T_456,1'h0};
  assign GEN_37 = {{11'd0}, 1'h1};
  assign T_461 = 12'h0 - GEN_37;
  assign T_462 = T_461[11:0];
  assign GEN_38 = {{6'd0}, T_454};
  assign T_463 = GEN_38 ^ T_462;
  assign T_464 = T_261 ? T_463 : {{1'd0}, T_258};
  assign T_468 = T_261 ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_39 = {{9'd0}, T_468};
  assign T_469 = 11'h400 | GEN_39;
  assign GEN_40 = {{1'd0}, T_469};
  assign T_470 = T_464 + GEN_40;
  assign T_471 = T_470[11:0];
  assign T_472 = T_471[11:10];
  assign T_474 = T_472 == 2'h3;
  assign T_476 = T_263 == 1'h0;
  assign T_477 = T_474 & T_476;
  assign GEN_41 = {{2'd0}, T_264};
  assign T_479 = 3'h0 - GEN_41;
  assign T_480 = T_479[2:0];
  assign GEN_42 = {{9'd0}, T_480};
  assign T_481 = GEN_42 << 9;
  assign T_482 = ~ T_481;
  assign T_483 = T_471 & T_482;
  assign GEN_43 = {{9'd0}, T_477};
  assign T_484 = GEN_43 << 9;
  assign GEN_44 = {{2'd0}, T_484};
  assign T_485 = T_483 | GEN_44;
  assign T_486 = T_261 ? T_458 : T_259;
  assign T_487 = {T_257,T_485};
  assign T_488 = {T_487,T_486};
  assign T_490 = in_bits_in1[31];
  assign T_491 = in_bits_in1[30:23];
  assign T_492 = in_bits_in1[22:0];
  assign GEN_45 = {{7'd0}, 1'h0};
  assign T_494 = T_491 == GEN_45;
  assign GEN_46 = {{22'd0}, 1'h0};
  assign T_496 = T_492 == GEN_46;
  assign T_497 = T_494 & T_496;
  assign GEN_47 = {{9'd0}, T_492};
  assign T_498 = GEN_47 << 9;
  assign T_499 = T_498[31];
  assign T_501 = T_498[30];
  assign T_503 = T_498[29];
  assign T_505 = T_498[28];
  assign T_507 = T_498[27];
  assign T_509 = T_498[26];
  assign T_511 = T_498[25];
  assign T_513 = T_498[24];
  assign T_515 = T_498[23];
  assign T_517 = T_498[22];
  assign T_519 = T_498[21];
  assign T_521 = T_498[20];
  assign T_523 = T_498[19];
  assign T_525 = T_498[18];
  assign T_527 = T_498[17];
  assign T_529 = T_498[16];
  assign T_531 = T_498[15];
  assign T_533 = T_498[14];
  assign T_535 = T_498[13];
  assign T_537 = T_498[12];
  assign T_539 = T_498[11];
  assign T_541 = T_498[10];
  assign T_543 = T_498[9];
  assign T_545 = T_498[8];
  assign T_547 = T_498[7];
  assign T_549 = T_498[6];
  assign T_551 = T_498[5];
  assign T_553 = T_498[4];
  assign T_555 = T_498[3];
  assign T_557 = T_498[2];
  assign T_559 = T_498[1];
  assign T_561 = T_557 ? 2'h2 : {{1'd0}, T_559};
  assign T_562 = T_555 ? 2'h3 : T_561;
  assign T_563 = T_553 ? 3'h4 : {{1'd0}, T_562};
  assign T_564 = T_551 ? 3'h5 : T_563;
  assign T_565 = T_549 ? 3'h6 : T_564;
  assign T_566 = T_547 ? 3'h7 : T_565;
  assign T_567 = T_545 ? 4'h8 : {{1'd0}, T_566};
  assign T_568 = T_543 ? 4'h9 : T_567;
  assign T_569 = T_541 ? 4'ha : T_568;
  assign T_570 = T_539 ? 4'hb : T_569;
  assign T_571 = T_537 ? 4'hc : T_570;
  assign T_572 = T_535 ? 4'hd : T_571;
  assign T_573 = T_533 ? 4'he : T_572;
  assign T_574 = T_531 ? 4'hf : T_573;
  assign T_575 = T_529 ? 5'h10 : {{1'd0}, T_574};
  assign T_576 = T_527 ? 5'h11 : T_575;
  assign T_577 = T_525 ? 5'h12 : T_576;
  assign T_578 = T_523 ? 5'h13 : T_577;
  assign T_579 = T_521 ? 5'h14 : T_578;
  assign T_580 = T_519 ? 5'h15 : T_579;
  assign T_581 = T_517 ? 5'h16 : T_580;
  assign T_582 = T_515 ? 5'h17 : T_581;
  assign T_583 = T_513 ? 5'h18 : T_582;
  assign T_584 = T_511 ? 5'h19 : T_583;
  assign T_585 = T_509 ? 5'h1a : T_584;
  assign T_586 = T_507 ? 5'h1b : T_585;
  assign T_587 = T_505 ? 5'h1c : T_586;
  assign T_588 = T_503 ? 5'h1d : T_587;
  assign T_589 = T_501 ? 5'h1e : T_588;
  assign T_590 = T_499 ? 5'h1f : T_589;
  assign T_591 = ~ T_590;
  assign GEN_48 = {{31'd0}, T_492};
  assign T_592 = GEN_48 << T_591;
  assign T_593 = T_592[21:0];
  assign T_595 = {T_593,1'h0};
  assign GEN_49 = {{8'd0}, 1'h1};
  assign T_598 = 9'h0 - GEN_49;
  assign T_599 = T_598[8:0];
  assign GEN_50 = {{4'd0}, T_591};
  assign T_600 = GEN_50 ^ T_599;
  assign T_601 = T_494 ? T_600 : {{1'd0}, T_491};
  assign T_605 = T_494 ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_51 = {{6'd0}, T_605};
  assign T_606 = 8'h80 | GEN_51;
  assign GEN_52 = {{1'd0}, T_606};
  assign T_607 = T_601 + GEN_52;
  assign T_608 = T_607[8:0];
  assign T_609 = T_608[8:7];
  assign T_611 = T_609 == 2'h3;
  assign T_613 = T_496 == 1'h0;
  assign T_614 = T_611 & T_613;
  assign GEN_53 = {{2'd0}, T_497};
  assign T_616 = 3'h0 - GEN_53;
  assign T_617 = T_616[2:0];
  assign GEN_54 = {{6'd0}, T_617};
  assign T_618 = GEN_54 << 6;
  assign T_619 = ~ T_618;
  assign T_620 = T_608 & T_619;
  assign GEN_55 = {{6'd0}, T_614};
  assign T_621 = GEN_55 << 6;
  assign GEN_56 = {{2'd0}, T_621};
  assign T_622 = T_620 | GEN_56;
  assign T_623 = T_494 ? T_595 : T_492;
  assign T_624 = {T_490,T_622};
  assign T_625 = {T_624,T_623};
  assign GEN_57 = $signed(32'hffffffff);
  assign T_626 = $unsigned(GEN_57);
  assign T_627 = {T_626,T_625};
  assign GEN_22 = in_bits_single ? T_627 : T_488;
  assign T_628 = in_bits_typ[1];
  assign T_629 = $signed(in_bits_in1);
  assign T_630 = in_bits_typ[0];
  assign T_631 = in_bits_in1[31:0];
  assign T_632 = {1'b0,$signed(T_631)};
  assign T_634 = $signed(T_631);
  assign T_635 = T_630 ? $signed(T_632) : $signed({{1{T_634[31]}},T_634});
  assign longValue = T_628 ? $signed(T_629) : $signed({{32{T_635[32]}},T_635});
  assign l2s_clk = clk;
  assign l2s_reset = reset;
  assign l2s_io_signedIn = T_637;
  assign l2s_io_in = T_638[63:0];
  assign l2s_io_roundingMode = in_bits_rm[1:0];
  assign T_637 = ~ T_630;
  assign T_638 = $unsigned(longValue);
  assign l2d_clk = clk;
  assign l2d_reset = reset;
  assign l2d_io_signedIn = T_637;
  assign l2d_io_in = T_638[63:0];
  assign l2d_io_roundingMode = in_bits_rm[1:0];
  assign GEN_58 = {{2'd0}, 3'h4};
  assign T_644 = in_bits_cmd & GEN_58;
  assign GEN_59 = {{4'd0}, 1'h0};
  assign T_645 = GEN_59 == T_644;
  assign T_648 = {T_626,l2s_io_out};
  assign GEN_23 = in_bits_single ? T_648 : GEN_22;
  assign GEN_24 = in_bits_single ? l2s_io_exceptionFlags : {{4'd0}, 1'h0};
  assign T_650 = in_bits_single == 1'h0;
  assign GEN_25 = T_650 ? l2d_io_out : GEN_23;
  assign GEN_26 = T_650 ? l2d_io_exceptionFlags : GEN_24;
  assign GEN_27 = T_645 ? GEN_25 : GEN_22;
  assign GEN_28 = T_645 ? GEN_26 : {{4'd0}, 1'h0};
  assign GEN_29 = in_valid ? mux_data : T_654_data;
  assign GEN_30 = in_valid ? mux_exc : T_654_exc;
  assign GEN_31 = T_653 ? T_654_data : T_660_data;
  assign GEN_32 = T_653 ? T_654_exc : T_660_exc;
  assign T_671_valid = T_659;
  assign T_671_bits_data = T_660_data;
  assign T_671_bits_exc = T_660_exc;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_60 = {1{$random}};
  T_132 = GEN_60[0:0];
  GEN_61 = {1{$random}};
  T_133_cmd = GEN_61[4:0];
  GEN_62 = {1{$random}};
  T_133_ldst = GEN_62[0:0];
  GEN_63 = {1{$random}};
  T_133_wen = GEN_63[0:0];
  GEN_64 = {1{$random}};
  T_133_ren1 = GEN_64[0:0];
  GEN_65 = {1{$random}};
  T_133_ren2 = GEN_65[0:0];
  GEN_66 = {1{$random}};
  T_133_ren3 = GEN_66[0:0];
  GEN_67 = {1{$random}};
  T_133_swap12 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  T_133_swap23 = GEN_68[0:0];
  GEN_69 = {1{$random}};
  T_133_single = GEN_69[0:0];
  GEN_70 = {1{$random}};
  T_133_fromint = GEN_70[0:0];
  GEN_71 = {1{$random}};
  T_133_toint = GEN_71[0:0];
  GEN_72 = {1{$random}};
  T_133_fastpipe = GEN_72[0:0];
  GEN_73 = {1{$random}};
  T_133_fma = GEN_73[0:0];
  GEN_74 = {1{$random}};
  T_133_div = GEN_74[0:0];
  GEN_75 = {1{$random}};
  T_133_sqrt = GEN_75[0:0];
  GEN_76 = {1{$random}};
  T_133_round = GEN_76[0:0];
  GEN_77 = {1{$random}};
  T_133_wflags = GEN_77[0:0];
  GEN_78 = {1{$random}};
  T_133_rm = GEN_78[2:0];
  GEN_79 = {1{$random}};
  T_133_typ = GEN_79[1:0];
  GEN_80 = {3{$random}};
  T_133_in1 = GEN_80[64:0];
  GEN_81 = {3{$random}};
  T_133_in2 = GEN_81[64:0];
  GEN_82 = {3{$random}};
  T_133_in3 = GEN_82[64:0];
  GEN_83 = {1{$random}};
  T_653 = GEN_83[0:0];
  GEN_84 = {3{$random}};
  T_654_data = GEN_84[64:0];
  GEN_85 = {1{$random}};
  T_654_exc = GEN_85[4:0];
  GEN_86 = {1{$random}};
  T_659 = GEN_86[0:0];
  GEN_87 = {3{$random}};
  T_660_data = GEN_87[64:0];
  GEN_88 = {1{$random}};
  T_660_exc = GEN_88[4:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_132 <= 1'h0;
    end else begin
      T_132 <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      T_133_cmd <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      T_133_ldst <= GEN_1;
    end
    if(1'h0) begin
    end else begin
      T_133_wen <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      T_133_ren1 <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      T_133_ren2 <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      T_133_ren3 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      T_133_swap12 <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      T_133_swap23 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      T_133_single <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      T_133_fromint <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      T_133_toint <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      T_133_fastpipe <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      T_133_fma <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      T_133_div <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      T_133_sqrt <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      T_133_round <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_133_wflags <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      T_133_rm <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      T_133_typ <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      T_133_in1 <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      T_133_in2 <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      T_133_in3 <= GEN_21;
    end
    if(reset) begin
      T_653 <= 1'h0;
    end else begin
      T_653 <= in_valid;
    end
    if(1'h0) begin
    end else begin
      T_654_data <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      T_654_exc <= GEN_30;
    end
    if(reset) begin
      T_659 <= 1'h0;
    end else begin
      T_659 <= T_653;
    end
    if(1'h0) begin
    end else begin
      T_660_data <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      T_660_exc <= GEN_32;
    end
  end
endmodule
module RoundRawFNToRecFN(
  input   clk,
  input   reset,
  input   io_invalidExc,
  input   io_infiniteExc,
  input   io_in_sign,
  input   io_in_isNaN,
  input   io_in_isInf,
  input   io_in_isZero,
  input  [9:0] io_in_sExp,
  input  [26:0] io_in_sig,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  roundingMode_nearest_even;
  wire  roundingMode_min;
  wire  roundingMode_max;
  wire  T_19;
  wire  T_21;
  wire  T_22;
  wire  roundMagUp;
  wire  doShiftSigDown1;
  wire  GEN_0;
  wire [9:0] GEN_1;
  wire  T_24;
  wire [24:0] GEN_2;
  wire [25:0] T_26;
  wire [24:0] T_27;
  wire [8:0] T_28;
  wire [8:0] T_29;
  wire [512:0] GEN_3;
  wire [512:0] T_31;
  wire [24:0] T_32;
  wire [15:0] T_33;
  wire [7:0] T_38;
  wire [15:0] GEN_4;
  wire [15:0] T_39;
  wire [7:0] T_40;
  wire [15:0] GEN_5;
  wire [15:0] T_41;
  wire [15:0] T_43;
  wire [15:0] T_44;
  wire [11:0] T_48;
  wire [15:0] GEN_6;
  wire [15:0] T_49;
  wire [11:0] T_50;
  wire [15:0] GEN_7;
  wire [15:0] T_51;
  wire [15:0] T_53;
  wire [15:0] T_54;
  wire [13:0] T_58;
  wire [15:0] GEN_8;
  wire [15:0] T_59;
  wire [13:0] T_60;
  wire [15:0] GEN_9;
  wire [15:0] T_61;
  wire [15:0] T_63;
  wire [15:0] T_64;
  wire [14:0] T_68;
  wire [15:0] GEN_10;
  wire [15:0] T_69;
  wire [14:0] T_70;
  wire [15:0] GEN_11;
  wire [15:0] T_71;
  wire [15:0] T_73;
  wire [15:0] T_74;
  wire [8:0] T_75;
  wire [7:0] T_76;
  wire [3:0] T_81;
  wire [7:0] GEN_12;
  wire [7:0] T_82;
  wire [3:0] T_83;
  wire [7:0] GEN_13;
  wire [7:0] T_84;
  wire [7:0] T_86;
  wire [7:0] T_87;
  wire [5:0] T_91;
  wire [7:0] GEN_14;
  wire [7:0] T_92;
  wire [5:0] T_93;
  wire [7:0] GEN_15;
  wire [7:0] T_94;
  wire [7:0] T_96;
  wire [7:0] T_97;
  wire [6:0] T_101;
  wire [7:0] GEN_16;
  wire [7:0] T_102;
  wire [6:0] T_103;
  wire [7:0] GEN_17;
  wire [7:0] T_104;
  wire [7:0] T_106;
  wire [7:0] T_107;
  wire  T_108;
  wire [8:0] T_109;
  wire [24:0] T_110;
  wire [24:0] T_111;
  wire [24:0] GEN_18;
  wire [24:0] T_112;
  wire [26:0] roundMask;
  wire [25:0] T_114;
  wire [25:0] T_115;
  wire [26:0] GEN_19;
  wire [26:0] roundPosMask;
  wire [26:0] T_116;
  wire [26:0] GEN_20;
  wire  roundPosBit;
  wire [26:0] GEN_21;
  wire [26:0] T_119;
  wire  anyRoundExtra;
  wire  common_inexact;
  wire  T_121;
  wire  T_122;
  wire  T_123;
  wire [26:0] T_124;
  wire [24:0] T_125;
  wire [24:0] GEN_23;
  wire [25:0] T_127;
  wire [24:0] T_128;
  wire  T_131;
  wire  T_132;
  wire [25:0] T_135;
  wire [25:0] T_136;
  wire [25:0] GEN_24;
  wire [25:0] T_137;
  wire [26:0] T_138;
  wire [26:0] T_139;
  wire [24:0] T_140;
  wire [25:0] roundedSig;
  wire [1:0] T_141;
  wire [2:0] T_142;
  wire [9:0] GEN_25;
  wire [10:0] T_143;
  wire [9:0] T_144;
  wire [9:0] sRoundedExp;
  wire [8:0] common_expOut;
  wire [22:0] T_145;
  wire [22:0] T_146;
  wire [22:0] common_fractOut;
  wire [2:0] T_147;
  wire [2:0] GEN_26;
  wire  common_overflow;
  wire [7:0] GEN_27;
  wire [9:0] GEN_28;
  wire  common_totalUnderflow;
  wire [8:0] T_152;
  wire [9:0] GEN_29;
  wire  T_153;
  wire  common_underflow;
  wire  isNaNOut;
  wire  notNaN_isSpecialInfOut;
  wire  T_155;
  wire  T_157;
  wire  T_158;
  wire  T_160;
  wire  commonCase;
  wire  overflow;
  wire  underflow;
  wire  T_161;
  wire  inexact;
  wire  overflow_roundMagUp;
  wire  T_162;
  wire  pegMinNonzeroMagOut;
  wire  T_163;
  wire  T_165;
  wire  pegMaxFiniteMagOut;
  wire  T_166;
  wire  notNaN_isInfOut;
  wire  signOut;
  wire  T_168;
  wire [8:0] T_171;
  wire [8:0] T_172;
  wire [8:0] T_173;
  wire [8:0] T_177;
  wire [8:0] T_178;
  wire [8:0] T_179;
  wire [8:0] T_182;
  wire [8:0] T_183;
  wire [8:0] T_184;
  wire [8:0] T_187;
  wire [8:0] T_188;
  wire [8:0] T_189;
  wire [8:0] T_192;
  wire [8:0] T_193;
  wire [8:0] T_196;
  wire [8:0] T_197;
  wire [8:0] T_200;
  wire [8:0] T_201;
  wire [8:0] T_204;
  wire [8:0] expOut;
  wire  T_205;
  wire [22:0] T_209;
  wire [22:0] T_210;
  wire [22:0] GEN_30;
  wire [23:0] T_212;
  wire [22:0] T_213;
  wire [22:0] fractOut;
  wire [9:0] T_214;
  wire [32:0] T_215;
  wire [1:0] T_216;
  wire [1:0] T_217;
  wire [2:0] T_218;
  wire [4:0] T_219;
  assign io_out = T_215;
  assign io_exceptionFlags = T_219;
  assign roundingMode_nearest_even = io_roundingMode == 2'h0;
  assign roundingMode_min = io_roundingMode == 2'h2;
  assign roundingMode_max = io_roundingMode == 2'h3;
  assign T_19 = roundingMode_min & io_in_sign;
  assign T_21 = io_in_sign == 1'h0;
  assign T_22 = roundingMode_max & T_21;
  assign roundMagUp = T_19 | T_22;
  assign doShiftSigDown1 = io_in_sig[26];
  assign GEN_0 = $signed(1'h0);
  assign GEN_1 = {10{GEN_0}};
  assign T_24 = $signed(io_in_sExp) < $signed(GEN_1);
  assign GEN_2 = {{24'd0}, T_24};
  assign T_26 = 25'h0 - GEN_2;
  assign T_27 = T_26[24:0];
  assign T_28 = io_in_sExp[8:0];
  assign T_29 = ~ T_28;
  assign GEN_3 = $signed(513'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign T_31 = $signed(GEN_3) >>> T_29;
  assign T_32 = T_31[130:106];
  assign T_33 = T_32[15:0];
  assign T_38 = T_33[15:8];
  assign GEN_4 = {{8'd0}, T_38};
  assign T_39 = GEN_4 & 16'hff;
  assign T_40 = T_33[7:0];
  assign GEN_5 = {{8'd0}, T_40};
  assign T_41 = GEN_5 << 8;
  assign T_43 = T_41 & 16'hff00;
  assign T_44 = T_39 | T_43;
  assign T_48 = T_44[15:4];
  assign GEN_6 = {{4'd0}, T_48};
  assign T_49 = GEN_6 & 16'hf0f;
  assign T_50 = T_44[11:0];
  assign GEN_7 = {{4'd0}, T_50};
  assign T_51 = GEN_7 << 4;
  assign T_53 = T_51 & 16'hf0f0;
  assign T_54 = T_49 | T_53;
  assign T_58 = T_54[15:2];
  assign GEN_8 = {{2'd0}, T_58};
  assign T_59 = GEN_8 & 16'h3333;
  assign T_60 = T_54[13:0];
  assign GEN_9 = {{2'd0}, T_60};
  assign T_61 = GEN_9 << 2;
  assign T_63 = T_61 & 16'hcccc;
  assign T_64 = T_59 | T_63;
  assign T_68 = T_64[15:1];
  assign GEN_10 = {{1'd0}, T_68};
  assign T_69 = GEN_10 & 16'h5555;
  assign T_70 = T_64[14:0];
  assign GEN_11 = {{1'd0}, T_70};
  assign T_71 = GEN_11 << 1;
  assign T_73 = T_71 & 16'haaaa;
  assign T_74 = T_69 | T_73;
  assign T_75 = T_32[24:16];
  assign T_76 = T_75[7:0];
  assign T_81 = T_76[7:4];
  assign GEN_12 = {{4'd0}, T_81};
  assign T_82 = GEN_12 & 8'hf;
  assign T_83 = T_76[3:0];
  assign GEN_13 = {{4'd0}, T_83};
  assign T_84 = GEN_13 << 4;
  assign T_86 = T_84 & 8'hf0;
  assign T_87 = T_82 | T_86;
  assign T_91 = T_87[7:2];
  assign GEN_14 = {{2'd0}, T_91};
  assign T_92 = GEN_14 & 8'h33;
  assign T_93 = T_87[5:0];
  assign GEN_15 = {{2'd0}, T_93};
  assign T_94 = GEN_15 << 2;
  assign T_96 = T_94 & 8'hcc;
  assign T_97 = T_92 | T_96;
  assign T_101 = T_97[7:1];
  assign GEN_16 = {{1'd0}, T_101};
  assign T_102 = GEN_16 & 8'h55;
  assign T_103 = T_97[6:0];
  assign GEN_17 = {{1'd0}, T_103};
  assign T_104 = GEN_17 << 1;
  assign T_106 = T_104 & 8'haa;
  assign T_107 = T_102 | T_106;
  assign T_108 = T_75[8];
  assign T_109 = {T_107,T_108};
  assign T_110 = {T_74,T_109};
  assign T_111 = T_27 | T_110;
  assign GEN_18 = {{24'd0}, doShiftSigDown1};
  assign T_112 = T_111 | GEN_18;
  assign roundMask = {T_112,2'h3};
  assign T_114 = roundMask[26:1];
  assign T_115 = ~ T_114;
  assign GEN_19 = {{1'd0}, T_115};
  assign roundPosMask = GEN_19 & roundMask;
  assign T_116 = io_in_sig & roundPosMask;
  assign GEN_20 = {{26'd0}, 1'h0};
  assign roundPosBit = T_116 != GEN_20;
  assign GEN_21 = {{1'd0}, T_114};
  assign T_119 = io_in_sig & GEN_21;
  assign anyRoundExtra = T_119 != GEN_20;
  assign common_inexact = roundPosBit | anyRoundExtra;
  assign T_121 = roundingMode_nearest_even & roundPosBit;
  assign T_122 = roundMagUp & common_inexact;
  assign T_123 = T_121 | T_122;
  assign T_124 = io_in_sig | roundMask;
  assign T_125 = T_124[26:2];
  assign GEN_23 = {{24'd0}, 1'h1};
  assign T_127 = T_125 + GEN_23;
  assign T_128 = T_127[24:0];
  assign T_131 = anyRoundExtra == 1'h0;
  assign T_132 = T_121 & T_131;
  assign T_135 = T_132 ? T_114 : 26'h0;
  assign T_136 = ~ T_135;
  assign GEN_24 = {{1'd0}, T_128};
  assign T_137 = GEN_24 & T_136;
  assign T_138 = ~ roundMask;
  assign T_139 = io_in_sig & T_138;
  assign T_140 = T_139[26:2];
  assign roundedSig = T_123 ? T_137 : {{1'd0}, T_140};
  assign T_141 = roundedSig[25:24];
  assign T_142 = {1'b0,$signed(T_141)};
  assign GEN_25 = {{7{T_142[2]}},T_142};
  assign T_143 = $signed(io_in_sExp) + $signed(GEN_25);
  assign T_144 = T_143[9:0];
  assign sRoundedExp = $signed(T_144);
  assign common_expOut = sRoundedExp[8:0];
  assign T_145 = roundedSig[23:1];
  assign T_146 = roundedSig[22:0];
  assign common_fractOut = doShiftSigDown1 ? T_145 : T_146;
  assign T_147 = sRoundedExp[9:7];
  assign GEN_26 = $signed(3'h3);
  assign common_overflow = $signed(T_147) >= $signed(GEN_26);
  assign GEN_27 = $signed(8'h6b);
  assign GEN_28 = {{2{GEN_27[7]}},GEN_27};
  assign common_totalUnderflow = $signed(sRoundedExp) < $signed(GEN_28);
  assign T_152 = doShiftSigDown1 ? $signed($signed(9'h81)) : $signed($signed(9'h82));
  assign GEN_29 = {{1{T_152[8]}},T_152};
  assign T_153 = $signed(io_in_sExp) < $signed(GEN_29);
  assign common_underflow = common_inexact & T_153;
  assign isNaNOut = io_invalidExc | io_in_isNaN;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T_155 = isNaNOut == 1'h0;
  assign T_157 = notNaN_isSpecialInfOut == 1'h0;
  assign T_158 = T_155 & T_157;
  assign T_160 = io_in_isZero == 1'h0;
  assign commonCase = T_158 & T_160;
  assign overflow = commonCase & common_overflow;
  assign underflow = commonCase & common_underflow;
  assign T_161 = commonCase & common_inexact;
  assign inexact = overflow | T_161;
  assign overflow_roundMagUp = roundingMode_nearest_even | roundMagUp;
  assign T_162 = commonCase & common_totalUnderflow;
  assign pegMinNonzeroMagOut = T_162 & roundMagUp;
  assign T_163 = commonCase & overflow;
  assign T_165 = overflow_roundMagUp == 1'h0;
  assign pegMaxFiniteMagOut = T_163 & T_165;
  assign T_166 = overflow & overflow_roundMagUp;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T_166;
  assign signOut = isNaNOut ? 1'h0 : io_in_sign;
  assign T_168 = io_in_isZero | common_totalUnderflow;
  assign T_171 = T_168 ? 9'h1c0 : {{8'd0}, 1'h0};
  assign T_172 = ~ T_171;
  assign T_173 = common_expOut & T_172;
  assign T_177 = pegMinNonzeroMagOut ? 9'h194 : {{8'd0}, 1'h0};
  assign T_178 = ~ T_177;
  assign T_179 = T_173 & T_178;
  assign T_182 = pegMaxFiniteMagOut ? 9'h80 : {{8'd0}, 1'h0};
  assign T_183 = ~ T_182;
  assign T_184 = T_179 & T_183;
  assign T_187 = notNaN_isInfOut ? 9'h40 : {{8'd0}, 1'h0};
  assign T_188 = ~ T_187;
  assign T_189 = T_184 & T_188;
  assign T_192 = pegMinNonzeroMagOut ? 9'h6b : {{8'd0}, 1'h0};
  assign T_193 = T_189 | T_192;
  assign T_196 = pegMaxFiniteMagOut ? 9'h17f : {{8'd0}, 1'h0};
  assign T_197 = T_193 | T_196;
  assign T_200 = notNaN_isInfOut ? 9'h180 : {{8'd0}, 1'h0};
  assign T_201 = T_197 | T_200;
  assign T_204 = isNaNOut ? 9'h1c0 : {{8'd0}, 1'h0};
  assign expOut = T_201 | T_204;
  assign T_205 = common_totalUnderflow | isNaNOut;
  assign T_209 = isNaNOut ? 23'h400000 : {{22'd0}, 1'h0};
  assign T_210 = T_205 ? T_209 : common_fractOut;
  assign GEN_30 = {{22'd0}, pegMaxFiniteMagOut};
  assign T_212 = 23'h0 - GEN_30;
  assign T_213 = T_212[22:0];
  assign fractOut = T_210 | T_213;
  assign T_214 = {signOut,expOut};
  assign T_215 = {T_214,fractOut};
  assign T_216 = {underflow,inexact};
  assign T_217 = {io_invalidExc,io_infiniteExc};
  assign T_218 = {T_217,overflow};
  assign T_219 = {T_218,T_216};
endmodule
module RecFNToRecFN_98(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_4;
  wire [1:0] T_5;
  wire  T_7;
  wire  T_15_sign;
  wire  T_15_isNaN;
  wire  T_15_isInf;
  wire  T_15_isZero;
  wire [12:0] T_15_sExp;
  wire [55:0] T_15_sig;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire [2:0] T_29;
  wire [2:0] GEN_0;
  wire  T_31;
  wire [12:0] T_32;
  wire [51:0] T_34;
  wire [53:0] T_36;
  wire [55:0] T_37;
  wire [11:0] GEN_1;
  wire [12:0] GEN_2;
  wire [13:0] T_39;
  wire [12:0] T_40;
  wire [12:0] T_41;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [9:0] outRawFloat_sExp;
  wire [26:0] outRawFloat_sig;
  wire  GEN_3;
  wire [12:0] GEN_4;
  wire  T_56;
  wire [2:0] T_57;
  wire  T_59;
  wire [8:0] T_67;
  wire [8:0] T_68;
  wire [9:0] T_69;
  wire [9:0] T_70;
  wire [25:0] T_71;
  wire [29:0] T_72;
  wire [29:0] GEN_6;
  wire  T_74;
  wire [26:0] T_75;
  wire  T_76;
  wire  T_78;
  wire  invalidExc;
  wire  RoundRawFNToRecFN_79_clk;
  wire  RoundRawFNToRecFN_79_reset;
  wire  RoundRawFNToRecFN_79_io_invalidExc;
  wire  RoundRawFNToRecFN_79_io_infiniteExc;
  wire  RoundRawFNToRecFN_79_io_in_sign;
  wire  RoundRawFNToRecFN_79_io_in_isNaN;
  wire  RoundRawFNToRecFN_79_io_in_isInf;
  wire  RoundRawFNToRecFN_79_io_in_isZero;
  wire [9:0] RoundRawFNToRecFN_79_io_in_sExp;
  wire [26:0] RoundRawFNToRecFN_79_io_in_sig;
  wire [1:0] RoundRawFNToRecFN_79_io_roundingMode;
  wire [32:0] RoundRawFNToRecFN_79_io_out;
  wire [4:0] RoundRawFNToRecFN_79_io_exceptionFlags;
  RoundRawFNToRecFN RoundRawFNToRecFN_79 (
    .clk(RoundRawFNToRecFN_79_clk),
    .reset(RoundRawFNToRecFN_79_reset),
    .io_invalidExc(RoundRawFNToRecFN_79_io_invalidExc),
    .io_infiniteExc(RoundRawFNToRecFN_79_io_infiniteExc),
    .io_in_sign(RoundRawFNToRecFN_79_io_in_sign),
    .io_in_isNaN(RoundRawFNToRecFN_79_io_in_isNaN),
    .io_in_isInf(RoundRawFNToRecFN_79_io_in_isInf),
    .io_in_isZero(RoundRawFNToRecFN_79_io_in_isZero),
    .io_in_sExp(RoundRawFNToRecFN_79_io_in_sExp),
    .io_in_sig(RoundRawFNToRecFN_79_io_in_sig),
    .io_roundingMode(RoundRawFNToRecFN_79_io_roundingMode),
    .io_out(RoundRawFNToRecFN_79_io_out),
    .io_exceptionFlags(RoundRawFNToRecFN_79_io_exceptionFlags)
  );
  assign io_out = RoundRawFNToRecFN_79_io_out;
  assign io_exceptionFlags = RoundRawFNToRecFN_79_io_exceptionFlags;
  assign T_4 = io_in[63:52];
  assign T_5 = T_4[11:10];
  assign T_7 = T_5 == 2'h3;
  assign T_15_sign = T_22;
  assign T_15_isNaN = T_24;
  assign T_15_isInf = T_28;
  assign T_15_isZero = T_31;
  assign T_15_sExp = T_32;
  assign T_15_sig = T_37;
  assign T_22 = io_in[64];
  assign T_23 = T_4[9];
  assign T_24 = T_7 & T_23;
  assign T_27 = T_23 == 1'h0;
  assign T_28 = T_7 & T_27;
  assign T_29 = T_4[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_31 = T_29 == GEN_0;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_34 = io_in[51:0];
  assign T_36 = {2'h1,T_34};
  assign T_37 = {T_36,2'h0};
  assign GEN_1 = $signed(12'h900);
  assign GEN_2 = {{1{GEN_1[11]}},GEN_1};
  assign T_39 = $signed(T_15_sExp) + $signed(GEN_2);
  assign T_40 = T_39[12:0];
  assign T_41 = $signed(T_40);
  assign outRawFloat_sign = T_15_sign;
  assign outRawFloat_isNaN = T_15_isNaN;
  assign outRawFloat_isInf = T_15_isInf;
  assign outRawFloat_isZero = T_15_isZero;
  assign outRawFloat_sExp = T_70;
  assign outRawFloat_sig = T_75;
  assign GEN_3 = $signed(1'h0);
  assign GEN_4 = {13{GEN_3}};
  assign T_56 = $signed(T_41) < $signed(GEN_4);
  assign T_57 = T_41[11:9];
  assign T_59 = T_57 != GEN_0;
  assign T_67 = T_41[8:0];
  assign T_68 = T_59 ? 9'h1fc : T_67;
  assign T_69 = {T_56,T_68};
  assign T_70 = $signed(T_69);
  assign T_71 = T_15_sig[55:30];
  assign T_72 = T_15_sig[29:0];
  assign GEN_6 = {{29'd0}, 1'h0};
  assign T_74 = T_72 != GEN_6;
  assign T_75 = {T_71,T_74};
  assign T_76 = outRawFloat_sig[24];
  assign T_78 = T_76 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_78;
  assign RoundRawFNToRecFN_79_clk = clk;
  assign RoundRawFNToRecFN_79_reset = reset;
  assign RoundRawFNToRecFN_79_io_invalidExc = invalidExc;
  assign RoundRawFNToRecFN_79_io_infiniteExc = 1'h0;
  assign RoundRawFNToRecFN_79_io_in_sign = outRawFloat_sign;
  assign RoundRawFNToRecFN_79_io_in_isNaN = outRawFloat_isNaN;
  assign RoundRawFNToRecFN_79_io_in_isInf = outRawFloat_isInf;
  assign RoundRawFNToRecFN_79_io_in_isZero = outRawFloat_isZero;
  assign RoundRawFNToRecFN_79_io_in_sExp = outRawFloat_sExp;
  assign RoundRawFNToRecFN_79_io_in_sig = outRawFloat_sig;
  assign RoundRawFNToRecFN_79_io_roundingMode = io_roundingMode;
endmodule
module FPToFP(
  input   clk,
  input   reset,
  input   io_in_valid,
  input  [4:0] io_in_bits_cmd,
  input   io_in_bits_ldst,
  input   io_in_bits_wen,
  input   io_in_bits_ren1,
  input   io_in_bits_ren2,
  input   io_in_bits_ren3,
  input   io_in_bits_swap12,
  input   io_in_bits_swap23,
  input   io_in_bits_single,
  input   io_in_bits_fromint,
  input   io_in_bits_toint,
  input   io_in_bits_fastpipe,
  input   io_in_bits_fma,
  input   io_in_bits_div,
  input   io_in_bits_sqrt,
  input   io_in_bits_round,
  input   io_in_bits_wflags,
  input  [2:0] io_in_bits_rm,
  input  [1:0] io_in_bits_typ,
  input  [64:0] io_in_bits_in1,
  input  [64:0] io_in_bits_in2,
  input  [64:0] io_in_bits_in3,
  output  io_out_valid,
  output [64:0] io_out_bits_data,
  output [4:0] io_out_bits_exc,
  input   io_lt
);
  reg  T_133;
  reg [31:0] GEN_35;
  reg [4:0] T_134_cmd;
  reg [31:0] GEN_36;
  reg  T_134_ldst;
  reg [31:0] GEN_37;
  reg  T_134_wen;
  reg [31:0] GEN_38;
  reg  T_134_ren1;
  reg [31:0] GEN_41;
  reg  T_134_ren2;
  reg [31:0] GEN_42;
  reg  T_134_ren3;
  reg [31:0] GEN_43;
  reg  T_134_swap12;
  reg [31:0] GEN_44;
  reg  T_134_swap23;
  reg [31:0] GEN_45;
  reg  T_134_single;
  reg [31:0] GEN_46;
  reg  T_134_fromint;
  reg [31:0] GEN_47;
  reg  T_134_toint;
  reg [31:0] GEN_48;
  reg  T_134_fastpipe;
  reg [31:0] GEN_49;
  reg  T_134_fma;
  reg [31:0] GEN_50;
  reg  T_134_div;
  reg [31:0] GEN_51;
  reg  T_134_sqrt;
  reg [31:0] GEN_52;
  reg  T_134_round;
  reg [31:0] GEN_53;
  reg  T_134_wflags;
  reg [31:0] GEN_54;
  reg [2:0] T_134_rm;
  reg [31:0] GEN_55;
  reg [1:0] T_134_typ;
  reg [31:0] GEN_56;
  reg [64:0] T_134_in1;
  reg [95:0] GEN_57;
  reg [64:0] T_134_in2;
  reg [95:0] GEN_58;
  reg [64:0] T_134_in3;
  reg [95:0] GEN_59;
  wire [4:0] GEN_0;
  wire  GEN_1;
  wire  GEN_2;
  wire  GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire [2:0] GEN_17;
  wire [1:0] GEN_18;
  wire [64:0] GEN_19;
  wire [64:0] GEN_20;
  wire [64:0] GEN_21;
  wire  in_valid;
  wire [4:0] in_bits_cmd;
  wire  in_bits_ldst;
  wire  in_bits_wen;
  wire  in_bits_ren1;
  wire  in_bits_ren2;
  wire  in_bits_ren3;
  wire  in_bits_swap12;
  wire  in_bits_swap23;
  wire  in_bits_single;
  wire  in_bits_fromint;
  wire  in_bits_toint;
  wire  in_bits_fastpipe;
  wire  in_bits_fma;
  wire  in_bits_div;
  wire  in_bits_sqrt;
  wire  in_bits_round;
  wire  in_bits_wflags;
  wire [2:0] in_bits_rm;
  wire [1:0] in_bits_typ;
  wire [64:0] in_bits_in1;
  wire [64:0] in_bits_in2;
  wire [64:0] in_bits_in3;
  wire [4:0] GEN_32;
  wire [4:0] T_254;
  wire [4:0] GEN_33;
  wire  isSgnj;
  wire  T_255;
  wire  T_256;
  wire  T_258;
  wire  T_259;
  wire  T_260;
  wire  T_261;
  wire  T_262;
  wire  T_263;
  wire  T_264;
  wire  sign_s;
  wire  T_266;
  wire  T_267;
  wire  T_270;
  wire  T_271;
  wire  T_272;
  wire  T_274;
  wire  T_275;
  wire  T_276;
  wire  sign_d;
  wire [30:0] T_277;
  wire [31:0] T_278;
  wire [32:0] T_279;
  wire [31:0] T_280;
  wire [64:0] fsgnj;
  wire  s2d_clk;
  wire  s2d_reset;
  wire [32:0] s2d_io_in;
  wire [1:0] s2d_io_roundingMode;
  wire [64:0] s2d_io_out;
  wire [4:0] s2d_io_exceptionFlags;
  wire  d2s_clk;
  wire  d2s_reset;
  wire [64:0] d2s_io_in;
  wire [1:0] d2s_io_roundingMode;
  wire [32:0] d2s_io_out;
  wire [4:0] d2s_io_exceptionFlags;
  wire [2:0] T_281;
  wire [2:0] T_282;
  wire [2:0] GEN_34;
  wire  T_284;
  wire [2:0] T_285;
  wire [2:0] T_286;
  wire  T_288;
  wire  isnan1;
  wire [2:0] T_289;
  wire [2:0] T_290;
  wire  T_292;
  wire [2:0] T_293;
  wire [2:0] T_294;
  wire  T_296;
  wire  isnan2;
  wire  T_297;
  wire  T_298;
  wire  T_299;
  wire  T_300;
  wire  issnan1;
  wire  T_301;
  wire  T_302;
  wire  T_303;
  wire  T_304;
  wire  issnan2;
  wire  T_305;
  wire [4:0] minmax_exc;
  wire  T_307;
  wire  T_309;
  wire  T_310;
  wire  isLHS;
  wire [64:0] mux_data;
  wire [4:0] mux_exc;
  wire [4:0] GEN_22;
  wire  T_317;
  wire [64:0] GEN_23;
  wire [4:0] T_320;
  wire [4:0] GEN_39;
  wire  T_321;
  wire [31:0] GEN_40;
  wire [31:0] T_323;
  wire [64:0] T_324;
  wire [64:0] GEN_24;
  wire [4:0] GEN_25;
  wire [64:0] GEN_26;
  wire [4:0] GEN_27;
  wire [64:0] GEN_28;
  wire [4:0] GEN_29;
  reg  T_329;
  reg [31:0] GEN_60;
  reg [64:0] T_330_data;
  reg [95:0] GEN_61;
  reg [4:0] T_330_exc;
  reg [31:0] GEN_62;
  wire [64:0] GEN_30;
  wire [4:0] GEN_31;
  wire  T_341_valid;
  wire [64:0] T_341_bits_data;
  wire [4:0] T_341_bits_exc;
  RecFNToRecFN s2d (
    .clk(s2d_clk),
    .reset(s2d_reset),
    .io_in(s2d_io_in),
    .io_roundingMode(s2d_io_roundingMode),
    .io_out(s2d_io_out),
    .io_exceptionFlags(s2d_io_exceptionFlags)
  );
  RecFNToRecFN_98 d2s (
    .clk(d2s_clk),
    .reset(d2s_reset),
    .io_in(d2s_io_in),
    .io_roundingMode(d2s_io_roundingMode),
    .io_out(d2s_io_out),
    .io_exceptionFlags(d2s_io_exceptionFlags)
  );
  assign io_out_valid = T_341_valid;
  assign io_out_bits_data = T_341_bits_data;
  assign io_out_bits_exc = T_341_bits_exc;
  assign GEN_0 = io_in_valid ? io_in_bits_cmd : T_134_cmd;
  assign GEN_1 = io_in_valid ? io_in_bits_ldst : T_134_ldst;
  assign GEN_2 = io_in_valid ? io_in_bits_wen : T_134_wen;
  assign GEN_3 = io_in_valid ? io_in_bits_ren1 : T_134_ren1;
  assign GEN_4 = io_in_valid ? io_in_bits_ren2 : T_134_ren2;
  assign GEN_5 = io_in_valid ? io_in_bits_ren3 : T_134_ren3;
  assign GEN_6 = io_in_valid ? io_in_bits_swap12 : T_134_swap12;
  assign GEN_7 = io_in_valid ? io_in_bits_swap23 : T_134_swap23;
  assign GEN_8 = io_in_valid ? io_in_bits_single : T_134_single;
  assign GEN_9 = io_in_valid ? io_in_bits_fromint : T_134_fromint;
  assign GEN_10 = io_in_valid ? io_in_bits_toint : T_134_toint;
  assign GEN_11 = io_in_valid ? io_in_bits_fastpipe : T_134_fastpipe;
  assign GEN_12 = io_in_valid ? io_in_bits_fma : T_134_fma;
  assign GEN_13 = io_in_valid ? io_in_bits_div : T_134_div;
  assign GEN_14 = io_in_valid ? io_in_bits_sqrt : T_134_sqrt;
  assign GEN_15 = io_in_valid ? io_in_bits_round : T_134_round;
  assign GEN_16 = io_in_valid ? io_in_bits_wflags : T_134_wflags;
  assign GEN_17 = io_in_valid ? io_in_bits_rm : T_134_rm;
  assign GEN_18 = io_in_valid ? io_in_bits_typ : T_134_typ;
  assign GEN_19 = io_in_valid ? io_in_bits_in1 : T_134_in1;
  assign GEN_20 = io_in_valid ? io_in_bits_in2 : T_134_in2;
  assign GEN_21 = io_in_valid ? io_in_bits_in3 : T_134_in3;
  assign in_valid = T_133;
  assign in_bits_cmd = T_134_cmd;
  assign in_bits_ldst = T_134_ldst;
  assign in_bits_wen = T_134_wen;
  assign in_bits_ren1 = T_134_ren1;
  assign in_bits_ren2 = T_134_ren2;
  assign in_bits_ren3 = T_134_ren3;
  assign in_bits_swap12 = T_134_swap12;
  assign in_bits_swap23 = T_134_swap23;
  assign in_bits_single = T_134_single;
  assign in_bits_fromint = T_134_fromint;
  assign in_bits_toint = T_134_toint;
  assign in_bits_fastpipe = T_134_fastpipe;
  assign in_bits_fma = T_134_fma;
  assign in_bits_div = T_134_div;
  assign in_bits_sqrt = T_134_sqrt;
  assign in_bits_round = T_134_round;
  assign in_bits_wflags = T_134_wflags;
  assign in_bits_rm = T_134_rm;
  assign in_bits_typ = T_134_typ;
  assign in_bits_in1 = T_134_in1;
  assign in_bits_in2 = T_134_in2;
  assign in_bits_in3 = T_134_in3;
  assign GEN_32 = {{2'd0}, 3'h5};
  assign T_254 = in_bits_cmd & GEN_32;
  assign GEN_33 = {{2'd0}, 3'h4};
  assign isSgnj = GEN_33 == T_254;
  assign T_255 = in_bits_single & isSgnj;
  assign T_256 = in_bits_rm[1];
  assign T_258 = T_255 == 1'h0;
  assign T_259 = T_256 | T_258;
  assign T_260 = in_bits_in1[32];
  assign T_261 = in_bits_rm[0];
  assign T_262 = T_259 ? T_260 : T_261;
  assign T_263 = in_bits_in2[32];
  assign T_264 = T_255 & T_263;
  assign sign_s = T_262 ^ T_264;
  assign T_266 = in_bits_single == 1'h0;
  assign T_267 = T_266 & isSgnj;
  assign T_270 = T_267 == 1'h0;
  assign T_271 = T_256 | T_270;
  assign T_272 = in_bits_in1[64];
  assign T_274 = T_271 ? T_272 : T_261;
  assign T_275 = in_bits_in2[64];
  assign T_276 = T_267 & T_275;
  assign sign_d = T_274 ^ T_276;
  assign T_277 = in_bits_in1[63:33];
  assign T_278 = in_bits_in1[31:0];
  assign T_279 = {sign_s,T_278};
  assign T_280 = {sign_d,T_277};
  assign fsgnj = {T_280,T_279};
  assign s2d_clk = clk;
  assign s2d_reset = reset;
  assign s2d_io_in = in_bits_in1[32:0];
  assign s2d_io_roundingMode = in_bits_rm[1:0];
  assign d2s_clk = clk;
  assign d2s_reset = reset;
  assign d2s_io_in = in_bits_in1;
  assign d2s_io_roundingMode = in_bits_rm[1:0];
  assign T_281 = in_bits_in1[31:29];
  assign T_282 = ~ T_281;
  assign GEN_34 = {{2'd0}, 1'h0};
  assign T_284 = T_282 == GEN_34;
  assign T_285 = in_bits_in1[63:61];
  assign T_286 = ~ T_285;
  assign T_288 = T_286 == GEN_34;
  assign isnan1 = in_bits_single ? T_284 : T_288;
  assign T_289 = in_bits_in2[31:29];
  assign T_290 = ~ T_289;
  assign T_292 = T_290 == GEN_34;
  assign T_293 = in_bits_in2[63:61];
  assign T_294 = ~ T_293;
  assign T_296 = T_294 == GEN_34;
  assign isnan2 = in_bits_single ? T_292 : T_296;
  assign T_297 = in_bits_in1[22];
  assign T_298 = in_bits_in1[51];
  assign T_299 = in_bits_single ? T_297 : T_298;
  assign T_300 = ~ T_299;
  assign issnan1 = isnan1 & T_300;
  assign T_301 = in_bits_in2[22];
  assign T_302 = in_bits_in2[51];
  assign T_303 = in_bits_single ? T_301 : T_302;
  assign T_304 = ~ T_303;
  assign issnan2 = isnan2 & T_304;
  assign T_305 = issnan1 | issnan2;
  assign minmax_exc = {T_305,4'h0};
  assign T_307 = T_261 != io_lt;
  assign T_309 = isnan1 == 1'h0;
  assign T_310 = T_307 & T_309;
  assign isLHS = isnan2 | T_310;
  assign mux_data = GEN_28;
  assign mux_exc = GEN_29;
  assign GEN_22 = isSgnj ? {{4'd0}, 1'h0} : minmax_exc;
  assign T_317 = isSgnj | isLHS;
  assign GEN_23 = T_317 ? fsgnj : in_bits_in2;
  assign T_320 = in_bits_cmd & GEN_33;
  assign GEN_39 = {{4'd0}, 1'h0};
  assign T_321 = GEN_39 == T_320;
  assign GEN_40 = $signed(32'hffffffff);
  assign T_323 = $unsigned(GEN_40);
  assign T_324 = {T_323,d2s_io_out};
  assign GEN_24 = in_bits_single ? T_324 : GEN_23;
  assign GEN_25 = in_bits_single ? d2s_io_exceptionFlags : GEN_22;
  assign GEN_26 = T_266 ? s2d_io_out : GEN_24;
  assign GEN_27 = T_266 ? s2d_io_exceptionFlags : GEN_25;
  assign GEN_28 = T_321 ? GEN_26 : GEN_23;
  assign GEN_29 = T_321 ? GEN_27 : GEN_22;
  assign GEN_30 = in_valid ? mux_data : T_330_data;
  assign GEN_31 = in_valid ? mux_exc : T_330_exc;
  assign T_341_valid = T_329;
  assign T_341_bits_data = T_330_data;
  assign T_341_bits_exc = T_330_exc;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_35 = {1{$random}};
  T_133 = GEN_35[0:0];
  GEN_36 = {1{$random}};
  T_134_cmd = GEN_36[4:0];
  GEN_37 = {1{$random}};
  T_134_ldst = GEN_37[0:0];
  GEN_38 = {1{$random}};
  T_134_wen = GEN_38[0:0];
  GEN_41 = {1{$random}};
  T_134_ren1 = GEN_41[0:0];
  GEN_42 = {1{$random}};
  T_134_ren2 = GEN_42[0:0];
  GEN_43 = {1{$random}};
  T_134_ren3 = GEN_43[0:0];
  GEN_44 = {1{$random}};
  T_134_swap12 = GEN_44[0:0];
  GEN_45 = {1{$random}};
  T_134_swap23 = GEN_45[0:0];
  GEN_46 = {1{$random}};
  T_134_single = GEN_46[0:0];
  GEN_47 = {1{$random}};
  T_134_fromint = GEN_47[0:0];
  GEN_48 = {1{$random}};
  T_134_toint = GEN_48[0:0];
  GEN_49 = {1{$random}};
  T_134_fastpipe = GEN_49[0:0];
  GEN_50 = {1{$random}};
  T_134_fma = GEN_50[0:0];
  GEN_51 = {1{$random}};
  T_134_div = GEN_51[0:0];
  GEN_52 = {1{$random}};
  T_134_sqrt = GEN_52[0:0];
  GEN_53 = {1{$random}};
  T_134_round = GEN_53[0:0];
  GEN_54 = {1{$random}};
  T_134_wflags = GEN_54[0:0];
  GEN_55 = {1{$random}};
  T_134_rm = GEN_55[2:0];
  GEN_56 = {1{$random}};
  T_134_typ = GEN_56[1:0];
  GEN_57 = {3{$random}};
  T_134_in1 = GEN_57[64:0];
  GEN_58 = {3{$random}};
  T_134_in2 = GEN_58[64:0];
  GEN_59 = {3{$random}};
  T_134_in3 = GEN_59[64:0];
  GEN_60 = {1{$random}};
  T_329 = GEN_60[0:0];
  GEN_61 = {3{$random}};
  T_330_data = GEN_61[64:0];
  GEN_62 = {1{$random}};
  T_330_exc = GEN_62[4:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      T_133 <= 1'h0;
    end else begin
      T_133 <= io_in_valid;
    end
    if(1'h0) begin
    end else begin
      T_134_cmd <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      T_134_ldst <= GEN_1;
    end
    if(1'h0) begin
    end else begin
      T_134_wen <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      T_134_ren1 <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      T_134_ren2 <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      T_134_ren3 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      T_134_swap12 <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      T_134_swap23 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      T_134_single <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      T_134_fromint <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      T_134_toint <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      T_134_fastpipe <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      T_134_fma <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      T_134_div <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      T_134_sqrt <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      T_134_round <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_134_wflags <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      T_134_rm <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      T_134_typ <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      T_134_in1 <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      T_134_in2 <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      T_134_in3 <= GEN_21;
    end
    if(reset) begin
      T_329 <= 1'h0;
    end else begin
      T_329 <= in_valid;
    end
    if(1'h0) begin
    end else begin
      T_330_data <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      T_330_exc <= GEN_31;
    end
  end
endmodule
module DivSqrtRecF64_mulAddZ31(
  input   clk,
  input   reset,
  output  io_inReady_div,
  output  io_inReady_sqrt,
  input   io_inValid,
  input   io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [1:0] io_roundingMode,
  output  io_outValid_div,
  output  io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags,
  output [3:0] io_usingMulAdd,
  output  io_latchMulAddA_0,
  output [53:0] io_mulAddA_0,
  output  io_latchMulAddB_0,
  output [53:0] io_mulAddB_0,
  output [104:0] io_mulAddC_2,
  input  [104:0] io_mulAddResult_3
);
  reg  valid_PA;
  reg [31:0] GEN_61;
  reg  sqrtOp_PA;
  reg [31:0] GEN_70;
  reg  sign_PA;
  reg [31:0] GEN_71;
  reg [2:0] specialCodeB_PA;
  reg [31:0] GEN_72;
  reg  fractB_51_PA;
  reg [31:0] GEN_73;
  reg [1:0] roundingMode_PA;
  reg [31:0] GEN_74;
  reg [2:0] specialCodeA_PA;
  reg [31:0] GEN_75;
  reg  fractA_51_PA;
  reg [31:0] GEN_76;
  reg [13:0] exp_PA;
  reg [31:0] GEN_77;
  reg [50:0] fractB_other_PA;
  reg [63:0] GEN_78;
  reg [50:0] fractA_other_PA;
  reg [63:0] GEN_79;
  reg  valid_PB;
  reg [31:0] GEN_80;
  reg  sqrtOp_PB;
  reg [31:0] GEN_81;
  reg  sign_PB;
  reg [31:0] GEN_82;
  reg [2:0] specialCodeA_PB;
  reg [31:0] GEN_83;
  reg  fractA_51_PB;
  reg [31:0] GEN_84;
  reg [2:0] specialCodeB_PB;
  reg [31:0] GEN_157;
  reg  fractB_51_PB;
  reg [31:0] GEN_158;
  reg [1:0] roundingMode_PB;
  reg [31:0] GEN_159;
  reg [13:0] exp_PB;
  reg [31:0] GEN_163;
  reg  fractA_0_PB;
  reg [31:0] GEN_166;
  reg [50:0] fractB_other_PB;
  reg [63:0] GEN_167;
  reg  valid_PC;
  reg [31:0] GEN_168;
  reg  sqrtOp_PC;
  reg [31:0] GEN_169;
  reg  sign_PC;
  reg [31:0] GEN_170;
  reg [2:0] specialCodeA_PC;
  reg [31:0] GEN_171;
  reg  fractA_51_PC;
  reg [31:0] GEN_172;
  reg [2:0] specialCodeB_PC;
  reg [31:0] GEN_173;
  reg  fractB_51_PC;
  reg [31:0] GEN_174;
  reg [1:0] roundingMode_PC;
  reg [31:0] GEN_175;
  reg [13:0] exp_PC;
  reg [31:0] GEN_176;
  reg  fractA_0_PC;
  reg [31:0] GEN_177;
  reg [50:0] fractB_other_PC;
  reg [63:0] GEN_178;
  reg [2:0] cycleNum_A;
  reg [31:0] GEN_179;
  reg [3:0] cycleNum_B;
  reg [31:0] GEN_180;
  reg [2:0] cycleNum_C;
  reg [31:0] GEN_181;
  reg [2:0] cycleNum_E;
  reg [31:0] GEN_182;
  reg [8:0] fractR0_A;
  reg [31:0] GEN_183;
  reg [9:0] hiSqrR0_A_sqrt;
  reg [31:0] GEN_184;
  reg [20:0] partNegSigma0_A;
  reg [31:0] GEN_185;
  reg [8:0] nextMulAdd9A_A;
  reg [31:0] GEN_186;
  reg [8:0] nextMulAdd9B_A;
  reg [31:0] GEN_187;
  reg [16:0] ER1_B_sqrt;
  reg [31:0] GEN_188;
  reg [31:0] ESqrR1_B_sqrt;
  reg [31:0] GEN_189;
  reg [57:0] sigX1_B;
  reg [63:0] GEN_190;
  reg [32:0] sqrSigma1_C;
  reg [63:0] GEN_191;
  reg [57:0] sigXN_C;
  reg [63:0] GEN_192;
  reg [30:0] u_C_sqrt;
  reg [31:0] GEN_193;
  reg  E_E_div;
  reg [31:0] GEN_194;
  reg [52:0] sigT_E;
  reg [63:0] GEN_195;
  reg  extraT_E;
  reg [31:0] GEN_196;
  reg  isNegRemT_E;
  reg [31:0] GEN_197;
  reg  trueEqX_E1;
  reg [31:0] GEN_198;
  wire  ready_PA;
  wire  ready_PB;
  wire  ready_PC;
  wire  leaving_PA;
  wire  leaving_PB;
  wire  leaving_PC;
  wire  cyc_B10_sqrt;
  wire  cyc_B9_sqrt;
  wire  cyc_B8_sqrt;
  wire  cyc_B7_sqrt;
  wire  cyc_B6;
  wire  cyc_B5;
  wire  cyc_B4;
  wire  cyc_B3;
  wire  cyc_B2;
  wire  cyc_B1;
  wire  cyc_B6_div;
  wire  cyc_B5_div;
  wire  cyc_B4_div;
  wire  cyc_B3_div;
  wire  cyc_B2_div;
  wire  cyc_B1_div;
  wire  cyc_B6_sqrt;
  wire  cyc_B5_sqrt;
  wire  cyc_B4_sqrt;
  wire  cyc_B3_sqrt;
  wire  cyc_B2_sqrt;
  wire  cyc_B1_sqrt;
  wire  cyc_C5;
  wire  cyc_C4;
  wire  valid_normalCase_leaving_PB;
  wire  cyc_C2;
  wire  cyc_C1;
  wire  cyc_E4;
  wire  cyc_E3;
  wire  cyc_E2;
  wire  cyc_E1;
  wire [45:0] zSigma1_B4;
  wire [57:0] sigXNU_B3_CX;
  wire [53:0] zComplSigT_C1_sqrt;
  wire [53:0] zComplSigT_C1;
  wire  T_113;
  wire  T_114;
  wire  T_116;
  wire  T_117;
  wire  T_119;
  wire  T_120;
  wire  T_122;
  wire  T_123;
  wire  T_125;
  wire  T_126;
  wire  T_128;
  wire  T_129;
  wire  T_131;
  wire  T_132;
  wire  T_134;
  wire  T_135;
  wire  T_137;
  wire  T_138;
  wire  T_141;
  wire  T_144;
  wire  T_147;
  wire  T_149;
  wire  T_150;
  wire  T_153;
  wire  T_154;
  wire  T_156;
  wire  cyc_S_div;
  wire  T_157;
  wire  cyc_S_sqrt;
  wire  cyc_S;
  wire  signA_S;
  wire [11:0] expA_S;
  wire [51:0] fractA_S;
  wire [2:0] specialCodeA_S;
  wire  isZeroA_S;
  wire [1:0] T_159;
  wire  isSpecialA_S;
  wire  signB_S;
  wire [11:0] expB_S;
  wire [51:0] fractB_S;
  wire [2:0] specialCodeB_S;
  wire  isZeroB_S;
  wire [1:0] T_162;
  wire  isSpecialB_S;
  wire  T_164;
  wire  sign_S;
  wire  T_166;
  wire  T_168;
  wire  T_169;
  wire  T_171;
  wire  T_172;
  wire  T_174;
  wire  normalCase_S_div;
  wire  T_179;
  wire  T_181;
  wire  normalCase_S_sqrt;
  wire  normalCase_S;
  wire  entering_PA_normalCase_div;
  wire  entering_PA_normalCase_sqrt;
  wire  entering_PA_normalCase;
  wire  T_183;
  wire  T_184;
  wire  T_185;
  wire  entering_PA;
  wire  T_187;
  wire  T_188;
  wire  T_190;
  wire  T_191;
  wire  T_193;
  wire  T_195;
  wire  T_196;
  wire  T_197;
  wire  entering_PB_S;
  wire  T_206;
  wire  entering_PC_S;
  wire  T_207;
  wire  GEN_0;
  wire  T_208;
  wire  GEN_1;
  wire  GEN_2;
  wire [2:0] GEN_3;
  wire  GEN_4;
  wire [1:0] GEN_5;
  wire  T_211;
  wire  T_212;
  wire [2:0] GEN_6;
  wire  GEN_7;
  wire  T_213;
  wire [2:0] GEN_53;
  wire [3:0] T_215;
  wire [2:0] T_216;
  wire [10:0] T_217;
  wire [10:0] T_218;
  wire [13:0] T_219;
  wire [13:0] GEN_54;
  wire [14:0] T_220;
  wire [13:0] T_221;
  wire [13:0] T_222;
  wire [50:0] T_223;
  wire [13:0] GEN_8;
  wire [50:0] GEN_9;
  wire [50:0] T_224;
  wire [50:0] GEN_10;
  wire  isZeroA_PA;
  wire [1:0] T_226;
  wire  isSpecialA_PA;
  wire [1:0] T_229;
  wire [52:0] sigA_PA;
  wire  isZeroB_PA;
  wire [1:0] T_231;
  wire  isSpecialB_PA;
  wire [1:0] T_234;
  wire [52:0] sigB_PA;
  wire  T_236;
  wire  T_238;
  wire  T_239;
  wire  T_241;
  wire  T_242;
  wire  T_244;
  wire  T_247;
  wire  T_249;
  wire  T_250;
  wire  T_253;
  wire  normalCase_PA;
  wire  valid_normalCase_leaving_PA;
  wire  valid_leaving_PA;
  wire  T_254;
  wire  T_257;
  wire  T_258;
  wire  entering_PB_normalCase;
  wire  entering_PB;
  wire  T_259;
  wire  GEN_11;
  wire  T_260;
  wire  T_261;
  wire [2:0] T_262;
  wire  T_264;
  wire [2:0] T_265;
  wire  T_267;
  wire [1:0] T_268;
  wire  GEN_12;
  wire  GEN_13;
  wire [2:0] GEN_14;
  wire  GEN_15;
  wire [2:0] GEN_16;
  wire  GEN_17;
  wire [1:0] GEN_18;
  wire  T_269;
  wire [13:0] GEN_19;
  wire  GEN_20;
  wire [50:0] GEN_21;
  wire  isZeroA_PB;
  wire [1:0] T_271;
  wire  isSpecialA_PB;
  wire  isZeroB_PB;
  wire [1:0] T_274;
  wire  isSpecialB_PB;
  wire  T_277;
  wire  T_279;
  wire  T_280;
  wire  T_282;
  wire  T_283;
  wire  T_285;
  wire  T_288;
  wire  T_290;
  wire  T_291;
  wire  T_294;
  wire  normalCase_PB;
  wire  valid_leaving_PB;
  wire  T_295;
  wire  T_298;
  wire  T_299;
  wire  entering_PC_normalCase;
  wire  entering_PC;
  wire  T_300;
  wire  GEN_22;
  wire  T_301;
  wire  T_302;
  wire [2:0] T_303;
  wire  T_305;
  wire [2:0] T_306;
  wire  T_308;
  wire [1:0] T_309;
  wire  GEN_23;
  wire  GEN_24;
  wire [2:0] GEN_25;
  wire  GEN_26;
  wire [2:0] GEN_27;
  wire  GEN_28;
  wire [1:0] GEN_29;
  wire [13:0] GEN_30;
  wire  GEN_31;
  wire [50:0] GEN_32;
  wire  isZeroA_PC;
  wire [1:0] T_311;
  wire  isSpecialA_PC;
  wire  T_313;
  wire  T_315;
  wire  isInfA_PC;
  wire  isNaNA_PC;
  wire  T_318;
  wire  isSigNaNA_PC;
  wire  isZeroB_PC;
  wire [1:0] T_320;
  wire  isSpecialB_PC;
  wire  T_322;
  wire  T_324;
  wire  isInfB_PC;
  wire  isNaNB_PC;
  wire  T_327;
  wire  isSigNaNB_PC;
  wire [1:0] T_329;
  wire [52:0] sigB_PC;
  wire  T_331;
  wire  T_333;
  wire  T_334;
  wire  T_336;
  wire  T_337;
  wire  T_339;
  wire  T_342;
  wire  T_344;
  wire  T_345;
  wire  T_348;
  wire  normalCase_PC;
  wire [13:0] GEN_55;
  wire [14:0] T_350;
  wire [13:0] expP2_PC;
  wire  T_351;
  wire [12:0] T_352;
  wire [13:0] T_354;
  wire [12:0] T_355;
  wire [13:0] T_357;
  wire [13:0] expP1_PC;
  wire  roundingMode_near_even_PC;
  wire  roundingMode_min_PC;
  wire  roundingMode_max_PC;
  wire  roundMagUp_PC;
  wire  overflowY_roundMagUp_PC;
  wire  T_359;
  wire  T_361;
  wire  roundMagDown_PC;
  wire  T_363;
  wire  valid_leaving_PC;
  wire  T_364;
  wire  T_366;
  wire  T_367;
  wire  T_369;
  wire  T_370;
  wire  T_371;
  wire [2:0] GEN_56;
  wire  T_373;
  wire  T_374;
  wire [1:0] T_377;
  wire [2:0] T_380;
  wire [2:0] GEN_57;
  wire [2:0] T_381;
  wire  T_383;
  wire [2:0] GEN_58;
  wire [3:0] T_385;
  wire [2:0] T_386;
  wire [2:0] T_388;
  wire [2:0] T_389;
  wire [2:0] GEN_33;
  wire  cyc_A6_sqrt;
  wire  cyc_A5_sqrt;
  wire  cyc_A4_sqrt;
  wire  cyc_A4;
  wire [2:0] GEN_59;
  wire  cyc_A3;
  wire [2:0] GEN_60;
  wire  cyc_A2;
  wire  cyc_A1;
  wire  T_397;
  wire  cyc_A3_div;
  wire  cyc_A2_div;
  wire  cyc_A1_div;
  wire  cyc_A3_sqrt;
  wire  cyc_A1_sqrt;
  wire [3:0] GEN_62;
  wire  T_403;
  wire  T_404;
  wire [3:0] T_407;
  wire [3:0] GEN_63;
  wire [4:0] T_409;
  wire [3:0] T_410;
  wire [3:0] T_411;
  wire [3:0] GEN_34;
  wire  T_413;
  wire  T_415;
  wire  T_417;
  wire [3:0] GEN_64;
  wire  T_419;
  wire [3:0] GEN_65;
  wire  T_421;
  wire [3:0] GEN_66;
  wire  T_423;
  wire [3:0] GEN_67;
  wire  T_425;
  wire [3:0] GEN_68;
  wire  T_427;
  wire [3:0] GEN_69;
  wire  T_429;
  wire  T_431;
  wire  T_432;
  wire  T_435;
  wire  T_436;
  wire  T_439;
  wire  T_440;
  wire  T_443;
  wire  T_445;
  wire  T_446;
  wire  T_449;
  wire  T_452;
  wire  T_453;
  wire  T_454;
  wire  T_455;
  wire  T_456;
  wire  T_457;
  wire  T_458;
  wire  T_459;
  wire  T_460;
  wire  T_461;
  wire  T_463;
  wire  T_464;
  wire [2:0] T_467;
  wire [3:0] T_469;
  wire [2:0] T_470;
  wire [2:0] T_471;
  wire [2:0] GEN_35;
  wire  cyc_C6_sqrt;
  wire  T_474;
  wire  T_476;
  wire  T_478;
  wire  T_480;
  wire  T_482;
  wire  cyc_C5_div;
  wire  cyc_C4_div;
  wire  cyc_C1_div;
  wire  cyc_C5_sqrt;
  wire  cyc_C4_sqrt;
  wire  cyc_C3_sqrt;
  wire  cyc_C1_sqrt;
  wire  T_494;
  wire  T_495;
  wire [3:0] T_498;
  wire [2:0] T_499;
  wire [2:0] T_500;
  wire [2:0] GEN_36;
  wire  T_502;
  wire  T_504;
  wire  T_506;
  wire  T_508;
  wire  cyc_E3_div;
  wire  cyc_E3_sqrt;
  wire [51:0] zFractB_A4_div;
  wire [2:0] T_518;
  wire  T_520;
  wire  zLinPiece_0_A4_div;
  wire  T_523;
  wire  zLinPiece_1_A4_div;
  wire  T_526;
  wire  zLinPiece_2_A4_div;
  wire  T_529;
  wire  zLinPiece_3_A4_div;
  wire  T_532;
  wire  zLinPiece_4_A4_div;
  wire  T_535;
  wire  zLinPiece_5_A4_div;
  wire  T_538;
  wire  zLinPiece_6_A4_div;
  wire  T_541;
  wire  zLinPiece_7_A4_div;
  wire [8:0] T_544;
  wire [8:0] T_547;
  wire [8:0] T_548;
  wire [8:0] T_551;
  wire [8:0] T_552;
  wire [8:0] T_555;
  wire [8:0] T_556;
  wire [8:0] T_559;
  wire [8:0] T_560;
  wire [8:0] T_563;
  wire [8:0] T_564;
  wire [8:0] T_567;
  wire [8:0] T_568;
  wire [8:0] T_571;
  wire [8:0] zK1_A4_div;
  wire [11:0] T_575;
  wire [11:0] T_579;
  wire [11:0] T_580;
  wire [11:0] T_584;
  wire [11:0] T_585;
  wire [11:0] T_589;
  wire [11:0] T_590;
  wire [11:0] T_594;
  wire [11:0] T_595;
  wire [11:0] T_599;
  wire [11:0] T_600;
  wire [11:0] T_604;
  wire [11:0] T_605;
  wire [11:0] T_609;
  wire [11:0] zComplFractK0_A4_div;
  wire [51:0] zFractB_A7_sqrt;
  wire  T_611;
  wire  T_613;
  wire  T_614;
  wire  T_617;
  wire  zQuadPiece_0_A7_sqrt;
  wire  zQuadPiece_1_A7_sqrt;
  wire  T_624;
  wire  zQuadPiece_2_A7_sqrt;
  wire  zQuadPiece_3_A7_sqrt;
  wire [8:0] T_633;
  wire [8:0] T_636;
  wire [8:0] T_637;
  wire [8:0] T_640;
  wire [8:0] T_641;
  wire [8:0] T_644;
  wire [8:0] zK2_A7_sqrt;
  wire [9:0] T_648;
  wire [9:0] T_652;
  wire [9:0] T_653;
  wire [9:0] T_657;
  wire [9:0] T_658;
  wire [9:0] T_662;
  wire [9:0] zComplK1_A7_sqrt;
  wire  T_663;
  wire  T_665;
  wire  T_666;
  wire  T_667;
  wire  T_669;
  wire  zQuadPiece_0_A6_sqrt;
  wire  zQuadPiece_1_A6_sqrt;
  wire  T_676;
  wire  zQuadPiece_2_A6_sqrt;
  wire  zQuadPiece_3_A6_sqrt;
  wire [12:0] T_686;
  wire [12:0] T_690;
  wire [12:0] T_691;
  wire [12:0] T_695;
  wire [12:0] T_696;
  wire [12:0] T_700;
  wire [12:0] zComplFractK0_A6_sqrt;
  wire [8:0] T_701;
  wire [8:0] T_702;
  wire  T_704;
  wire [8:0] T_706;
  wire [8:0] mulAdd9A_A;
  wire [8:0] T_707;
  wire [8:0] T_708;
  wire [8:0] T_712;
  wire [8:0] mulAdd9B_A;
  wire [9:0] GEN_85;
  wire [10:0] T_714;
  wire [9:0] T_715;
  wire [19:0] T_716;
  wire [5:0] GEN_86;
  wire [6:0] T_718;
  wire [5:0] T_719;
  wire [13:0] T_720;
  wire [19:0] T_721;
  wire [19:0] T_722;
  wire [7:0] GEN_87;
  wire [8:0] T_724;
  wire [7:0] T_725;
  wire [12:0] T_726;
  wire [20:0] T_727;
  wire [20:0] GEN_88;
  wire [20:0] T_728;
  wire [18:0] GEN_89;
  wire [18:0] T_730;
  wire [19:0] GEN_90;
  wire [20:0] T_731;
  wire [19:0] T_732;
  wire [19:0] T_734;
  wire [20:0] GEN_91;
  wire [20:0] T_735;
  wire  T_736;
  wire  T_738;
  wire  T_739;
  wire [10:0] T_742;
  wire [20:0] GEN_92;
  wire [20:0] T_743;
  wire  T_745;
  wire  T_746;
  wire [20:0] T_747;
  wire [20:0] GEN_93;
  wire [21:0] T_749;
  wire [20:0] T_750;
  wire [20:0] T_752;
  wire [20:0] T_753;
  wire  T_754;
  wire [20:0] T_756;
  wire [20:0] T_757;
  wire [24:0] GEN_94;
  wire [24:0] T_758;
  wire [24:0] T_760;
  wire [24:0] GEN_95;
  wire [24:0] T_761;
  wire [23:0] GEN_96;
  wire [23:0] T_762;
  wire [23:0] T_764;
  wire [24:0] GEN_97;
  wire [24:0] mulAdd9C_A;
  wire [17:0] T_765;
  wire [17:0] T_767;
  wire [18:0] T_768;
  wire [18:0] GEN_98;
  wire [19:0] T_769;
  wire [18:0] loMulAdd9Out_A;
  wire  T_770;
  wire [6:0] T_771;
  wire [6:0] GEN_99;
  wire [7:0] T_773;
  wire [6:0] T_774;
  wire [6:0] T_776;
  wire [17:0] T_777;
  wire [24:0] mulAdd9Out_A;
  wire  T_778;
  wire  T_779;
  wire [24:0] T_780;
  wire [14:0] T_781;
  wire [14:0] T_783;
  wire [8:0] zFractR0_A6_sqrt;
  wire [25:0] GEN_100;
  wire [25:0] T_785;
  wire [25:0] sqrR0_A5_sqrt;
  wire  T_786;
  wire  T_787;
  wire [13:0] T_789;
  wire [13:0] T_791;
  wire [8:0] zFractR0_A4_div;
  wire  T_792;
  wire  T_793;
  wire [22:0] T_795;
  wire [22:0] T_797;
  wire [8:0] zSigma0_A2;
  wire [14:0] T_798;
  wire [15:0] T_799;
  wire [15:0] T_800;
  wire [14:0] fractR1_A1;
  wire [15:0] r1_A1;
  wire [16:0] GEN_101;
  wire [16:0] T_803;
  wire [16:0] ER1_A1_sqrt;
  wire  T_804;
  wire [8:0] T_805;
  wire [8:0] GEN_37;
  wire [15:0] T_806;
  wire [15:0] GEN_38;
  wire  T_807;
  wire [24:0] T_809;
  wire [20:0] T_810;
  wire [20:0] GEN_39;
  wire  T_811;
  wire  T_812;
  wire  T_813;
  wire  T_814;
  wire  T_815;
  wire [13:0] T_819;
  wire [13:0] GEN_102;
  wire [13:0] T_820;
  wire [8:0] T_821;
  wire [8:0] T_823;
  wire [13:0] GEN_103;
  wire [13:0] T_824;
  wire [8:0] T_825;
  wire [13:0] GEN_104;
  wire [13:0] T_826;
  wire  T_827;
  wire [8:0] T_828;
  wire [8:0] T_830;
  wire [13:0] GEN_105;
  wire [13:0] T_831;
  wire [13:0] GEN_106;
  wire [13:0] T_832;
  wire [13:0] GEN_40;
  wire  T_836;
  wire [8:0] T_838;
  wire [8:0] T_839;
  wire [8:0] T_841;
  wire [8:0] T_842;
  wire [8:0] T_843;
  wire [8:0] T_844;
  wire [8:0] T_846;
  wire [8:0] T_847;
  wire [7:0] T_849;
  wire [8:0] T_850;
  wire [8:0] T_852;
  wire [8:0] T_853;
  wire [8:0] GEN_41;
  wire [16:0] GEN_42;
  wire  T_854;
  wire  T_855;
  wire  T_856;
  wire  T_857;
  wire  T_858;
  wire  T_859;
  wire  T_860;
  wire [52:0] GEN_107;
  wire [52:0] T_861;
  wire [52:0] T_863;
  wire  T_864;
  wire [52:0] T_866;
  wire [52:0] T_867;
  wire [52:0] T_869;
  wire [52:0] T_870;
  wire [33:0] T_871;
  wire [52:0] GEN_108;
  wire [52:0] T_872;
  wire  T_873;
  wire [45:0] T_874;
  wire [45:0] T_876;
  wire [52:0] GEN_109;
  wire [52:0] T_877;
  wire [32:0] T_878;
  wire [45:0] GEN_110;
  wire [45:0] T_879;
  wire [45:0] T_881;
  wire [52:0] GEN_111;
  wire [52:0] T_882;
  wire [45:0] GEN_112;
  wire [45:0] T_883;
  wire [45:0] T_885;
  wire [52:0] GEN_113;
  wire [52:0] T_886;
  wire [52:0] T_888;
  wire [52:0] T_889;
  wire [53:0] GEN_114;
  wire [53:0] T_890;
  wire  T_892;
  wire  T_893;
  wire  T_894;
  wire  T_895;
  wire  T_896;
  wire [51:0] GEN_115;
  wire [51:0] T_897;
  wire [51:0] T_899;
  wire [50:0] GEN_116;
  wire [50:0] T_900;
  wire [50:0] T_902;
  wire [51:0] GEN_117;
  wire [51:0] T_903;
  wire [52:0] GEN_118;
  wire [52:0] T_904;
  wire [52:0] T_906;
  wire [52:0] GEN_119;
  wire [52:0] T_907;
  wire [52:0] GEN_120;
  wire [52:0] T_908;
  wire [29:0] T_909;
  wire [29:0] T_911;
  wire [52:0] GEN_121;
  wire [52:0] T_912;
  wire [32:0] T_914;
  wire [52:0] GEN_122;
  wire [52:0] T_915;
  wire [53:0] GEN_123;
  wire [53:0] T_916;
  wire  T_917;
  wire  T_918;
  wire  T_919;
  wire  T_920;
  wire  T_921;
  wire  T_922;
  wire  T_923;
  wire  T_924;
  wire  T_925;
  wire  T_926;
  wire  T_927;
  wire  T_928;
  wire  T_929;
  wire  T_930;
  wire  T_931;
  wire  T_932;
  wire  T_933;
  wire  T_934;
  wire  T_935;
  wire  T_936;
  wire  T_937;
  wire  T_938;
  wire  T_939;
  wire  T_940;
  wire  T_941;
  wire  T_942;
  wire  T_943;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_947;
  wire  T_948;
  wire [1:0] T_949;
  wire [1:0] T_950;
  wire [3:0] T_951;
  wire [104:0] GEN_124;
  wire [104:0] T_952;
  wire [104:0] T_954;
  wire [103:0] GEN_125;
  wire [103:0] T_955;
  wire [103:0] T_957;
  wire [104:0] GEN_126;
  wire [104:0] T_958;
  wire  T_959;
  wire [104:0] GEN_127;
  wire [104:0] T_960;
  wire [104:0] T_962;
  wire [104:0] T_963;
  wire  T_965;
  wire  T_966;
  wire [53:0] GEN_128;
  wire [53:0] T_967;
  wire [53:0] T_969;
  wire [104:0] GEN_129;
  wire [104:0] T_970;
  wire  T_972;
  wire [1:0] T_974;
  wire  T_975;
  wire  T_977;
  wire [1:0] T_979;
  wire [1:0] T_980;
  wire  T_982;
  wire [1:0] T_984;
  wire [1:0] T_985;
  wire [55:0] GEN_130;
  wire [55:0] T_986;
  wire [55:0] T_988;
  wire [104:0] GEN_131;
  wire [104:0] T_989;
  wire [31:0] ESqrR1_B8_sqrt;
  wire [45:0] T_990;
  wire [45:0] T_991;
  wire [45:0] T_993;
  wire [32:0] sqrSigma1_B1;
  wire [57:0] T_994;
  wire  T_995;
  wire  E_C1_div;
  wire  T_998;
  wire  T_999;
  wire  T_1000;
  wire [53:0] T_1001;
  wire [53:0] T_1002;
  wire [53:0] T_1004;
  wire  T_1005;
  wire [52:0] T_1007;
  wire [52:0] T_1008;
  wire [53:0] T_1009;
  wire [53:0] T_1011;
  wire [53:0] T_1012;
  wire [53:0] T_1016;
  wire [53:0] sigT_C1;
  wire [55:0] remT_E2;
  wire [31:0] GEN_43;
  wire [57:0] GEN_44;
  wire [32:0] GEN_45;
  wire  T_1017;
  wire  T_1018;
  wire [57:0] GEN_46;
  wire [30:0] T_1019;
  wire [30:0] GEN_47;
  wire [52:0] T_1020;
  wire  T_1021;
  wire  GEN_48;
  wire [52:0] GEN_49;
  wire  GEN_50;
  wire  T_1022;
  wire  T_1023;
  wire  T_1024;
  wire [53:0] T_1025;
  wire [53:0] GEN_132;
  wire  T_1027;
  wire [1:0] T_1030;
  wire [1:0] GEN_133;
  wire  T_1032;
  wire  T_1033;
  wire  T_1034;
  wire  GEN_51;
  wire  GEN_52;
  wire  T_1037;
  wire [13:0] T_1039;
  wire  T_1044;
  wire [13:0] T_1046;
  wire [13:0] T_1047;
  wire [12:0] T_1048;
  wire [12:0] GEN_134;
  wire [13:0] T_1050;
  wire [12:0] T_1051;
  wire [12:0] T_1053;
  wire [13:0] GEN_135;
  wire [13:0] sExpX_E;
  wire [12:0] posExpX_E;
  wire [12:0] T_1054;
  wire [8192:0] GEN_136;
  wire [8192:0] T_1056;
  wire [52:0] T_1057;
  wire [31:0] T_1058;
  wire [15:0] T_1063;
  wire [31:0] GEN_137;
  wire [31:0] T_1064;
  wire [15:0] T_1065;
  wire [31:0] GEN_138;
  wire [31:0] T_1066;
  wire [31:0] T_1068;
  wire [31:0] T_1069;
  wire [23:0] T_1073;
  wire [31:0] GEN_139;
  wire [31:0] T_1074;
  wire [23:0] T_1075;
  wire [31:0] GEN_140;
  wire [31:0] T_1076;
  wire [31:0] T_1078;
  wire [31:0] T_1079;
  wire [27:0] T_1083;
  wire [31:0] GEN_141;
  wire [31:0] T_1084;
  wire [27:0] T_1085;
  wire [31:0] GEN_142;
  wire [31:0] T_1086;
  wire [31:0] T_1088;
  wire [31:0] T_1089;
  wire [29:0] T_1093;
  wire [31:0] GEN_143;
  wire [31:0] T_1094;
  wire [29:0] T_1095;
  wire [31:0] GEN_144;
  wire [31:0] T_1096;
  wire [31:0] T_1098;
  wire [31:0] T_1099;
  wire [30:0] T_1103;
  wire [31:0] GEN_145;
  wire [31:0] T_1104;
  wire [30:0] T_1105;
  wire [31:0] GEN_146;
  wire [31:0] T_1106;
  wire [31:0] T_1108;
  wire [31:0] T_1109;
  wire [20:0] T_1110;
  wire [15:0] T_1111;
  wire [7:0] T_1116;
  wire [15:0] GEN_147;
  wire [15:0] T_1117;
  wire [7:0] T_1118;
  wire [15:0] GEN_148;
  wire [15:0] T_1119;
  wire [15:0] T_1121;
  wire [15:0] T_1122;
  wire [11:0] T_1126;
  wire [15:0] GEN_149;
  wire [15:0] T_1127;
  wire [11:0] T_1128;
  wire [15:0] GEN_150;
  wire [15:0] T_1129;
  wire [15:0] T_1131;
  wire [15:0] T_1132;
  wire [13:0] T_1136;
  wire [15:0] GEN_151;
  wire [15:0] T_1137;
  wire [13:0] T_1138;
  wire [15:0] GEN_152;
  wire [15:0] T_1139;
  wire [15:0] T_1141;
  wire [15:0] T_1142;
  wire [14:0] T_1146;
  wire [15:0] GEN_153;
  wire [15:0] T_1147;
  wire [14:0] T_1148;
  wire [15:0] GEN_154;
  wire [15:0] T_1149;
  wire [15:0] T_1151;
  wire [15:0] T_1152;
  wire [4:0] T_1153;
  wire [3:0] T_1154;
  wire [1:0] T_1155;
  wire  T_1156;
  wire  T_1157;
  wire [1:0] T_1158;
  wire [1:0] T_1159;
  wire  T_1160;
  wire  T_1161;
  wire [1:0] T_1162;
  wire [3:0] T_1163;
  wire  T_1164;
  wire [4:0] T_1165;
  wire [20:0] T_1166;
  wire [52:0] roundMask_E;
  wire [53:0] T_1168;
  wire [53:0] T_1169;
  wire [53:0] T_1171;
  wire [53:0] incrPosMask_E;
  wire [52:0] T_1172;
  wire [52:0] T_1173;
  wire [52:0] GEN_155;
  wire  hiRoundPosBitT_E;
  wire [51:0] T_1175;
  wire [52:0] GEN_156;
  wire [52:0] T_1178;
  wire [52:0] T_1180;
  wire  all1sHiRoundExtraT_E;
  wire  T_1182;
  wire  T_1184;
  wire  T_1185;
  wire  all1sHiRoundT_E;
  wire [53:0] GEN_160;
  wire [54:0] T_1187;
  wire [53:0] T_1188;
  wire [53:0] GEN_161;
  wire [54:0] T_1189;
  wire [53:0] sigAdjT_E;
  wire [52:0] T_1191;
  wire [53:0] T_1192;
  wire [53:0] sigY0_E;
  wire [53:0] T_1195;
  wire [53:0] GEN_162;
  wire [54:0] T_1197;
  wire [53:0] sigY1_E;
  wire  T_1199;
  wire  T_1201;
  wire  T_1202;
  wire  trueLtX_E1;
  wire  T_1205;
  wire  T_1206;
  wire  T_1207;
  wire  T_1208;
  wire  hiRoundPosBit_E1;
  wire  T_1213;
  wire  T_1215;
  wire  anyRoundExtra_E1;
  wire  T_1216;
  wire  T_1218;
  wire  T_1219;
  wire [53:0] roundEvenMask_E1;
  wire  T_1221;
  wire  T_1224;
  wire  T_1225;
  wire  T_1228;
  wire  T_1231;
  wire  T_1233;
  wire  T_1234;
  wire  T_1235;
  wire  T_1236;
  wire  T_1239;
  wire  T_1243;
  wire  T_1244;
  wire  T_1248;
  wire  T_1249;
  wire  T_1250;
  wire  T_1251;
  wire [53:0] T_1252;
  wire [53:0] T_1253;
  wire [53:0] sigY_E1;
  wire [51:0] fractY_E1;
  wire  inexactY_E1;
  wire  T_1254;
  wire  T_1256;
  wire [13:0] T_1258;
  wire  T_1262;
  wire  T_1263;
  wire [13:0] T_1265;
  wire [13:0] T_1266;
  wire  T_1273;
  wire [13:0] T_1275;
  wire [13:0] T_1276;
  wire  T_1278;
  wire [12:0] T_1279;
  wire [13:0] T_1281;
  wire [12:0] T_1282;
  wire [12:0] T_1284;
  wire [13:0] GEN_164;
  wire [13:0] sExpY_E1;
  wire [11:0] expY_E1;
  wire  T_1285;
  wire  T_1287;
  wire [2:0] T_1289;
  wire  T_1290;
  wire  overflowY_E1;
  wire [12:0] T_1292;
  wire  T_1294;
  wire  totalUnderflowY_E1;
  wire  T_1296;
  wire  T_1297;
  wire  underflowY_E1;
  wire  T_1299;
  wire  T_1302;
  wire  T_1303;
  wire  T_1304;
  wire  T_1305;
  wire  T_1306;
  wire  notSigNaN_invalid_PC;
  wire  T_1309;
  wire  T_1310;
  wire  invalid_PC;
  wire  T_1315;
  wire  T_1318;
  wire  infinity_PC;
  wire  overflow_E1;
  wire  underflow_E1;
  wire  T_1319;
  wire  T_1320;
  wire  inexact_E1;
  wire  T_1321;
  wire  T_1324;
  wire  T_1325;
  wire  notSpecial_isZeroOut_E1;
  wire  T_1326;
  wire  pegMinFiniteMagOut_E1;
  wire  T_1328;
  wire  pegMaxFiniteMagOut_E1;
  wire  T_1329;
  wire  T_1330;
  wire  T_1331;
  wire  notNaN_isInfOut_E1;
  wire  T_1334;
  wire  T_1335;
  wire  isNaNOut_PC;
  wire  T_1337;
  wire  T_1338;
  wire  T_1339;
  wire  signOut_PC;
  wire [11:0] T_1343;
  wire [11:0] T_1344;
  wire [11:0] T_1345;
  wire [11:0] T_1349;
  wire [11:0] T_1350;
  wire [11:0] T_1351;
  wire [11:0] T_1355;
  wire [11:0] T_1356;
  wire [11:0] T_1357;
  wire [11:0] T_1361;
  wire [11:0] T_1362;
  wire [11:0] T_1363;
  wire [11:0] T_1366;
  wire [11:0] T_1367;
  wire [11:0] T_1370;
  wire [11:0] T_1371;
  wire [11:0] T_1374;
  wire [11:0] T_1375;
  wire [11:0] T_1378;
  wire [11:0] expOut_E1;
  wire  T_1379;
  wire  T_1380;
  wire [51:0] T_1384;
  wire [51:0] T_1385;
  wire [51:0] GEN_165;
  wire [52:0] T_1387;
  wire [51:0] T_1388;
  wire [51:0] fractOut_E1;
  wire [12:0] T_1389;
  wire [64:0] T_1390;
  wire [1:0] T_1391;
  wire [1:0] T_1392;
  wire [2:0] T_1393;
  wire [4:0] T_1394;
  assign io_inReady_div = T_138;
  assign io_inReady_sqrt = T_153;
  assign io_outValid_div = T_370;
  assign io_outValid_sqrt = T_371;
  assign io_out = T_1390;
  assign io_exceptionFlags = T_1394;
  assign io_usingMulAdd = T_951;
  assign io_latchMulAddA_0 = T_860;
  assign io_mulAddA_0 = T_890;
  assign io_latchMulAddB_0 = T_896;
  assign io_mulAddB_0 = T_916;
  assign io_mulAddC_2 = T_989;
  assign ready_PA = T_257;
  assign ready_PB = T_298;
  assign ready_PC = T_367;
  assign leaving_PA = T_254;
  assign leaving_PB = T_295;
  assign leaving_PC = T_364;
  assign cyc_B10_sqrt = T_413;
  assign cyc_B9_sqrt = T_415;
  assign cyc_B8_sqrt = T_417;
  assign cyc_B7_sqrt = T_419;
  assign cyc_B6 = T_421;
  assign cyc_B5 = T_423;
  assign cyc_B4 = T_425;
  assign cyc_B3 = T_427;
  assign cyc_B2 = T_429;
  assign cyc_B1 = T_431;
  assign cyc_B6_div = T_435;
  assign cyc_B5_div = T_439;
  assign cyc_B4_div = T_443;
  assign cyc_B3_div = T_446;
  assign cyc_B2_div = T_449;
  assign cyc_B1_div = T_452;
  assign cyc_B6_sqrt = T_454;
  assign cyc_B5_sqrt = T_456;
  assign cyc_B4_sqrt = T_458;
  assign cyc_B3_sqrt = T_459;
  assign cyc_B2_sqrt = T_460;
  assign cyc_B1_sqrt = T_461;
  assign cyc_C5 = T_474;
  assign cyc_C4 = T_476;
  assign valid_normalCase_leaving_PB = T_478;
  assign cyc_C2 = T_480;
  assign cyc_C1 = T_482;
  assign cyc_E4 = T_502;
  assign cyc_E3 = T_504;
  assign cyc_E2 = T_506;
  assign cyc_E1 = T_508;
  assign zSigma1_B4 = T_993;
  assign sigXNU_B3_CX = T_994;
  assign zComplSigT_C1_sqrt = T_1016;
  assign zComplSigT_C1 = T_1012;
  assign T_113 = cyc_B7_sqrt == 1'h0;
  assign T_114 = ready_PA & T_113;
  assign T_116 = cyc_B6_sqrt == 1'h0;
  assign T_117 = T_114 & T_116;
  assign T_119 = cyc_B5_sqrt == 1'h0;
  assign T_120 = T_117 & T_119;
  assign T_122 = cyc_B4_sqrt == 1'h0;
  assign T_123 = T_120 & T_122;
  assign T_125 = cyc_B3 == 1'h0;
  assign T_126 = T_123 & T_125;
  assign T_128 = cyc_B2 == 1'h0;
  assign T_129 = T_126 & T_128;
  assign T_131 = cyc_B1_sqrt == 1'h0;
  assign T_132 = T_129 & T_131;
  assign T_134 = cyc_C5 == 1'h0;
  assign T_135 = T_132 & T_134;
  assign T_137 = cyc_C4 == 1'h0;
  assign T_138 = T_135 & T_137;
  assign T_141 = ready_PA & T_116;
  assign T_144 = T_141 & T_119;
  assign T_147 = T_144 & T_122;
  assign T_149 = cyc_B2_div == 1'h0;
  assign T_150 = T_147 & T_149;
  assign T_153 = T_150 & T_131;
  assign T_154 = io_inReady_div & io_inValid;
  assign T_156 = io_sqrtOp == 1'h0;
  assign cyc_S_div = T_154 & T_156;
  assign T_157 = io_inReady_sqrt & io_inValid;
  assign cyc_S_sqrt = T_157 & io_sqrtOp;
  assign cyc_S = cyc_S_div | cyc_S_sqrt;
  assign signA_S = io_a[64];
  assign expA_S = io_a[63:52];
  assign fractA_S = io_a[51:0];
  assign specialCodeA_S = expA_S[11:9];
  assign isZeroA_S = specialCodeA_S == 3'h0;
  assign T_159 = specialCodeA_S[2:1];
  assign isSpecialA_S = T_159 == 2'h3;
  assign signB_S = io_b[64];
  assign expB_S = io_b[63:52];
  assign fractB_S = io_b[51:0];
  assign specialCodeB_S = expB_S[11:9];
  assign isZeroB_S = specialCodeB_S == 3'h0;
  assign T_162 = specialCodeB_S[2:1];
  assign isSpecialB_S = T_162 == 2'h3;
  assign T_164 = signA_S ^ signB_S;
  assign sign_S = io_sqrtOp ? signB_S : T_164;
  assign T_166 = isSpecialA_S == 1'h0;
  assign T_168 = isSpecialB_S == 1'h0;
  assign T_169 = T_166 & T_168;
  assign T_171 = isZeroA_S == 1'h0;
  assign T_172 = T_169 & T_171;
  assign T_174 = isZeroB_S == 1'h0;
  assign normalCase_S_div = T_172 & T_174;
  assign T_179 = T_168 & T_174;
  assign T_181 = signB_S == 1'h0;
  assign normalCase_S_sqrt = T_179 & T_181;
  assign normalCase_S = io_sqrtOp ? normalCase_S_sqrt : normalCase_S_div;
  assign entering_PA_normalCase_div = cyc_S_div & normalCase_S_div;
  assign entering_PA_normalCase_sqrt = cyc_S_sqrt & normalCase_S_sqrt;
  assign entering_PA_normalCase = entering_PA_normalCase_div | entering_PA_normalCase_sqrt;
  assign T_183 = ready_PB == 1'h0;
  assign T_184 = valid_PA | T_183;
  assign T_185 = cyc_S & T_184;
  assign entering_PA = entering_PA_normalCase | T_185;
  assign T_187 = normalCase_S == 1'h0;
  assign T_188 = cyc_S & T_187;
  assign T_190 = valid_PA == 1'h0;
  assign T_191 = T_188 & T_190;
  assign T_193 = valid_PB == 1'h0;
  assign T_195 = ready_PC == 1'h0;
  assign T_196 = T_193 & T_195;
  assign T_197 = leaving_PB | T_196;
  assign entering_PB_S = T_191 & T_197;
  assign T_206 = T_191 & T_193;
  assign entering_PC_S = T_206 & ready_PC;
  assign T_207 = entering_PA | leaving_PA;
  assign GEN_0 = T_207 ? entering_PA : valid_PA;
  assign T_208 = fractB_S[51];
  assign GEN_1 = entering_PA ? io_sqrtOp : sqrtOp_PA;
  assign GEN_2 = entering_PA ? sign_S : sign_PA;
  assign GEN_3 = entering_PA ? specialCodeB_S : specialCodeB_PA;
  assign GEN_4 = entering_PA ? T_208 : fractB_51_PA;
  assign GEN_5 = entering_PA ? io_roundingMode : roundingMode_PA;
  assign T_211 = entering_PA & T_156;
  assign T_212 = fractA_S[51];
  assign GEN_6 = T_211 ? specialCodeA_S : specialCodeA_PA;
  assign GEN_7 = T_211 ? T_212 : fractA_51_PA;
  assign T_213 = expB_S[11];
  assign GEN_53 = {{2'd0}, T_213};
  assign T_215 = 3'h0 - GEN_53;
  assign T_216 = T_215[2:0];
  assign T_217 = expB_S[10:0];
  assign T_218 = ~ T_217;
  assign T_219 = {T_216,T_218};
  assign GEN_54 = {{2'd0}, expA_S};
  assign T_220 = GEN_54 + T_219;
  assign T_221 = T_220[13:0];
  assign T_222 = io_sqrtOp ? {{2'd0}, expB_S} : T_221;
  assign T_223 = fractB_S[50:0];
  assign GEN_8 = entering_PA_normalCase ? T_222 : exp_PA;
  assign GEN_9 = entering_PA_normalCase ? T_223 : fractB_other_PA;
  assign T_224 = fractA_S[50:0];
  assign GEN_10 = entering_PA_normalCase_div ? T_224 : fractA_other_PA;
  assign isZeroA_PA = specialCodeA_PA == 3'h0;
  assign T_226 = specialCodeA_PA[2:1];
  assign isSpecialA_PA = T_226 == 2'h3;
  assign T_229 = {1'h1,fractA_51_PA};
  assign sigA_PA = {T_229,fractA_other_PA};
  assign isZeroB_PA = specialCodeB_PA == 3'h0;
  assign T_231 = specialCodeB_PA[2:1];
  assign isSpecialB_PA = T_231 == 2'h3;
  assign T_234 = {1'h1,fractB_51_PA};
  assign sigB_PA = {T_234,fractB_other_PA};
  assign T_236 = isSpecialB_PA == 1'h0;
  assign T_238 = isZeroB_PA == 1'h0;
  assign T_239 = T_236 & T_238;
  assign T_241 = sign_PA == 1'h0;
  assign T_242 = T_239 & T_241;
  assign T_244 = isSpecialA_PA == 1'h0;
  assign T_247 = T_244 & T_236;
  assign T_249 = isZeroA_PA == 1'h0;
  assign T_250 = T_247 & T_249;
  assign T_253 = T_250 & T_238;
  assign normalCase_PA = sqrtOp_PA ? T_242 : T_253;
  assign valid_normalCase_leaving_PA = cyc_B4_div | cyc_B7_sqrt;
  assign valid_leaving_PA = normalCase_PA ? valid_normalCase_leaving_PA : ready_PB;
  assign T_254 = valid_PA & valid_leaving_PA;
  assign T_257 = T_190 | valid_leaving_PA;
  assign T_258 = valid_PA & normalCase_PA;
  assign entering_PB_normalCase = T_258 & valid_normalCase_leaving_PA;
  assign entering_PB = entering_PB_S | leaving_PA;
  assign T_259 = entering_PB | leaving_PB;
  assign GEN_11 = T_259 ? entering_PB : valid_PB;
  assign T_260 = valid_PA ? sqrtOp_PA : io_sqrtOp;
  assign T_261 = valid_PA ? sign_PA : sign_S;
  assign T_262 = valid_PA ? specialCodeA_PA : specialCodeA_S;
  assign T_264 = valid_PA ? fractA_51_PA : T_212;
  assign T_265 = valid_PA ? specialCodeB_PA : specialCodeB_S;
  assign T_267 = valid_PA ? fractB_51_PA : T_208;
  assign T_268 = valid_PA ? roundingMode_PA : io_roundingMode;
  assign GEN_12 = entering_PB ? T_260 : sqrtOp_PB;
  assign GEN_13 = entering_PB ? T_261 : sign_PB;
  assign GEN_14 = entering_PB ? T_262 : specialCodeA_PB;
  assign GEN_15 = entering_PB ? T_264 : fractA_51_PB;
  assign GEN_16 = entering_PB ? T_265 : specialCodeB_PB;
  assign GEN_17 = entering_PB ? T_267 : fractB_51_PB;
  assign GEN_18 = entering_PB ? T_268 : roundingMode_PB;
  assign T_269 = fractA_other_PA[0];
  assign GEN_19 = entering_PB_normalCase ? exp_PA : exp_PB;
  assign GEN_20 = entering_PB_normalCase ? T_269 : fractA_0_PB;
  assign GEN_21 = entering_PB_normalCase ? fractB_other_PA : fractB_other_PB;
  assign isZeroA_PB = specialCodeA_PB == 3'h0;
  assign T_271 = specialCodeA_PB[2:1];
  assign isSpecialA_PB = T_271 == 2'h3;
  assign isZeroB_PB = specialCodeB_PB == 3'h0;
  assign T_274 = specialCodeB_PB[2:1];
  assign isSpecialB_PB = T_274 == 2'h3;
  assign T_277 = isSpecialB_PB == 1'h0;
  assign T_279 = isZeroB_PB == 1'h0;
  assign T_280 = T_277 & T_279;
  assign T_282 = sign_PB == 1'h0;
  assign T_283 = T_280 & T_282;
  assign T_285 = isSpecialA_PB == 1'h0;
  assign T_288 = T_285 & T_277;
  assign T_290 = isZeroA_PB == 1'h0;
  assign T_291 = T_288 & T_290;
  assign T_294 = T_291 & T_279;
  assign normalCase_PB = sqrtOp_PB ? T_283 : T_294;
  assign valid_leaving_PB = normalCase_PB ? valid_normalCase_leaving_PB : ready_PC;
  assign T_295 = valid_PB & valid_leaving_PB;
  assign T_298 = T_193 | valid_leaving_PB;
  assign T_299 = valid_PB & normalCase_PB;
  assign entering_PC_normalCase = T_299 & valid_normalCase_leaving_PB;
  assign entering_PC = entering_PC_S | leaving_PB;
  assign T_300 = entering_PC | leaving_PC;
  assign GEN_22 = T_300 ? entering_PC : valid_PC;
  assign T_301 = valid_PB ? sqrtOp_PB : io_sqrtOp;
  assign T_302 = valid_PB ? sign_PB : sign_S;
  assign T_303 = valid_PB ? specialCodeA_PB : specialCodeA_S;
  assign T_305 = valid_PB ? fractA_51_PB : T_212;
  assign T_306 = valid_PB ? specialCodeB_PB : specialCodeB_S;
  assign T_308 = valid_PB ? fractB_51_PB : T_208;
  assign T_309 = valid_PB ? roundingMode_PB : io_roundingMode;
  assign GEN_23 = entering_PC ? T_301 : sqrtOp_PC;
  assign GEN_24 = entering_PC ? T_302 : sign_PC;
  assign GEN_25 = entering_PC ? T_303 : specialCodeA_PC;
  assign GEN_26 = entering_PC ? T_305 : fractA_51_PC;
  assign GEN_27 = entering_PC ? T_306 : specialCodeB_PC;
  assign GEN_28 = entering_PC ? T_308 : fractB_51_PC;
  assign GEN_29 = entering_PC ? T_309 : roundingMode_PC;
  assign GEN_30 = entering_PC_normalCase ? exp_PB : exp_PC;
  assign GEN_31 = entering_PC_normalCase ? fractA_0_PB : fractA_0_PC;
  assign GEN_32 = entering_PC_normalCase ? fractB_other_PB : fractB_other_PC;
  assign isZeroA_PC = specialCodeA_PC == 3'h0;
  assign T_311 = specialCodeA_PC[2:1];
  assign isSpecialA_PC = T_311 == 2'h3;
  assign T_313 = specialCodeA_PC[0];
  assign T_315 = T_313 == 1'h0;
  assign isInfA_PC = isSpecialA_PC & T_315;
  assign isNaNA_PC = isSpecialA_PC & T_313;
  assign T_318 = fractA_51_PC == 1'h0;
  assign isSigNaNA_PC = isNaNA_PC & T_318;
  assign isZeroB_PC = specialCodeB_PC == 3'h0;
  assign T_320 = specialCodeB_PC[2:1];
  assign isSpecialB_PC = T_320 == 2'h3;
  assign T_322 = specialCodeB_PC[0];
  assign T_324 = T_322 == 1'h0;
  assign isInfB_PC = isSpecialB_PC & T_324;
  assign isNaNB_PC = isSpecialB_PC & T_322;
  assign T_327 = fractB_51_PC == 1'h0;
  assign isSigNaNB_PC = isNaNB_PC & T_327;
  assign T_329 = {1'h1,fractB_51_PC};
  assign sigB_PC = {T_329,fractB_other_PC};
  assign T_331 = isSpecialB_PC == 1'h0;
  assign T_333 = isZeroB_PC == 1'h0;
  assign T_334 = T_331 & T_333;
  assign T_336 = sign_PC == 1'h0;
  assign T_337 = T_334 & T_336;
  assign T_339 = isSpecialA_PC == 1'h0;
  assign T_342 = T_339 & T_331;
  assign T_344 = isZeroA_PC == 1'h0;
  assign T_345 = T_342 & T_344;
  assign T_348 = T_345 & T_333;
  assign normalCase_PC = sqrtOp_PC ? T_337 : T_348;
  assign GEN_55 = {{12'd0}, 2'h2};
  assign T_350 = exp_PC + GEN_55;
  assign expP2_PC = T_350[13:0];
  assign T_351 = exp_PC[0];
  assign T_352 = expP2_PC[13:1];
  assign T_354 = {T_352,1'h0};
  assign T_355 = exp_PC[13:1];
  assign T_357 = {T_355,1'h1};
  assign expP1_PC = T_351 ? T_354 : T_357;
  assign roundingMode_near_even_PC = roundingMode_PC == 2'h0;
  assign roundingMode_min_PC = roundingMode_PC == 2'h2;
  assign roundingMode_max_PC = roundingMode_PC == 2'h3;
  assign roundMagUp_PC = sign_PC ? roundingMode_min_PC : roundingMode_max_PC;
  assign overflowY_roundMagUp_PC = roundingMode_near_even_PC | roundMagUp_PC;
  assign T_359 = roundMagUp_PC == 1'h0;
  assign T_361 = roundingMode_near_even_PC == 1'h0;
  assign roundMagDown_PC = T_359 & T_361;
  assign T_363 = normalCase_PC == 1'h0;
  assign valid_leaving_PC = T_363 | cyc_E1;
  assign T_364 = valid_PC & valid_leaving_PC;
  assign T_366 = valid_PC == 1'h0;
  assign T_367 = T_366 | valid_leaving_PC;
  assign T_369 = sqrtOp_PC == 1'h0;
  assign T_370 = leaving_PC & T_369;
  assign T_371 = leaving_PC & sqrtOp_PC;
  assign GEN_56 = {{2'd0}, 1'h0};
  assign T_373 = cycleNum_A != GEN_56;
  assign T_374 = entering_PA_normalCase | T_373;
  assign T_377 = entering_PA_normalCase_div ? 2'h3 : {{1'd0}, 1'h0};
  assign T_380 = entering_PA_normalCase_sqrt ? 3'h6 : {{2'd0}, 1'h0};
  assign GEN_57 = {{1'd0}, T_377};
  assign T_381 = GEN_57 | T_380;
  assign T_383 = entering_PA_normalCase == 1'h0;
  assign GEN_58 = {{2'd0}, 1'h1};
  assign T_385 = cycleNum_A - GEN_58;
  assign T_386 = T_385[2:0];
  assign T_388 = T_383 ? T_386 : {{2'd0}, 1'h0};
  assign T_389 = T_381 | T_388;
  assign GEN_33 = T_374 ? T_389 : cycleNum_A;
  assign cyc_A6_sqrt = cycleNum_A == 3'h6;
  assign cyc_A5_sqrt = cycleNum_A == 3'h5;
  assign cyc_A4_sqrt = cycleNum_A == 3'h4;
  assign cyc_A4 = cyc_A4_sqrt | entering_PA_normalCase_div;
  assign GEN_59 = {{1'd0}, 2'h3};
  assign cyc_A3 = cycleNum_A == GEN_59;
  assign GEN_60 = {{1'd0}, 2'h2};
  assign cyc_A2 = cycleNum_A == GEN_60;
  assign cyc_A1 = cycleNum_A == GEN_58;
  assign T_397 = sqrtOp_PA == 1'h0;
  assign cyc_A3_div = cyc_A3 & T_397;
  assign cyc_A2_div = cyc_A2 & T_397;
  assign cyc_A1_div = cyc_A1 & T_397;
  assign cyc_A3_sqrt = cyc_A3 & sqrtOp_PA;
  assign cyc_A1_sqrt = cyc_A1 & sqrtOp_PA;
  assign GEN_62 = {{3'd0}, 1'h0};
  assign T_403 = cycleNum_B != GEN_62;
  assign T_404 = cyc_A1 | T_403;
  assign T_407 = sqrtOp_PA ? 4'ha : {{1'd0}, 3'h6};
  assign GEN_63 = {{3'd0}, 1'h1};
  assign T_409 = cycleNum_B - GEN_63;
  assign T_410 = T_409[3:0];
  assign T_411 = cyc_A1 ? T_407 : T_410;
  assign GEN_34 = T_404 ? T_411 : cycleNum_B;
  assign T_413 = cycleNum_B == 4'ha;
  assign T_415 = cycleNum_B == 4'h9;
  assign T_417 = cycleNum_B == 4'h8;
  assign GEN_64 = {{1'd0}, 3'h7};
  assign T_419 = cycleNum_B == GEN_64;
  assign GEN_65 = {{1'd0}, 3'h6};
  assign T_421 = cycleNum_B == GEN_65;
  assign GEN_66 = {{1'd0}, 3'h5};
  assign T_423 = cycleNum_B == GEN_66;
  assign GEN_67 = {{1'd0}, 3'h4};
  assign T_425 = cycleNum_B == GEN_67;
  assign GEN_68 = {{2'd0}, 2'h3};
  assign T_427 = cycleNum_B == GEN_68;
  assign GEN_69 = {{2'd0}, 2'h2};
  assign T_429 = cycleNum_B == GEN_69;
  assign T_431 = cycleNum_B == GEN_63;
  assign T_432 = cyc_B6 & valid_PA;
  assign T_435 = T_432 & T_397;
  assign T_436 = cyc_B5 & valid_PA;
  assign T_439 = T_436 & T_397;
  assign T_440 = cyc_B4 & valid_PA;
  assign T_443 = T_440 & T_397;
  assign T_445 = sqrtOp_PB == 1'h0;
  assign T_446 = cyc_B3 & T_445;
  assign T_449 = cyc_B2 & T_445;
  assign T_452 = cyc_B1 & T_445;
  assign T_453 = cyc_B6 & valid_PB;
  assign T_454 = T_453 & sqrtOp_PB;
  assign T_455 = cyc_B5 & valid_PB;
  assign T_456 = T_455 & sqrtOp_PB;
  assign T_457 = cyc_B4 & valid_PB;
  assign T_458 = T_457 & sqrtOp_PB;
  assign T_459 = cyc_B3 & sqrtOp_PB;
  assign T_460 = cyc_B2 & sqrtOp_PB;
  assign T_461 = cyc_B1 & sqrtOp_PB;
  assign T_463 = cycleNum_C != GEN_56;
  assign T_464 = cyc_B1 | T_463;
  assign T_467 = sqrtOp_PB ? 3'h6 : 3'h5;
  assign T_469 = cycleNum_C - GEN_58;
  assign T_470 = T_469[2:0];
  assign T_471 = cyc_B1 ? T_467 : T_470;
  assign GEN_35 = T_464 ? T_471 : cycleNum_C;
  assign cyc_C6_sqrt = cycleNum_C == 3'h6;
  assign T_474 = cycleNum_C == 3'h5;
  assign T_476 = cycleNum_C == 3'h4;
  assign T_478 = cycleNum_C == GEN_59;
  assign T_480 = cycleNum_C == GEN_60;
  assign T_482 = cycleNum_C == GEN_58;
  assign cyc_C5_div = cyc_C5 & T_445;
  assign cyc_C4_div = cyc_C4 & T_445;
  assign cyc_C1_div = cyc_C1 & T_369;
  assign cyc_C5_sqrt = cyc_C5 & sqrtOp_PB;
  assign cyc_C4_sqrt = cyc_C4 & sqrtOp_PB;
  assign cyc_C3_sqrt = valid_normalCase_leaving_PB & sqrtOp_PB;
  assign cyc_C1_sqrt = cyc_C1 & sqrtOp_PC;
  assign T_494 = cycleNum_E != GEN_56;
  assign T_495 = cyc_C1 | T_494;
  assign T_498 = cycleNum_E - GEN_58;
  assign T_499 = T_498[2:0];
  assign T_500 = cyc_C1 ? 3'h4 : T_499;
  assign GEN_36 = T_495 ? T_500 : cycleNum_E;
  assign T_502 = cycleNum_E == 3'h4;
  assign T_504 = cycleNum_E == GEN_59;
  assign T_506 = cycleNum_E == GEN_60;
  assign T_508 = cycleNum_E == GEN_58;
  assign cyc_E3_div = cyc_E3 & T_369;
  assign cyc_E3_sqrt = cyc_E3 & sqrtOp_PC;
  assign zFractB_A4_div = entering_PA_normalCase_div ? fractB_S : {{51'd0}, 1'h0};
  assign T_518 = fractB_S[51:49];
  assign T_520 = T_518 == GEN_56;
  assign zLinPiece_0_A4_div = entering_PA_normalCase_div & T_520;
  assign T_523 = T_518 == GEN_58;
  assign zLinPiece_1_A4_div = entering_PA_normalCase_div & T_523;
  assign T_526 = T_518 == GEN_60;
  assign zLinPiece_2_A4_div = entering_PA_normalCase_div & T_526;
  assign T_529 = T_518 == GEN_59;
  assign zLinPiece_3_A4_div = entering_PA_normalCase_div & T_529;
  assign T_532 = T_518 == 3'h4;
  assign zLinPiece_4_A4_div = entering_PA_normalCase_div & T_532;
  assign T_535 = T_518 == 3'h5;
  assign zLinPiece_5_A4_div = entering_PA_normalCase_div & T_535;
  assign T_538 = T_518 == 3'h6;
  assign zLinPiece_6_A4_div = entering_PA_normalCase_div & T_538;
  assign T_541 = T_518 == 3'h7;
  assign zLinPiece_7_A4_div = entering_PA_normalCase_div & T_541;
  assign T_544 = zLinPiece_0_A4_div ? 9'h1c7 : {{8'd0}, 1'h0};
  assign T_547 = zLinPiece_1_A4_div ? 9'h16c : {{8'd0}, 1'h0};
  assign T_548 = T_544 | T_547;
  assign T_551 = zLinPiece_2_A4_div ? 9'h12a : {{8'd0}, 1'h0};
  assign T_552 = T_548 | T_551;
  assign T_555 = zLinPiece_3_A4_div ? 9'hf8 : {{8'd0}, 1'h0};
  assign T_556 = T_552 | T_555;
  assign T_559 = zLinPiece_4_A4_div ? 9'hd2 : {{8'd0}, 1'h0};
  assign T_560 = T_556 | T_559;
  assign T_563 = zLinPiece_5_A4_div ? 9'hb4 : {{8'd0}, 1'h0};
  assign T_564 = T_560 | T_563;
  assign T_567 = zLinPiece_6_A4_div ? 9'h9c : {{8'd0}, 1'h0};
  assign T_568 = T_564 | T_567;
  assign T_571 = zLinPiece_7_A4_div ? 9'h89 : {{8'd0}, 1'h0};
  assign zK1_A4_div = T_568 | T_571;
  assign T_575 = zLinPiece_0_A4_div ? 12'h1c : {{11'd0}, 1'h0};
  assign T_579 = zLinPiece_1_A4_div ? 12'h3a2 : {{11'd0}, 1'h0};
  assign T_580 = T_575 | T_579;
  assign T_584 = zLinPiece_2_A4_div ? 12'h675 : {{11'd0}, 1'h0};
  assign T_585 = T_580 | T_584;
  assign T_589 = zLinPiece_3_A4_div ? 12'h8c6 : {{11'd0}, 1'h0};
  assign T_590 = T_585 | T_589;
  assign T_594 = zLinPiece_4_A4_div ? 12'hab4 : {{11'd0}, 1'h0};
  assign T_595 = T_590 | T_594;
  assign T_599 = zLinPiece_5_A4_div ? 12'hc56 : {{11'd0}, 1'h0};
  assign T_600 = T_595 | T_599;
  assign T_604 = zLinPiece_6_A4_div ? 12'hdbd : {{11'd0}, 1'h0};
  assign T_605 = T_600 | T_604;
  assign T_609 = zLinPiece_7_A4_div ? 12'hef4 : {{11'd0}, 1'h0};
  assign zComplFractK0_A4_div = T_605 | T_609;
  assign zFractB_A7_sqrt = entering_PA_normalCase_sqrt ? fractB_S : {{51'd0}, 1'h0};
  assign T_611 = expB_S[0];
  assign T_613 = T_611 == 1'h0;
  assign T_614 = entering_PA_normalCase_sqrt & T_613;
  assign T_617 = T_208 == 1'h0;
  assign zQuadPiece_0_A7_sqrt = T_614 & T_617;
  assign zQuadPiece_1_A7_sqrt = T_614 & T_208;
  assign T_624 = entering_PA_normalCase_sqrt & T_611;
  assign zQuadPiece_2_A7_sqrt = T_624 & T_617;
  assign zQuadPiece_3_A7_sqrt = T_624 & T_208;
  assign T_633 = zQuadPiece_0_A7_sqrt ? 9'h1c8 : {{8'd0}, 1'h0};
  assign T_636 = zQuadPiece_1_A7_sqrt ? 9'hc1 : {{8'd0}, 1'h0};
  assign T_637 = T_633 | T_636;
  assign T_640 = zQuadPiece_2_A7_sqrt ? 9'h143 : {{8'd0}, 1'h0};
  assign T_641 = T_637 | T_640;
  assign T_644 = zQuadPiece_3_A7_sqrt ? 9'h89 : {{8'd0}, 1'h0};
  assign zK2_A7_sqrt = T_641 | T_644;
  assign T_648 = zQuadPiece_0_A7_sqrt ? 10'h2f : {{9'd0}, 1'h0};
  assign T_652 = zQuadPiece_1_A7_sqrt ? 10'h1df : {{9'd0}, 1'h0};
  assign T_653 = T_648 | T_652;
  assign T_657 = zQuadPiece_2_A7_sqrt ? 10'h14d : {{9'd0}, 1'h0};
  assign T_658 = T_653 | T_657;
  assign T_662 = zQuadPiece_3_A7_sqrt ? 10'h27e : {{9'd0}, 1'h0};
  assign zComplK1_A7_sqrt = T_658 | T_662;
  assign T_663 = exp_PA[0];
  assign T_665 = T_663 == 1'h0;
  assign T_666 = cyc_A6_sqrt & T_665;
  assign T_667 = sigB_PA[51];
  assign T_669 = T_667 == 1'h0;
  assign zQuadPiece_0_A6_sqrt = T_666 & T_669;
  assign zQuadPiece_1_A6_sqrt = T_666 & T_667;
  assign T_676 = cyc_A6_sqrt & T_663;
  assign zQuadPiece_2_A6_sqrt = T_676 & T_669;
  assign zQuadPiece_3_A6_sqrt = T_676 & T_667;
  assign T_686 = zQuadPiece_0_A6_sqrt ? 13'h1a : {{12'd0}, 1'h0};
  assign T_690 = zQuadPiece_1_A6_sqrt ? 13'hbca : {{12'd0}, 1'h0};
  assign T_691 = T_686 | T_690;
  assign T_695 = zQuadPiece_2_A6_sqrt ? 13'h12d3 : {{12'd0}, 1'h0};
  assign T_696 = T_691 | T_695;
  assign T_700 = zQuadPiece_3_A6_sqrt ? 13'h1b17 : {{12'd0}, 1'h0};
  assign zComplFractK0_A6_sqrt = T_696 | T_700;
  assign T_701 = zFractB_A4_div[48:40];
  assign T_702 = T_701 | zK2_A7_sqrt;
  assign T_704 = cyc_S == 1'h0;
  assign T_706 = T_704 ? nextMulAdd9A_A : {{8'd0}, 1'h0};
  assign mulAdd9A_A = T_702 | T_706;
  assign T_707 = zFractB_A7_sqrt[50:42];
  assign T_708 = zK1_A4_div | T_707;
  assign T_712 = T_704 ? nextMulAdd9B_A : {{8'd0}, 1'h0};
  assign mulAdd9B_A = T_708 | T_712;
  assign GEN_85 = {{9'd0}, entering_PA_normalCase_sqrt};
  assign T_714 = 10'h0 - GEN_85;
  assign T_715 = T_714[9:0];
  assign T_716 = {zComplK1_A7_sqrt,T_715};
  assign GEN_86 = {{5'd0}, cyc_A6_sqrt};
  assign T_718 = 6'h0 - GEN_86;
  assign T_719 = T_718[5:0];
  assign T_720 = {cyc_A6_sqrt,zComplFractK0_A6_sqrt};
  assign T_721 = {T_720,T_719};
  assign T_722 = T_716 | T_721;
  assign GEN_87 = {{7'd0}, entering_PA_normalCase_div};
  assign T_724 = 8'h0 - GEN_87;
  assign T_725 = T_724[7:0];
  assign T_726 = {entering_PA_normalCase_div,zComplFractK0_A4_div};
  assign T_727 = {T_726,T_725};
  assign GEN_88 = {{1'd0}, T_722};
  assign T_728 = GEN_88 | T_727;
  assign GEN_89 = {{10'd0}, fractR0_A};
  assign T_730 = GEN_89 << 10;
  assign GEN_90 = {{1'd0}, T_730};
  assign T_731 = 20'h40000 + GEN_90;
  assign T_732 = T_731[19:0];
  assign T_734 = cyc_A5_sqrt ? T_732 : {{19'd0}, 1'h0};
  assign GEN_91 = {{1'd0}, T_734};
  assign T_735 = T_728 | GEN_91;
  assign T_736 = hiSqrR0_A_sqrt[9];
  assign T_738 = T_736 == 1'h0;
  assign T_739 = cyc_A4_sqrt & T_738;
  assign T_742 = T_739 ? 11'h400 : {{10'd0}, 1'h0};
  assign GEN_92 = {{10'd0}, T_742};
  assign T_743 = T_735 | GEN_92;
  assign T_745 = cyc_A4_sqrt & T_736;
  assign T_746 = T_745 | cyc_A3_div;
  assign T_747 = sigB_PA[46:26];
  assign GEN_93 = {{10'd0}, 11'h400};
  assign T_749 = T_747 + GEN_93;
  assign T_750 = T_749[20:0];
  assign T_752 = T_746 ? T_750 : {{20'd0}, 1'h0};
  assign T_753 = T_743 | T_752;
  assign T_754 = cyc_A3_sqrt | cyc_A2;
  assign T_756 = T_754 ? partNegSigma0_A : {{20'd0}, 1'h0};
  assign T_757 = T_753 | T_756;
  assign GEN_94 = {{16'd0}, fractR0_A};
  assign T_758 = GEN_94 << 16;
  assign T_760 = cyc_A1_sqrt ? T_758 : {{24'd0}, 1'h0};
  assign GEN_95 = {{4'd0}, T_757};
  assign T_761 = GEN_95 | T_760;
  assign GEN_96 = {{15'd0}, fractR0_A};
  assign T_762 = GEN_96 << 15;
  assign T_764 = cyc_A1_div ? T_762 : {{23'd0}, 1'h0};
  assign GEN_97 = {{1'd0}, T_764};
  assign mulAdd9C_A = T_761 | GEN_97;
  assign T_765 = mulAdd9A_A * mulAdd9B_A;
  assign T_767 = mulAdd9C_A[17:0];
  assign T_768 = {1'h0,T_767};
  assign GEN_98 = {{1'd0}, T_765};
  assign T_769 = GEN_98 + T_768;
  assign loMulAdd9Out_A = T_769[18:0];
  assign T_770 = loMulAdd9Out_A[18];
  assign T_771 = mulAdd9C_A[24:18];
  assign GEN_99 = {{6'd0}, 1'h1};
  assign T_773 = T_771 + GEN_99;
  assign T_774 = T_773[6:0];
  assign T_776 = T_770 ? T_774 : T_771;
  assign T_777 = loMulAdd9Out_A[17:0];
  assign mulAdd9Out_A = {T_776,T_777};
  assign T_778 = mulAdd9Out_A[19];
  assign T_779 = cyc_A6_sqrt & T_778;
  assign T_780 = ~ mulAdd9Out_A;
  assign T_781 = T_780[24:10];
  assign T_783 = T_779 ? T_781 : {{14'd0}, 1'h0};
  assign zFractR0_A6_sqrt = T_783[8:0];
  assign GEN_100 = {{1'd0}, mulAdd9Out_A};
  assign T_785 = GEN_100 << 1;
  assign sqrR0_A5_sqrt = T_663 ? T_785 : {{1'd0}, mulAdd9Out_A};
  assign T_786 = mulAdd9Out_A[20];
  assign T_787 = entering_PA_normalCase_div & T_786;
  assign T_789 = T_780[24:11];
  assign T_791 = T_787 ? T_789 : {{13'd0}, 1'h0};
  assign zFractR0_A4_div = T_791[8:0];
  assign T_792 = mulAdd9Out_A[11];
  assign T_793 = cyc_A2 & T_792;
  assign T_795 = T_780[24:2];
  assign T_797 = T_793 ? T_795 : {{22'd0}, 1'h0};
  assign zSigma0_A2 = T_797[8:0];
  assign T_798 = mulAdd9Out_A[24:10];
  assign T_799 = mulAdd9Out_A[24:9];
  assign T_800 = sqrtOp_PA ? {{1'd0}, T_798} : T_799;
  assign fractR1_A1 = T_800[14:0];
  assign r1_A1 = {1'h1,fractR1_A1};
  assign GEN_101 = {{1'd0}, r1_A1};
  assign T_803 = GEN_101 << 1;
  assign ER1_A1_sqrt = T_663 ? T_803 : {{1'd0}, r1_A1};
  assign T_804 = cyc_A6_sqrt | entering_PA_normalCase_div;
  assign T_805 = zFractR0_A6_sqrt | zFractR0_A4_div;
  assign GEN_37 = T_804 ? T_805 : fractR0_A;
  assign T_806 = sqrR0_A5_sqrt[25:10];
  assign GEN_38 = cyc_A5_sqrt ? T_806 : {{6'd0}, hiSqrR0_A_sqrt};
  assign T_807 = cyc_A4_sqrt | cyc_A3;
  assign T_809 = cyc_A4_sqrt ? mulAdd9Out_A : {{9'd0}, T_799};
  assign T_810 = T_809[20:0];
  assign GEN_39 = T_807 ? T_810 : partNegSigma0_A;
  assign T_811 = entering_PA_normalCase_sqrt | cyc_A6_sqrt;
  assign T_812 = T_811 | cyc_A5_sqrt;
  assign T_813 = T_812 | cyc_A4;
  assign T_814 = T_813 | cyc_A3;
  assign T_815 = T_814 | cyc_A2;
  assign T_819 = entering_PA_normalCase_sqrt ? T_789 : {{13'd0}, 1'h0};
  assign GEN_102 = {{5'd0}, zFractR0_A6_sqrt};
  assign T_820 = T_819 | GEN_102;
  assign T_821 = sigB_PA[43:35];
  assign T_823 = cyc_A4_sqrt ? T_821 : {{8'd0}, 1'h0};
  assign GEN_103 = {{5'd0}, T_823};
  assign T_824 = T_820 | GEN_103;
  assign T_825 = zFractB_A4_div[43:35];
  assign GEN_104 = {{5'd0}, T_825};
  assign T_826 = T_824 | GEN_104;
  assign T_827 = cyc_A5_sqrt | cyc_A3;
  assign T_828 = sigB_PA[52:44];
  assign T_830 = T_827 ? T_828 : {{8'd0}, 1'h0};
  assign GEN_105 = {{5'd0}, T_830};
  assign T_831 = T_826 | GEN_105;
  assign GEN_106 = {{5'd0}, zSigma0_A2};
  assign T_832 = T_831 | GEN_106;
  assign GEN_40 = T_815 ? T_832 : {{5'd0}, nextMulAdd9A_A};
  assign T_836 = T_813 | cyc_A2;
  assign T_838 = T_707 | zFractR0_A6_sqrt;
  assign T_839 = sqrR0_A5_sqrt[9:1];
  assign T_841 = cyc_A5_sqrt ? T_839 : {{8'd0}, 1'h0};
  assign T_842 = T_838 | T_841;
  assign T_843 = T_842 | zFractR0_A4_div;
  assign T_844 = hiSqrR0_A_sqrt[8:0];
  assign T_846 = cyc_A4_sqrt ? T_844 : {{8'd0}, 1'h0};
  assign T_847 = T_843 | T_846;
  assign T_849 = fractR0_A[8:1];
  assign T_850 = {1'h1,T_849};
  assign T_852 = cyc_A2 ? T_850 : {{8'd0}, 1'h0};
  assign T_853 = T_847 | T_852;
  assign GEN_41 = T_836 ? T_853 : nextMulAdd9B_A;
  assign GEN_42 = cyc_A1_sqrt ? ER1_A1_sqrt : ER1_B_sqrt;
  assign T_854 = cyc_A1 | cyc_B7_sqrt;
  assign T_855 = T_854 | cyc_B6_div;
  assign T_856 = T_855 | cyc_B4;
  assign T_857 = T_856 | cyc_B3;
  assign T_858 = T_857 | cyc_C6_sqrt;
  assign T_859 = T_858 | cyc_C4;
  assign T_860 = T_859 | cyc_C1;
  assign GEN_107 = {{36'd0}, ER1_A1_sqrt};
  assign T_861 = GEN_107 << 36;
  assign T_863 = cyc_A1_sqrt ? T_861 : {{52'd0}, 1'h0};
  assign T_864 = cyc_B7_sqrt | cyc_A1_div;
  assign T_866 = T_864 ? sigB_PA : {{52'd0}, 1'h0};
  assign T_867 = T_863 | T_866;
  assign T_869 = cyc_B6_div ? sigA_PA : {{52'd0}, 1'h0};
  assign T_870 = T_867 | T_869;
  assign T_871 = zSigma1_B4[45:12];
  assign GEN_108 = {{19'd0}, T_871};
  assign T_872 = T_870 | GEN_108;
  assign T_873 = cyc_B3 | cyc_C6_sqrt;
  assign T_874 = sigXNU_B3_CX[57:12];
  assign T_876 = T_873 ? T_874 : {{45'd0}, 1'h0};
  assign GEN_109 = {{7'd0}, T_876};
  assign T_877 = T_872 | GEN_109;
  assign T_878 = sigXN_C[57:25];
  assign GEN_110 = {{13'd0}, T_878};
  assign T_879 = GEN_110 << 13;
  assign T_881 = cyc_C4_div ? T_879 : {{45'd0}, 1'h0};
  assign GEN_111 = {{7'd0}, T_881};
  assign T_882 = T_877 | GEN_111;
  assign GEN_112 = {{15'd0}, u_C_sqrt};
  assign T_883 = GEN_112 << 15;
  assign T_885 = cyc_C4_sqrt ? T_883 : {{45'd0}, 1'h0};
  assign GEN_113 = {{7'd0}, T_885};
  assign T_886 = T_882 | GEN_113;
  assign T_888 = cyc_C1_div ? sigB_PC : {{52'd0}, 1'h0};
  assign T_889 = T_886 | T_888;
  assign GEN_114 = {{1'd0}, T_889};
  assign T_890 = GEN_114 | zComplSigT_C1_sqrt;
  assign T_892 = T_854 | cyc_B6_sqrt;
  assign T_893 = T_892 | cyc_B4;
  assign T_894 = T_893 | cyc_C6_sqrt;
  assign T_895 = T_894 | cyc_C4;
  assign T_896 = T_895 | cyc_C1;
  assign GEN_115 = {{36'd0}, r1_A1};
  assign T_897 = GEN_115 << 36;
  assign T_899 = cyc_A1 ? T_897 : {{51'd0}, 1'h0};
  assign GEN_116 = {{19'd0}, ESqrR1_B_sqrt};
  assign T_900 = GEN_116 << 19;
  assign T_902 = cyc_B7_sqrt ? T_900 : {{50'd0}, 1'h0};
  assign GEN_117 = {{1'd0}, T_902};
  assign T_903 = T_899 | GEN_117;
  assign GEN_118 = {{36'd0}, ER1_B_sqrt};
  assign T_904 = GEN_118 << 36;
  assign T_906 = cyc_B6_sqrt ? T_904 : {{52'd0}, 1'h0};
  assign GEN_119 = {{1'd0}, T_903};
  assign T_907 = GEN_119 | T_906;
  assign GEN_120 = {{7'd0}, zSigma1_B4};
  assign T_908 = T_907 | GEN_120;
  assign T_909 = sqrSigma1_C[30:1];
  assign T_911 = cyc_C6_sqrt ? T_909 : {{29'd0}, 1'h0};
  assign GEN_121 = {{23'd0}, T_911};
  assign T_912 = T_908 | GEN_121;
  assign T_914 = cyc_C4 ? sqrSigma1_C : {{32'd0}, 1'h0};
  assign GEN_122 = {{20'd0}, T_914};
  assign T_915 = T_912 | GEN_122;
  assign GEN_123 = {{1'd0}, T_915};
  assign T_916 = GEN_123 | zComplSigT_C1;
  assign T_917 = cyc_A4 | cyc_A3_div;
  assign T_918 = T_917 | cyc_A1_div;
  assign T_919 = T_918 | cyc_B10_sqrt;
  assign T_920 = T_919 | cyc_B9_sqrt;
  assign T_921 = T_920 | cyc_B7_sqrt;
  assign T_922 = T_921 | cyc_B6;
  assign T_923 = T_922 | cyc_B5_sqrt;
  assign T_924 = T_923 | cyc_B3_sqrt;
  assign T_925 = T_924 | cyc_B2_div;
  assign T_926 = T_925 | cyc_B1_sqrt;
  assign T_927 = T_926 | cyc_C4;
  assign T_928 = cyc_A3 | cyc_A2_div;
  assign T_929 = T_928 | cyc_B9_sqrt;
  assign T_930 = T_929 | cyc_B8_sqrt;
  assign T_931 = T_930 | cyc_B6;
  assign T_932 = T_931 | cyc_B5;
  assign T_933 = T_932 | cyc_B4_sqrt;
  assign T_934 = T_933 | cyc_B2_sqrt;
  assign T_935 = T_934 | cyc_B1_div;
  assign T_936 = T_935 | cyc_C6_sqrt;
  assign T_937 = T_936 | valid_normalCase_leaving_PB;
  assign T_938 = cyc_A2 | cyc_A1_div;
  assign T_939 = T_938 | cyc_B8_sqrt;
  assign T_940 = T_939 | cyc_B7_sqrt;
  assign T_941 = T_940 | cyc_B5;
  assign T_942 = T_941 | cyc_B4;
  assign T_943 = T_942 | cyc_B3_sqrt;
  assign T_944 = T_943 | cyc_B1_sqrt;
  assign T_945 = T_944 | cyc_C5;
  assign T_946 = T_945 | cyc_C2;
  assign T_947 = io_latchMulAddA_0 | cyc_B6;
  assign T_948 = T_947 | cyc_B2_sqrt;
  assign T_949 = {T_946,T_948};
  assign T_950 = {T_927,T_937};
  assign T_951 = {T_950,T_949};
  assign GEN_124 = {{47'd0}, sigX1_B};
  assign T_952 = GEN_124 << 47;
  assign T_954 = cyc_B1 ? T_952 : {{104'd0}, 1'h0};
  assign GEN_125 = {{46'd0}, sigX1_B};
  assign T_955 = GEN_125 << 46;
  assign T_957 = cyc_C6_sqrt ? T_955 : {{103'd0}, 1'h0};
  assign GEN_126 = {{1'd0}, T_957};
  assign T_958 = T_954 | GEN_126;
  assign T_959 = cyc_C4_sqrt | cyc_C2;
  assign GEN_127 = {{47'd0}, sigXN_C};
  assign T_960 = GEN_127 << 47;
  assign T_962 = T_959 ? T_960 : {{104'd0}, 1'h0};
  assign T_963 = T_958 | T_962;
  assign T_965 = E_E_div == 1'h0;
  assign T_966 = cyc_E3_div & T_965;
  assign GEN_128 = {{53'd0}, fractA_0_PC};
  assign T_967 = GEN_128 << 53;
  assign T_969 = T_966 ? T_967 : {{53'd0}, 1'h0};
  assign GEN_129 = {{51'd0}, T_969};
  assign T_970 = T_963 | GEN_129;
  assign T_972 = sigB_PC[0];
  assign T_974 = {T_972,1'h0};
  assign T_975 = sigB_PC[1];
  assign T_977 = T_975 ^ T_972;
  assign T_979 = {T_977,T_972};
  assign T_980 = T_351 ? T_974 : T_979;
  assign T_982 = extraT_E == 1'h0;
  assign T_984 = {T_982,1'h0};
  assign T_985 = T_980 ^ T_984;
  assign GEN_130 = {{54'd0}, T_985};
  assign T_986 = GEN_130 << 54;
  assign T_988 = cyc_E3_sqrt ? T_986 : {{55'd0}, 1'h0};
  assign GEN_131 = {{49'd0}, T_988};
  assign T_989 = T_970 | GEN_131;
  assign ESqrR1_B8_sqrt = io_mulAddResult_3[103:72];
  assign T_990 = io_mulAddResult_3[90:45];
  assign T_991 = ~ T_990;
  assign T_993 = cyc_B4 ? T_991 : {{45'd0}, 1'h0};
  assign sqrSigma1_B1 = io_mulAddResult_3[79:47];
  assign T_994 = io_mulAddResult_3[104:47];
  assign T_995 = io_mulAddResult_3[104];
  assign E_C1_div = T_995 == 1'h0;
  assign T_998 = E_C1_div == 1'h0;
  assign T_999 = cyc_C1_div & T_998;
  assign T_1000 = T_999 | cyc_C1_sqrt;
  assign T_1001 = io_mulAddResult_3[104:51];
  assign T_1002 = ~ T_1001;
  assign T_1004 = T_1000 ? T_1002 : {{53'd0}, 1'h0};
  assign T_1005 = cyc_C1_div & E_C1_div;
  assign T_1007 = io_mulAddResult_3[102:50];
  assign T_1008 = ~ T_1007;
  assign T_1009 = {1'h0,T_1008};
  assign T_1011 = T_1005 ? T_1009 : {{53'd0}, 1'h0};
  assign T_1012 = T_1004 | T_1011;
  assign T_1016 = cyc_C1_sqrt ? T_1002 : {{53'd0}, 1'h0};
  assign sigT_C1 = ~ zComplSigT_C1;
  assign remT_E2 = io_mulAddResult_3[55:0];
  assign GEN_43 = cyc_B8_sqrt ? ESqrR1_B8_sqrt : ESqrR1_B_sqrt;
  assign GEN_44 = cyc_B3 ? sigXNU_B3_CX : sigX1_B;
  assign GEN_45 = cyc_B1 ? sqrSigma1_B1 : sqrSigma1_C;
  assign T_1017 = cyc_C6_sqrt | cyc_C5_div;
  assign T_1018 = T_1017 | cyc_C3_sqrt;
  assign GEN_46 = T_1018 ? sigXNU_B3_CX : sigXN_C;
  assign T_1019 = sigXNU_B3_CX[56:26];
  assign GEN_47 = cyc_C5_sqrt ? T_1019 : u_C_sqrt;
  assign T_1020 = sigT_C1[53:1];
  assign T_1021 = sigT_C1[0];
  assign GEN_48 = cyc_C1 ? E_C1_div : E_E_div;
  assign GEN_49 = cyc_C1 ? T_1020 : sigT_E;
  assign GEN_50 = cyc_C1 ? T_1021 : extraT_E;
  assign T_1022 = remT_E2[55];
  assign T_1023 = remT_E2[53];
  assign T_1024 = sqrtOp_PC ? T_1022 : T_1023;
  assign T_1025 = remT_E2[53:0];
  assign GEN_132 = {{53'd0}, 1'h0};
  assign T_1027 = T_1025 == GEN_132;
  assign T_1030 = remT_E2[55:54];
  assign GEN_133 = {{1'd0}, 1'h0};
  assign T_1032 = T_1030 == GEN_133;
  assign T_1033 = T_369 | T_1032;
  assign T_1034 = T_1027 & T_1033;
  assign GEN_51 = cyc_E2 ? T_1024 : isNegRemT_E;
  assign GEN_52 = cyc_E2 ? T_1034 : trueEqX_E1;
  assign T_1037 = T_369 & E_E_div;
  assign T_1039 = T_1037 ? exp_PC : {{13'd0}, 1'h0};
  assign T_1044 = T_369 & T_965;
  assign T_1046 = T_1044 ? expP1_PC : {{13'd0}, 1'h0};
  assign T_1047 = T_1039 | T_1046;
  assign T_1048 = exp_PC[13:1];
  assign GEN_134 = {{1'd0}, 12'h400};
  assign T_1050 = T_1048 + GEN_134;
  assign T_1051 = T_1050[12:0];
  assign T_1053 = sqrtOp_PC ? T_1051 : {{12'd0}, 1'h0};
  assign GEN_135 = {{1'd0}, T_1053};
  assign sExpX_E = T_1047 | GEN_135;
  assign posExpX_E = sExpX_E[12:0];
  assign T_1054 = ~ posExpX_E;
  assign GEN_136 = $signed(8193'h100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000);
  assign T_1056 = $signed(GEN_136) >>> T_1054;
  assign T_1057 = T_1056[1026:974];
  assign T_1058 = T_1057[31:0];
  assign T_1063 = T_1058[31:16];
  assign GEN_137 = {{16'd0}, T_1063};
  assign T_1064 = GEN_137 & 32'hffff;
  assign T_1065 = T_1058[15:0];
  assign GEN_138 = {{16'd0}, T_1065};
  assign T_1066 = GEN_138 << 16;
  assign T_1068 = T_1066 & 32'hffff0000;
  assign T_1069 = T_1064 | T_1068;
  assign T_1073 = T_1069[31:8];
  assign GEN_139 = {{8'd0}, T_1073};
  assign T_1074 = GEN_139 & 32'hff00ff;
  assign T_1075 = T_1069[23:0];
  assign GEN_140 = {{8'd0}, T_1075};
  assign T_1076 = GEN_140 << 8;
  assign T_1078 = T_1076 & 32'hff00ff00;
  assign T_1079 = T_1074 | T_1078;
  assign T_1083 = T_1079[31:4];
  assign GEN_141 = {{4'd0}, T_1083};
  assign T_1084 = GEN_141 & 32'hf0f0f0f;
  assign T_1085 = T_1079[27:0];
  assign GEN_142 = {{4'd0}, T_1085};
  assign T_1086 = GEN_142 << 4;
  assign T_1088 = T_1086 & 32'hf0f0f0f0;
  assign T_1089 = T_1084 | T_1088;
  assign T_1093 = T_1089[31:2];
  assign GEN_143 = {{2'd0}, T_1093};
  assign T_1094 = GEN_143 & 32'h33333333;
  assign T_1095 = T_1089[29:0];
  assign GEN_144 = {{2'd0}, T_1095};
  assign T_1096 = GEN_144 << 2;
  assign T_1098 = T_1096 & 32'hcccccccc;
  assign T_1099 = T_1094 | T_1098;
  assign T_1103 = T_1099[31:1];
  assign GEN_145 = {{1'd0}, T_1103};
  assign T_1104 = GEN_145 & 32'h55555555;
  assign T_1105 = T_1099[30:0];
  assign GEN_146 = {{1'd0}, T_1105};
  assign T_1106 = GEN_146 << 1;
  assign T_1108 = T_1106 & 32'haaaaaaaa;
  assign T_1109 = T_1104 | T_1108;
  assign T_1110 = T_1057[52:32];
  assign T_1111 = T_1110[15:0];
  assign T_1116 = T_1111[15:8];
  assign GEN_147 = {{8'd0}, T_1116};
  assign T_1117 = GEN_147 & 16'hff;
  assign T_1118 = T_1111[7:0];
  assign GEN_148 = {{8'd0}, T_1118};
  assign T_1119 = GEN_148 << 8;
  assign T_1121 = T_1119 & 16'hff00;
  assign T_1122 = T_1117 | T_1121;
  assign T_1126 = T_1122[15:4];
  assign GEN_149 = {{4'd0}, T_1126};
  assign T_1127 = GEN_149 & 16'hf0f;
  assign T_1128 = T_1122[11:0];
  assign GEN_150 = {{4'd0}, T_1128};
  assign T_1129 = GEN_150 << 4;
  assign T_1131 = T_1129 & 16'hf0f0;
  assign T_1132 = T_1127 | T_1131;
  assign T_1136 = T_1132[15:2];
  assign GEN_151 = {{2'd0}, T_1136};
  assign T_1137 = GEN_151 & 16'h3333;
  assign T_1138 = T_1132[13:0];
  assign GEN_152 = {{2'd0}, T_1138};
  assign T_1139 = GEN_152 << 2;
  assign T_1141 = T_1139 & 16'hcccc;
  assign T_1142 = T_1137 | T_1141;
  assign T_1146 = T_1142[15:1];
  assign GEN_153 = {{1'd0}, T_1146};
  assign T_1147 = GEN_153 & 16'h5555;
  assign T_1148 = T_1142[14:0];
  assign GEN_154 = {{1'd0}, T_1148};
  assign T_1149 = GEN_154 << 1;
  assign T_1151 = T_1149 & 16'haaaa;
  assign T_1152 = T_1147 | T_1151;
  assign T_1153 = T_1110[20:16];
  assign T_1154 = T_1153[3:0];
  assign T_1155 = T_1154[1:0];
  assign T_1156 = T_1155[0];
  assign T_1157 = T_1155[1];
  assign T_1158 = {T_1156,T_1157};
  assign T_1159 = T_1154[3:2];
  assign T_1160 = T_1159[0];
  assign T_1161 = T_1159[1];
  assign T_1162 = {T_1160,T_1161};
  assign T_1163 = {T_1158,T_1162};
  assign T_1164 = T_1153[4];
  assign T_1165 = {T_1163,T_1164};
  assign T_1166 = {T_1152,T_1165};
  assign roundMask_E = {T_1109,T_1166};
  assign T_1168 = {1'h0,roundMask_E};
  assign T_1169 = ~ T_1168;
  assign T_1171 = {roundMask_E,1'h1};
  assign incrPosMask_E = T_1169 & T_1171;
  assign T_1172 = incrPosMask_E[53:1];
  assign T_1173 = sigT_E & T_1172;
  assign GEN_155 = {{52'd0}, 1'h0};
  assign hiRoundPosBitT_E = T_1173 != GEN_155;
  assign T_1175 = roundMask_E[52:1];
  assign GEN_156 = {{1'd0}, T_1175};
  assign T_1178 = ~ sigT_E;
  assign T_1180 = T_1178 & GEN_156;
  assign all1sHiRoundExtraT_E = T_1180 == GEN_155;
  assign T_1182 = roundMask_E[0];
  assign T_1184 = T_1182 == 1'h0;
  assign T_1185 = T_1184 | hiRoundPosBitT_E;
  assign all1sHiRoundT_E = T_1185 & all1sHiRoundExtraT_E;
  assign GEN_160 = {{1'd0}, sigT_E};
  assign T_1187 = 54'h0 + GEN_160;
  assign T_1188 = T_1187[53:0];
  assign GEN_161 = {{53'd0}, roundMagUp_PC};
  assign T_1189 = T_1188 + GEN_161;
  assign sigAdjT_E = T_1189[53:0];
  assign T_1191 = ~ roundMask_E;
  assign T_1192 = {1'h1,T_1191};
  assign sigY0_E = sigAdjT_E & T_1192;
  assign T_1195 = sigAdjT_E | T_1168;
  assign GEN_162 = {{53'd0}, 1'h1};
  assign T_1197 = T_1195 + GEN_162;
  assign sigY1_E = T_1197[53:0];
  assign T_1199 = isNegRemT_E == 1'h0;
  assign T_1201 = trueEqX_E1 == 1'h0;
  assign T_1202 = T_1199 & T_1201;
  assign trueLtX_E1 = sqrtOp_PC ? T_1202 : isNegRemT_E;
  assign T_1205 = trueLtX_E1 == 1'h0;
  assign T_1206 = T_1182 & T_1205;
  assign T_1207 = T_1206 & all1sHiRoundExtraT_E;
  assign T_1208 = T_1207 & extraT_E;
  assign hiRoundPosBit_E1 = hiRoundPosBitT_E ^ T_1208;
  assign T_1213 = T_1201 | T_982;
  assign T_1215 = all1sHiRoundExtraT_E == 1'h0;
  assign anyRoundExtra_E1 = T_1213 | T_1215;
  assign T_1216 = roundingMode_near_even_PC & hiRoundPosBit_E1;
  assign T_1218 = anyRoundExtra_E1 == 1'h0;
  assign T_1219 = T_1216 & T_1218;
  assign roundEvenMask_E1 = T_1219 ? incrPosMask_E : {{53'd0}, 1'h0};
  assign T_1221 = roundMagDown_PC & extraT_E;
  assign T_1224 = T_1221 & T_1205;
  assign T_1225 = T_1224 & all1sHiRoundT_E;
  assign T_1228 = extraT_E & T_1205;
  assign T_1231 = T_1228 & T_1201;
  assign T_1233 = all1sHiRoundT_E == 1'h0;
  assign T_1234 = T_1231 | T_1233;
  assign T_1235 = roundMagUp_PC & T_1234;
  assign T_1236 = T_1225 | T_1235;
  assign T_1239 = extraT_E | T_1205;
  assign T_1243 = T_1239 & T_1184;
  assign T_1244 = hiRoundPosBitT_E | T_1243;
  assign T_1248 = T_1228 & all1sHiRoundExtraT_E;
  assign T_1249 = T_1244 | T_1248;
  assign T_1250 = roundingMode_near_even_PC & T_1249;
  assign T_1251 = T_1236 | T_1250;
  assign T_1252 = T_1251 ? sigY1_E : sigY0_E;
  assign T_1253 = ~ roundEvenMask_E1;
  assign sigY_E1 = T_1252 & T_1253;
  assign fractY_E1 = sigY_E1[51:0];
  assign inexactY_E1 = hiRoundPosBit_E1 | anyRoundExtra_E1;
  assign T_1254 = sigY_E1[53];
  assign T_1256 = T_1254 == 1'h0;
  assign T_1258 = T_1256 ? sExpX_E : {{13'd0}, 1'h0};
  assign T_1262 = T_1254 & T_369;
  assign T_1263 = T_1262 & E_E_div;
  assign T_1265 = T_1263 ? expP1_PC : {{13'd0}, 1'h0};
  assign T_1266 = T_1258 | T_1265;
  assign T_1273 = T_1262 & T_965;
  assign T_1275 = T_1273 ? expP2_PC : {{13'd0}, 1'h0};
  assign T_1276 = T_1266 | T_1275;
  assign T_1278 = T_1254 & sqrtOp_PC;
  assign T_1279 = expP2_PC[13:1];
  assign T_1281 = T_1279 + GEN_134;
  assign T_1282 = T_1281[12:0];
  assign T_1284 = T_1278 ? T_1282 : {{12'd0}, 1'h0};
  assign GEN_164 = {{1'd0}, T_1284};
  assign sExpY_E1 = T_1276 | GEN_164;
  assign expY_E1 = sExpY_E1[11:0];
  assign T_1285 = sExpY_E1[13];
  assign T_1287 = T_1285 == 1'h0;
  assign T_1289 = sExpY_E1[12:10];
  assign T_1290 = 3'h3 <= T_1289;
  assign overflowY_E1 = T_1287 & T_1290;
  assign T_1292 = sExpY_E1[12:0];
  assign T_1294 = T_1292 < 13'h3ce;
  assign totalUnderflowY_E1 = T_1285 | T_1294;
  assign T_1296 = posExpX_E <= 13'h401;
  assign T_1297 = T_1296 & inexactY_E1;
  assign underflowY_E1 = totalUnderflowY_E1 | T_1297;
  assign T_1299 = isNaNB_PC == 1'h0;
  assign T_1302 = T_1299 & T_333;
  assign T_1303 = T_1302 & sign_PC;
  assign T_1304 = isZeroA_PC & isZeroB_PC;
  assign T_1305 = isInfA_PC & isInfB_PC;
  assign T_1306 = T_1304 | T_1305;
  assign notSigNaN_invalid_PC = sqrtOp_PC ? T_1303 : T_1306;
  assign T_1309 = T_369 & isSigNaNA_PC;
  assign T_1310 = T_1309 | isSigNaNB_PC;
  assign invalid_PC = T_1310 | notSigNaN_invalid_PC;
  assign T_1315 = T_369 & T_339;
  assign T_1318 = T_1315 & T_344;
  assign infinity_PC = T_1318 & isZeroB_PC;
  assign overflow_E1 = normalCase_PC & overflowY_E1;
  assign underflow_E1 = normalCase_PC & underflowY_E1;
  assign T_1319 = overflow_E1 | underflow_E1;
  assign T_1320 = normalCase_PC & inexactY_E1;
  assign inexact_E1 = T_1319 | T_1320;
  assign T_1321 = isZeroA_PC | isInfB_PC;
  assign T_1324 = totalUnderflowY_E1 & T_359;
  assign T_1325 = T_1321 | T_1324;
  assign notSpecial_isZeroOut_E1 = sqrtOp_PC ? isZeroB_PC : T_1325;
  assign T_1326 = normalCase_PC & totalUnderflowY_E1;
  assign pegMinFiniteMagOut_E1 = T_1326 & roundMagUp_PC;
  assign T_1328 = overflowY_roundMagUp_PC == 1'h0;
  assign pegMaxFiniteMagOut_E1 = overflow_E1 & T_1328;
  assign T_1329 = isInfA_PC | isZeroB_PC;
  assign T_1330 = overflow_E1 & overflowY_roundMagUp_PC;
  assign T_1331 = T_1329 | T_1330;
  assign notNaN_isInfOut_E1 = sqrtOp_PC ? isInfB_PC : T_1331;
  assign T_1334 = T_369 & isNaNA_PC;
  assign T_1335 = T_1334 | isNaNB_PC;
  assign isNaNOut_PC = T_1335 | notSigNaN_invalid_PC;
  assign T_1337 = isNaNOut_PC == 1'h0;
  assign T_1338 = isZeroB_PC & sign_PC;
  assign T_1339 = sqrtOp_PC ? T_1338 : sign_PC;
  assign signOut_PC = T_1337 & T_1339;
  assign T_1343 = notSpecial_isZeroOut_E1 ? 12'he00 : {{11'd0}, 1'h0};
  assign T_1344 = ~ T_1343;
  assign T_1345 = expY_E1 & T_1344;
  assign T_1349 = pegMinFiniteMagOut_E1 ? 12'hc31 : {{11'd0}, 1'h0};
  assign T_1350 = ~ T_1349;
  assign T_1351 = T_1345 & T_1350;
  assign T_1355 = pegMaxFiniteMagOut_E1 ? 12'h400 : {{11'd0}, 1'h0};
  assign T_1356 = ~ T_1355;
  assign T_1357 = T_1351 & T_1356;
  assign T_1361 = notNaN_isInfOut_E1 ? 12'h200 : {{11'd0}, 1'h0};
  assign T_1362 = ~ T_1361;
  assign T_1363 = T_1357 & T_1362;
  assign T_1366 = pegMinFiniteMagOut_E1 ? 12'h3ce : {{11'd0}, 1'h0};
  assign T_1367 = T_1363 | T_1366;
  assign T_1370 = pegMaxFiniteMagOut_E1 ? 12'hbff : {{11'd0}, 1'h0};
  assign T_1371 = T_1367 | T_1370;
  assign T_1374 = notNaN_isInfOut_E1 ? 12'hc00 : {{11'd0}, 1'h0};
  assign T_1375 = T_1371 | T_1374;
  assign T_1378 = isNaNOut_PC ? 12'he00 : {{11'd0}, 1'h0};
  assign expOut_E1 = T_1375 | T_1378;
  assign T_1379 = notSpecial_isZeroOut_E1 | totalUnderflowY_E1;
  assign T_1380 = T_1379 | isNaNOut_PC;
  assign T_1384 = isNaNOut_PC ? 52'h8000000000000 : {{51'd0}, 1'h0};
  assign T_1385 = T_1380 ? T_1384 : fractY_E1;
  assign GEN_165 = {{51'd0}, pegMaxFiniteMagOut_E1};
  assign T_1387 = 52'h0 - GEN_165;
  assign T_1388 = T_1387[51:0];
  assign fractOut_E1 = T_1385 | T_1388;
  assign T_1389 = {signOut_PC,expOut_E1};
  assign T_1390 = {T_1389,fractOut_E1};
  assign T_1391 = {underflow_E1,inexact_E1};
  assign T_1392 = {invalid_PC,infinity_PC};
  assign T_1393 = {T_1392,overflow_E1};
  assign T_1394 = {T_1393,T_1391};
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_61 = {1{$random}};
  valid_PA = GEN_61[0:0];
  GEN_70 = {1{$random}};
  sqrtOp_PA = GEN_70[0:0];
  GEN_71 = {1{$random}};
  sign_PA = GEN_71[0:0];
  GEN_72 = {1{$random}};
  specialCodeB_PA = GEN_72[2:0];
  GEN_73 = {1{$random}};
  fractB_51_PA = GEN_73[0:0];
  GEN_74 = {1{$random}};
  roundingMode_PA = GEN_74[1:0];
  GEN_75 = {1{$random}};
  specialCodeA_PA = GEN_75[2:0];
  GEN_76 = {1{$random}};
  fractA_51_PA = GEN_76[0:0];
  GEN_77 = {1{$random}};
  exp_PA = GEN_77[13:0];
  GEN_78 = {2{$random}};
  fractB_other_PA = GEN_78[50:0];
  GEN_79 = {2{$random}};
  fractA_other_PA = GEN_79[50:0];
  GEN_80 = {1{$random}};
  valid_PB = GEN_80[0:0];
  GEN_81 = {1{$random}};
  sqrtOp_PB = GEN_81[0:0];
  GEN_82 = {1{$random}};
  sign_PB = GEN_82[0:0];
  GEN_83 = {1{$random}};
  specialCodeA_PB = GEN_83[2:0];
  GEN_84 = {1{$random}};
  fractA_51_PB = GEN_84[0:0];
  GEN_157 = {1{$random}};
  specialCodeB_PB = GEN_157[2:0];
  GEN_158 = {1{$random}};
  fractB_51_PB = GEN_158[0:0];
  GEN_159 = {1{$random}};
  roundingMode_PB = GEN_159[1:0];
  GEN_163 = {1{$random}};
  exp_PB = GEN_163[13:0];
  GEN_166 = {1{$random}};
  fractA_0_PB = GEN_166[0:0];
  GEN_167 = {2{$random}};
  fractB_other_PB = GEN_167[50:0];
  GEN_168 = {1{$random}};
  valid_PC = GEN_168[0:0];
  GEN_169 = {1{$random}};
  sqrtOp_PC = GEN_169[0:0];
  GEN_170 = {1{$random}};
  sign_PC = GEN_170[0:0];
  GEN_171 = {1{$random}};
  specialCodeA_PC = GEN_171[2:0];
  GEN_172 = {1{$random}};
  fractA_51_PC = GEN_172[0:0];
  GEN_173 = {1{$random}};
  specialCodeB_PC = GEN_173[2:0];
  GEN_174 = {1{$random}};
  fractB_51_PC = GEN_174[0:0];
  GEN_175 = {1{$random}};
  roundingMode_PC = GEN_175[1:0];
  GEN_176 = {1{$random}};
  exp_PC = GEN_176[13:0];
  GEN_177 = {1{$random}};
  fractA_0_PC = GEN_177[0:0];
  GEN_178 = {2{$random}};
  fractB_other_PC = GEN_178[50:0];
  GEN_179 = {1{$random}};
  cycleNum_A = GEN_179[2:0];
  GEN_180 = {1{$random}};
  cycleNum_B = GEN_180[3:0];
  GEN_181 = {1{$random}};
  cycleNum_C = GEN_181[2:0];
  GEN_182 = {1{$random}};
  cycleNum_E = GEN_182[2:0];
  GEN_183 = {1{$random}};
  fractR0_A = GEN_183[8:0];
  GEN_184 = {1{$random}};
  hiSqrR0_A_sqrt = GEN_184[9:0];
  GEN_185 = {1{$random}};
  partNegSigma0_A = GEN_185[20:0];
  GEN_186 = {1{$random}};
  nextMulAdd9A_A = GEN_186[8:0];
  GEN_187 = {1{$random}};
  nextMulAdd9B_A = GEN_187[8:0];
  GEN_188 = {1{$random}};
  ER1_B_sqrt = GEN_188[16:0];
  GEN_189 = {1{$random}};
  ESqrR1_B_sqrt = GEN_189[31:0];
  GEN_190 = {2{$random}};
  sigX1_B = GEN_190[57:0];
  GEN_191 = {2{$random}};
  sqrSigma1_C = GEN_191[32:0];
  GEN_192 = {2{$random}};
  sigXN_C = GEN_192[57:0];
  GEN_193 = {1{$random}};
  u_C_sqrt = GEN_193[30:0];
  GEN_194 = {1{$random}};
  E_E_div = GEN_194[0:0];
  GEN_195 = {2{$random}};
  sigT_E = GEN_195[52:0];
  GEN_196 = {1{$random}};
  extraT_E = GEN_196[0:0];
  GEN_197 = {1{$random}};
  isNegRemT_E = GEN_197[0:0];
  GEN_198 = {1{$random}};
  trueEqX_E1 = GEN_198[0:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      valid_PA <= 1'h0;
    end else begin
      valid_PA <= GEN_0;
    end
    if(1'h0) begin
    end else begin
      sqrtOp_PA <= GEN_1;
    end
    if(1'h0) begin
    end else begin
      sign_PA <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      specialCodeB_PA <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      fractB_51_PA <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      roundingMode_PA <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      specialCodeA_PA <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      fractA_51_PA <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      exp_PA <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      fractB_other_PA <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      fractA_other_PA <= GEN_10;
    end
    if(reset) begin
      valid_PB <= 1'h0;
    end else begin
      valid_PB <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      sqrtOp_PB <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      sign_PB <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      specialCodeA_PB <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      fractA_51_PB <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      specialCodeB_PB <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      fractB_51_PB <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      roundingMode_PB <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      exp_PB <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      fractA_0_PB <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      fractB_other_PB <= GEN_21;
    end
    if(reset) begin
      valid_PC <= 1'h0;
    end else begin
      valid_PC <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      sqrtOp_PC <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      sign_PC <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      specialCodeA_PC <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      fractA_51_PC <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      specialCodeB_PC <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      fractB_51_PC <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      roundingMode_PC <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      exp_PC <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      fractA_0_PC <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      fractB_other_PC <= GEN_32;
    end
    if(reset) begin
      cycleNum_A <= 3'h0;
    end else begin
      cycleNum_A <= GEN_33;
    end
    if(reset) begin
      cycleNum_B <= 4'h0;
    end else begin
      cycleNum_B <= GEN_34;
    end
    if(reset) begin
      cycleNum_C <= 3'h0;
    end else begin
      cycleNum_C <= GEN_35;
    end
    if(reset) begin
      cycleNum_E <= 3'h0;
    end else begin
      cycleNum_E <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      fractR0_A <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      hiSqrR0_A_sqrt <= GEN_38[9:0];
    end
    if(1'h0) begin
    end else begin
      partNegSigma0_A <= GEN_39;
    end
    if(1'h0) begin
    end else begin
      nextMulAdd9A_A <= GEN_40[8:0];
    end
    if(1'h0) begin
    end else begin
      nextMulAdd9B_A <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      ER1_B_sqrt <= GEN_42;
    end
    if(1'h0) begin
    end else begin
      ESqrR1_B_sqrt <= GEN_43;
    end
    if(1'h0) begin
    end else begin
      sigX1_B <= GEN_44;
    end
    if(1'h0) begin
    end else begin
      sqrSigma1_C <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      sigXN_C <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      u_C_sqrt <= GEN_47;
    end
    if(1'h0) begin
    end else begin
      E_E_div <= GEN_48;
    end
    if(1'h0) begin
    end else begin
      sigT_E <= GEN_49;
    end
    if(1'h0) begin
    end else begin
      extraT_E <= GEN_50;
    end
    if(1'h0) begin
    end else begin
      isNegRemT_E <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      trueEqX_E1 <= GEN_52;
    end
  end
endmodule
module Mul54(
  input   clk,
  input   reset,
  input   io_val_s0,
  input   io_latch_a_s0,
  input  [53:0] io_a_s0,
  input   io_latch_b_s0,
  input  [53:0] io_b_s0,
  input  [104:0] io_c_s2,
  output [104:0] io_result_s3
);
  reg  val_s1;
  reg [31:0] GEN_7;
  reg  val_s2;
  reg [31:0] GEN_8;
  reg [53:0] reg_a_s1;
  reg [63:0] GEN_9;
  reg [53:0] reg_b_s1;
  reg [63:0] GEN_10;
  reg [53:0] reg_a_s2;
  reg [63:0] GEN_11;
  reg [53:0] reg_b_s2;
  reg [63:0] GEN_12;
  reg [104:0] reg_result_s3;
  reg [127:0] GEN_13;
  wire [53:0] GEN_0;
  wire [53:0] GEN_1;
  wire [53:0] GEN_2;
  wire [53:0] GEN_3;
  wire [53:0] GEN_4;
  wire [53:0] GEN_5;
  wire [107:0] T_14;
  wire [104:0] T_15;
  wire [105:0] T_16;
  wire [104:0] T_17;
  wire [104:0] GEN_6;
  assign io_result_s3 = reg_result_s3;
  assign GEN_0 = io_latch_a_s0 ? io_a_s0 : reg_a_s1;
  assign GEN_1 = io_latch_b_s0 ? io_b_s0 : reg_b_s1;
  assign GEN_2 = io_val_s0 ? GEN_0 : reg_a_s1;
  assign GEN_3 = io_val_s0 ? GEN_1 : reg_b_s1;
  assign GEN_4 = val_s1 ? reg_a_s1 : reg_a_s2;
  assign GEN_5 = val_s1 ? reg_b_s1 : reg_b_s2;
  assign T_14 = reg_a_s2 * reg_b_s2;
  assign T_15 = T_14[104:0];
  assign T_16 = T_15 + io_c_s2;
  assign T_17 = T_16[104:0];
  assign GEN_6 = val_s2 ? T_17 : reg_result_s3;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_7 = {1{$random}};
  val_s1 = GEN_7[0:0];
  GEN_8 = {1{$random}};
  val_s2 = GEN_8[0:0];
  GEN_9 = {2{$random}};
  reg_a_s1 = GEN_9[53:0];
  GEN_10 = {2{$random}};
  reg_b_s1 = GEN_10[53:0];
  GEN_11 = {2{$random}};
  reg_a_s2 = GEN_11[53:0];
  GEN_12 = {2{$random}};
  reg_b_s2 = GEN_12[53:0];
  GEN_13 = {4{$random}};
  reg_result_s3 = GEN_13[104:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      val_s1 <= io_val_s0;
    end
    if(1'h0) begin
    end else begin
      val_s2 <= val_s1;
    end
    if(1'h0) begin
    end else begin
      reg_a_s1 <= GEN_2;
    end
    if(1'h0) begin
    end else begin
      reg_b_s1 <= GEN_3;
    end
    if(1'h0) begin
    end else begin
      reg_a_s2 <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      reg_b_s2 <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      reg_result_s3 <= GEN_6;
    end
  end
endmodule
module DivSqrtRecF64(
  input   clk,
  input   reset,
  output  io_inReady_div,
  output  io_inReady_sqrt,
  input   io_inValid,
  input   io_sqrtOp,
  input  [64:0] io_a,
  input  [64:0] io_b,
  input  [1:0] io_roundingMode,
  output  io_outValid_div,
  output  io_outValid_sqrt,
  output [64:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire  ds_clk;
  wire  ds_reset;
  wire  ds_io_inReady_div;
  wire  ds_io_inReady_sqrt;
  wire  ds_io_inValid;
  wire  ds_io_sqrtOp;
  wire [64:0] ds_io_a;
  wire [64:0] ds_io_b;
  wire [1:0] ds_io_roundingMode;
  wire  ds_io_outValid_div;
  wire  ds_io_outValid_sqrt;
  wire [64:0] ds_io_out;
  wire [4:0] ds_io_exceptionFlags;
  wire [3:0] ds_io_usingMulAdd;
  wire  ds_io_latchMulAddA_0;
  wire [53:0] ds_io_mulAddA_0;
  wire  ds_io_latchMulAddB_0;
  wire [53:0] ds_io_mulAddB_0;
  wire [104:0] ds_io_mulAddC_2;
  wire [104:0] ds_io_mulAddResult_3;
  wire  mul_clk;
  wire  mul_reset;
  wire  mul_io_val_s0;
  wire  mul_io_latch_a_s0;
  wire [53:0] mul_io_a_s0;
  wire  mul_io_latch_b_s0;
  wire [53:0] mul_io_b_s0;
  wire [104:0] mul_io_c_s2;
  wire [104:0] mul_io_result_s3;
  wire  T_11;
  DivSqrtRecF64_mulAddZ31 ds (
    .clk(ds_clk),
    .reset(ds_reset),
    .io_inReady_div(ds_io_inReady_div),
    .io_inReady_sqrt(ds_io_inReady_sqrt),
    .io_inValid(ds_io_inValid),
    .io_sqrtOp(ds_io_sqrtOp),
    .io_a(ds_io_a),
    .io_b(ds_io_b),
    .io_roundingMode(ds_io_roundingMode),
    .io_outValid_div(ds_io_outValid_div),
    .io_outValid_sqrt(ds_io_outValid_sqrt),
    .io_out(ds_io_out),
    .io_exceptionFlags(ds_io_exceptionFlags),
    .io_usingMulAdd(ds_io_usingMulAdd),
    .io_latchMulAddA_0(ds_io_latchMulAddA_0),
    .io_mulAddA_0(ds_io_mulAddA_0),
    .io_latchMulAddB_0(ds_io_latchMulAddB_0),
    .io_mulAddB_0(ds_io_mulAddB_0),
    .io_mulAddC_2(ds_io_mulAddC_2),
    .io_mulAddResult_3(ds_io_mulAddResult_3)
  );
  Mul54 mul (
    .clk(mul_clk),
    .reset(mul_reset),
    .io_val_s0(mul_io_val_s0),
    .io_latch_a_s0(mul_io_latch_a_s0),
    .io_a_s0(mul_io_a_s0),
    .io_latch_b_s0(mul_io_latch_b_s0),
    .io_b_s0(mul_io_b_s0),
    .io_c_s2(mul_io_c_s2),
    .io_result_s3(mul_io_result_s3)
  );
  assign io_inReady_div = ds_io_inReady_div;
  assign io_inReady_sqrt = ds_io_inReady_sqrt;
  assign io_outValid_div = ds_io_outValid_div;
  assign io_outValid_sqrt = ds_io_outValid_sqrt;
  assign io_out = ds_io_out;
  assign io_exceptionFlags = ds_io_exceptionFlags;
  assign ds_clk = clk;
  assign ds_reset = reset;
  assign ds_io_inValid = io_inValid;
  assign ds_io_sqrtOp = io_sqrtOp;
  assign ds_io_a = io_a;
  assign ds_io_b = io_b;
  assign ds_io_roundingMode = io_roundingMode;
  assign ds_io_mulAddResult_3 = mul_io_result_s3;
  assign mul_clk = clk;
  assign mul_reset = reset;
  assign mul_io_val_s0 = T_11;
  assign mul_io_latch_a_s0 = ds_io_latchMulAddA_0;
  assign mul_io_a_s0 = ds_io_mulAddA_0;
  assign mul_io_latch_b_s0 = ds_io_latchMulAddB_0;
  assign mul_io_b_s0 = ds_io_mulAddB_0;
  assign mul_io_c_s2 = ds_io_mulAddC_2;
  assign T_11 = ds_io_usingMulAdd[0];
endmodule
module RecFNToRecFN_99(
  input   clk,
  input   reset,
  input  [64:0] io_in,
  input  [1:0] io_roundingMode,
  output [32:0] io_out,
  output [4:0] io_exceptionFlags
);
  wire [11:0] T_4;
  wire [1:0] T_5;
  wire  T_7;
  wire  T_15_sign;
  wire  T_15_isNaN;
  wire  T_15_isInf;
  wire  T_15_isZero;
  wire [12:0] T_15_sExp;
  wire [55:0] T_15_sig;
  wire  T_22;
  wire  T_23;
  wire  T_24;
  wire  T_27;
  wire  T_28;
  wire [2:0] T_29;
  wire [2:0] GEN_0;
  wire  T_31;
  wire [12:0] T_32;
  wire [51:0] T_34;
  wire [53:0] T_36;
  wire [55:0] T_37;
  wire [11:0] GEN_1;
  wire [12:0] GEN_2;
  wire [13:0] T_39;
  wire [12:0] T_40;
  wire [12:0] T_41;
  wire  outRawFloat_sign;
  wire  outRawFloat_isNaN;
  wire  outRawFloat_isInf;
  wire  outRawFloat_isZero;
  wire [9:0] outRawFloat_sExp;
  wire [26:0] outRawFloat_sig;
  wire  GEN_3;
  wire [12:0] GEN_4;
  wire  T_56;
  wire [2:0] T_57;
  wire  T_59;
  wire [8:0] T_67;
  wire [8:0] T_68;
  wire [9:0] T_69;
  wire [9:0] T_70;
  wire [25:0] T_71;
  wire [29:0] T_72;
  wire [29:0] GEN_6;
  wire  T_74;
  wire [26:0] T_75;
  wire  T_76;
  wire  T_78;
  wire  invalidExc;
  wire  RoundRawFNToRecFN_100_79_clk;
  wire  RoundRawFNToRecFN_100_79_reset;
  wire  RoundRawFNToRecFN_100_79_io_invalidExc;
  wire  RoundRawFNToRecFN_100_79_io_infiniteExc;
  wire  RoundRawFNToRecFN_100_79_io_in_sign;
  wire  RoundRawFNToRecFN_100_79_io_in_isNaN;
  wire  RoundRawFNToRecFN_100_79_io_in_isInf;
  wire  RoundRawFNToRecFN_100_79_io_in_isZero;
  wire [9:0] RoundRawFNToRecFN_100_79_io_in_sExp;
  wire [26:0] RoundRawFNToRecFN_100_79_io_in_sig;
  wire [1:0] RoundRawFNToRecFN_100_79_io_roundingMode;
  wire [32:0] RoundRawFNToRecFN_100_79_io_out;
  wire [4:0] RoundRawFNToRecFN_100_79_io_exceptionFlags;
  RoundRawFNToRecFN RoundRawFNToRecFN_100_79 (
    .clk(RoundRawFNToRecFN_100_79_clk),
    .reset(RoundRawFNToRecFN_100_79_reset),
    .io_invalidExc(RoundRawFNToRecFN_100_79_io_invalidExc),
    .io_infiniteExc(RoundRawFNToRecFN_100_79_io_infiniteExc),
    .io_in_sign(RoundRawFNToRecFN_100_79_io_in_sign),
    .io_in_isNaN(RoundRawFNToRecFN_100_79_io_in_isNaN),
    .io_in_isInf(RoundRawFNToRecFN_100_79_io_in_isInf),
    .io_in_isZero(RoundRawFNToRecFN_100_79_io_in_isZero),
    .io_in_sExp(RoundRawFNToRecFN_100_79_io_in_sExp),
    .io_in_sig(RoundRawFNToRecFN_100_79_io_in_sig),
    .io_roundingMode(RoundRawFNToRecFN_100_79_io_roundingMode),
    .io_out(RoundRawFNToRecFN_100_79_io_out),
    .io_exceptionFlags(RoundRawFNToRecFN_100_79_io_exceptionFlags)
  );
  assign io_out = RoundRawFNToRecFN_100_79_io_out;
  assign io_exceptionFlags = RoundRawFNToRecFN_100_79_io_exceptionFlags;
  assign T_4 = io_in[63:52];
  assign T_5 = T_4[11:10];
  assign T_7 = T_5 == 2'h3;
  assign T_15_sign = T_22;
  assign T_15_isNaN = T_24;
  assign T_15_isInf = T_28;
  assign T_15_isZero = T_31;
  assign T_15_sExp = T_32;
  assign T_15_sig = T_37;
  assign T_22 = io_in[64];
  assign T_23 = T_4[9];
  assign T_24 = T_7 & T_23;
  assign T_27 = T_23 == 1'h0;
  assign T_28 = T_7 & T_27;
  assign T_29 = T_4[11:9];
  assign GEN_0 = {{2'd0}, 1'h0};
  assign T_31 = T_29 == GEN_0;
  assign T_32 = {1'b0,$signed(T_4)};
  assign T_34 = io_in[51:0];
  assign T_36 = {2'h1,T_34};
  assign T_37 = {T_36,2'h0};
  assign GEN_1 = $signed(12'h900);
  assign GEN_2 = {{1{GEN_1[11]}},GEN_1};
  assign T_39 = $signed(T_15_sExp) + $signed(GEN_2);
  assign T_40 = T_39[12:0];
  assign T_41 = $signed(T_40);
  assign outRawFloat_sign = T_15_sign;
  assign outRawFloat_isNaN = T_15_isNaN;
  assign outRawFloat_isInf = T_15_isInf;
  assign outRawFloat_isZero = T_15_isZero;
  assign outRawFloat_sExp = T_70;
  assign outRawFloat_sig = T_75;
  assign GEN_3 = $signed(1'h0);
  assign GEN_4 = {13{GEN_3}};
  assign T_56 = $signed(T_41) < $signed(GEN_4);
  assign T_57 = T_41[11:9];
  assign T_59 = T_57 != GEN_0;
  assign T_67 = T_41[8:0];
  assign T_68 = T_59 ? 9'h1fc : T_67;
  assign T_69 = {T_56,T_68};
  assign T_70 = $signed(T_69);
  assign T_71 = T_15_sig[55:30];
  assign T_72 = T_15_sig[29:0];
  assign GEN_6 = {{29'd0}, 1'h0};
  assign T_74 = T_72 != GEN_6;
  assign T_75 = {T_71,T_74};
  assign T_76 = outRawFloat_sig[24];
  assign T_78 = T_76 == 1'h0;
  assign invalidExc = outRawFloat_isNaN & T_78;
  assign RoundRawFNToRecFN_100_79_clk = clk;
  assign RoundRawFNToRecFN_100_79_reset = reset;
  assign RoundRawFNToRecFN_100_79_io_invalidExc = invalidExc;
  assign RoundRawFNToRecFN_100_79_io_infiniteExc = 1'h0;
  assign RoundRawFNToRecFN_100_79_io_in_sign = outRawFloat_sign;
  assign RoundRawFNToRecFN_100_79_io_in_isNaN = outRawFloat_isNaN;
  assign RoundRawFNToRecFN_100_79_io_in_isInf = outRawFloat_isInf;
  assign RoundRawFNToRecFN_100_79_io_in_isZero = outRawFloat_isZero;
  assign RoundRawFNToRecFN_100_79_io_in_sExp = outRawFloat_sExp;
  assign RoundRawFNToRecFN_100_79_io_in_sig = outRawFloat_sig;
  assign RoundRawFNToRecFN_100_79_io_roundingMode = io_roundingMode;
endmodule
module FPU(
  input   clk,
  input   reset,
  input  [31:0] io_inst,
  input  [63:0] io_fromint_data,
  input  [2:0] io_fcsr_rm,
  output  io_fcsr_flags_valid,
  output [4:0] io_fcsr_flags_bits,
  output [63:0] io_store_data,
  output [63:0] io_toint_data,
  input   io_dmem_resp_val,
  input  [2:0] io_dmem_resp_type,
  input  [4:0] io_dmem_resp_tag,
  input  [63:0] io_dmem_resp_data,
  input   io_valid,
  output  io_fcsr_rdy,
  output  io_nack_mem,
  output  io_illegal_rm,
  input   io_killx,
  input   io_killm,
  output [4:0] io_dec_cmd,
  output  io_dec_ldst,
  output  io_dec_wen,
  output  io_dec_ren1,
  output  io_dec_ren2,
  output  io_dec_ren3,
  output  io_dec_swap12,
  output  io_dec_swap23,
  output  io_dec_single,
  output  io_dec_fromint,
  output  io_dec_toint,
  output  io_dec_fastpipe,
  output  io_dec_fma,
  output  io_dec_div,
  output  io_dec_sqrt,
  output  io_dec_round,
  output  io_dec_wflags,
  output  io_sboard_set,
  output  io_sboard_clr,
  output [4:0] io_sboard_clra,
  output  io_cp_req_ready,
  input   io_cp_req_valid,
  input  [4:0] io_cp_req_bits_cmd,
  input   io_cp_req_bits_ldst,
  input   io_cp_req_bits_wen,
  input   io_cp_req_bits_ren1,
  input   io_cp_req_bits_ren2,
  input   io_cp_req_bits_ren3,
  input   io_cp_req_bits_swap12,
  input   io_cp_req_bits_swap23,
  input   io_cp_req_bits_single,
  input   io_cp_req_bits_fromint,
  input   io_cp_req_bits_toint,
  input   io_cp_req_bits_fastpipe,
  input   io_cp_req_bits_fma,
  input   io_cp_req_bits_div,
  input   io_cp_req_bits_sqrt,
  input   io_cp_req_bits_round,
  input   io_cp_req_bits_wflags,
  input  [2:0] io_cp_req_bits_rm,
  input  [1:0] io_cp_req_bits_typ,
  input  [64:0] io_cp_req_bits_in1,
  input  [64:0] io_cp_req_bits_in2,
  input  [64:0] io_cp_req_bits_in3,
  input   io_cp_resp_ready,
  output  io_cp_resp_valid,
  output [64:0] io_cp_resp_bits_data,
  output [4:0] io_cp_resp_bits_exc
);
  reg  ex_reg_valid;
  reg [31:0] GEN_59;
  wire  req_valid;
  reg [31:0] ex_reg_inst;
  reg [31:0] GEN_60;
  wire [31:0] GEN_2;
  wire  T_193;
  wire  ex_cp_valid;
  wire  T_195;
  wire  T_196;
  wire  T_197;
  reg  mem_reg_valid;
  reg [31:0] GEN_61;
  reg [31:0] mem_reg_inst;
  reg [31:0] GEN_62;
  wire [31:0] GEN_3;
  reg  mem_cp_valid;
  reg [31:0] GEN_78;
  wire  T_200;
  wire  T_202;
  wire  killm;
  wire  T_204;
  wire  T_205;
  wire  T_206;
  reg  wb_reg_valid;
  reg [31:0] GEN_90;
  reg  wb_cp_valid;
  reg [31:0] GEN_91;
  wire  fp_decoder_clk;
  wire  fp_decoder_reset;
  wire [31:0] fp_decoder_io_inst;
  wire [4:0] fp_decoder_io_sigs_cmd;
  wire  fp_decoder_io_sigs_ldst;
  wire  fp_decoder_io_sigs_wen;
  wire  fp_decoder_io_sigs_ren1;
  wire  fp_decoder_io_sigs_ren2;
  wire  fp_decoder_io_sigs_ren3;
  wire  fp_decoder_io_sigs_swap12;
  wire  fp_decoder_io_sigs_swap23;
  wire  fp_decoder_io_sigs_single;
  wire  fp_decoder_io_sigs_fromint;
  wire  fp_decoder_io_sigs_toint;
  wire  fp_decoder_io_sigs_fastpipe;
  wire  fp_decoder_io_sigs_fma;
  wire  fp_decoder_io_sigs_div;
  wire  fp_decoder_io_sigs_sqrt;
  wire  fp_decoder_io_sigs_round;
  wire  fp_decoder_io_sigs_wflags;
  wire [4:0] cp_ctrl_cmd;
  wire  cp_ctrl_ldst;
  wire  cp_ctrl_wen;
  wire  cp_ctrl_ren1;
  wire  cp_ctrl_ren2;
  wire  cp_ctrl_ren3;
  wire  cp_ctrl_swap12;
  wire  cp_ctrl_swap23;
  wire  cp_ctrl_single;
  wire  cp_ctrl_fromint;
  wire  cp_ctrl_toint;
  wire  cp_ctrl_fastpipe;
  wire  cp_ctrl_fma;
  wire  cp_ctrl_div;
  wire  cp_ctrl_sqrt;
  wire  cp_ctrl_round;
  wire  cp_ctrl_wflags;
  reg [4:0] T_246_cmd;
  reg [31:0] GEN_92;
  reg  T_246_ldst;
  reg [31:0] GEN_93;
  reg  T_246_wen;
  reg [31:0] GEN_94;
  reg  T_246_ren1;
  reg [31:0] GEN_150;
  reg  T_246_ren2;
  reg [31:0] GEN_152;
  reg  T_246_ren3;
  reg [31:0] GEN_153;
  reg  T_246_swap12;
  reg [31:0] GEN_154;
  reg  T_246_swap23;
  reg [31:0] GEN_155;
  reg  T_246_single;
  reg [31:0] GEN_156;
  reg  T_246_fromint;
  reg [31:0] GEN_157;
  reg  T_246_toint;
  reg [31:0] GEN_158;
  reg  T_246_fastpipe;
  reg [31:0] GEN_159;
  reg  T_246_fma;
  reg [31:0] GEN_160;
  reg  T_246_div;
  reg [31:0] GEN_161;
  reg  T_246_sqrt;
  reg [31:0] GEN_162;
  reg  T_246_round;
  reg [31:0] GEN_163;
  reg  T_246_wflags;
  reg [31:0] GEN_164;
  wire [4:0] GEN_4;
  wire  GEN_5;
  wire  GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire  GEN_11;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_15;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  GEN_19;
  wire  GEN_20;
  wire [4:0] ex_ctrl_cmd;
  wire  ex_ctrl_ldst;
  wire  ex_ctrl_wen;
  wire  ex_ctrl_ren1;
  wire  ex_ctrl_ren2;
  wire  ex_ctrl_ren3;
  wire  ex_ctrl_swap12;
  wire  ex_ctrl_swap23;
  wire  ex_ctrl_single;
  wire  ex_ctrl_fromint;
  wire  ex_ctrl_toint;
  wire  ex_ctrl_fastpipe;
  wire  ex_ctrl_fma;
  wire  ex_ctrl_div;
  wire  ex_ctrl_sqrt;
  wire  ex_ctrl_round;
  wire  ex_ctrl_wflags;
  reg [4:0] mem_ctrl_cmd;
  reg [31:0] GEN_165;
  reg  mem_ctrl_ldst;
  reg [31:0] GEN_166;
  reg  mem_ctrl_wen;
  reg [31:0] GEN_167;
  reg  mem_ctrl_ren1;
  reg [31:0] GEN_168;
  reg  mem_ctrl_ren2;
  reg [31:0] GEN_169;
  reg  mem_ctrl_ren3;
  reg [31:0] GEN_170;
  reg  mem_ctrl_swap12;
  reg [31:0] GEN_171;
  reg  mem_ctrl_swap23;
  reg [31:0] GEN_172;
  reg  mem_ctrl_single;
  reg [31:0] GEN_173;
  reg  mem_ctrl_fromint;
  reg [31:0] GEN_174;
  reg  mem_ctrl_toint;
  reg [31:0] GEN_175;
  reg  mem_ctrl_fastpipe;
  reg [31:0] GEN_176;
  reg  mem_ctrl_fma;
  reg [31:0] GEN_177;
  reg  mem_ctrl_div;
  reg [31:0] GEN_178;
  reg  mem_ctrl_sqrt;
  reg [31:0] GEN_179;
  reg  mem_ctrl_round;
  reg [31:0] GEN_180;
  reg  mem_ctrl_wflags;
  reg [31:0] GEN_181;
  wire [4:0] GEN_21;
  wire  GEN_22;
  wire  GEN_23;
  wire  GEN_24;
  wire  GEN_25;
  wire  GEN_26;
  wire  GEN_27;
  wire  GEN_28;
  wire  GEN_29;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  GEN_33;
  wire  GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire  GEN_37;
  reg [4:0] wb_ctrl_cmd;
  reg [31:0] GEN_182;
  reg  wb_ctrl_ldst;
  reg [31:0] GEN_183;
  reg  wb_ctrl_wen;
  reg [31:0] GEN_184;
  reg  wb_ctrl_ren1;
  reg [31:0] GEN_185;
  reg  wb_ctrl_ren2;
  reg [31:0] GEN_186;
  reg  wb_ctrl_ren3;
  reg [31:0] GEN_187;
  reg  wb_ctrl_swap12;
  reg [31:0] GEN_188;
  reg  wb_ctrl_swap23;
  reg [31:0] GEN_189;
  reg  wb_ctrl_single;
  reg [31:0] GEN_190;
  reg  wb_ctrl_fromint;
  reg [31:0] GEN_191;
  reg  wb_ctrl_toint;
  reg [31:0] GEN_192;
  reg  wb_ctrl_fastpipe;
  reg [31:0] GEN_193;
  reg  wb_ctrl_fma;
  reg [31:0] GEN_194;
  reg  wb_ctrl_div;
  reg [31:0] GEN_195;
  reg  wb_ctrl_sqrt;
  reg [31:0] GEN_196;
  reg  wb_ctrl_round;
  reg [31:0] GEN_197;
  reg  wb_ctrl_wflags;
  reg [31:0] GEN_198;
  wire [4:0] GEN_38;
  wire  GEN_39;
  wire  GEN_40;
  wire  GEN_41;
  wire  GEN_42;
  wire  GEN_43;
  wire  GEN_44;
  wire  GEN_45;
  wire  GEN_46;
  wire  GEN_47;
  wire  GEN_48;
  wire  GEN_49;
  wire  GEN_50;
  wire  GEN_51;
  wire  GEN_52;
  wire  GEN_53;
  wire  GEN_54;
  reg  load_wb;
  reg [31:0] GEN_199;
  wire  T_315;
  wire  T_316;
  wire  T_317;
  reg  load_wb_single;
  reg [31:0] GEN_200;
  wire  GEN_55;
  reg [63:0] load_wb_data;
  reg [63:0] GEN_201;
  wire [63:0] GEN_56;
  reg [4:0] load_wb_tag;
  reg [31:0] GEN_202;
  wire [4:0] GEN_57;
  wire  T_318;
  wire [7:0] T_319;
  wire [22:0] T_320;
  wire [7:0] GEN_110;
  wire  T_322;
  wire [22:0] GEN_111;
  wire  T_324;
  wire  T_325;
  wire [31:0] GEN_112;
  wire [31:0] T_326;
  wire  T_327;
  wire  T_329;
  wire  T_331;
  wire  T_333;
  wire  T_335;
  wire  T_337;
  wire  T_339;
  wire  T_341;
  wire  T_343;
  wire  T_345;
  wire  T_347;
  wire  T_349;
  wire  T_351;
  wire  T_353;
  wire  T_355;
  wire  T_357;
  wire  T_359;
  wire  T_361;
  wire  T_363;
  wire  T_365;
  wire  T_367;
  wire  T_369;
  wire  T_371;
  wire  T_373;
  wire  T_375;
  wire  T_377;
  wire  T_379;
  wire  T_381;
  wire  T_383;
  wire  T_385;
  wire  T_387;
  wire [1:0] T_389;
  wire [1:0] T_390;
  wire [2:0] T_391;
  wire [2:0] T_392;
  wire [2:0] T_393;
  wire [2:0] T_394;
  wire [3:0] T_395;
  wire [3:0] T_396;
  wire [3:0] T_397;
  wire [3:0] T_398;
  wire [3:0] T_399;
  wire [3:0] T_400;
  wire [3:0] T_401;
  wire [3:0] T_402;
  wire [4:0] T_403;
  wire [4:0] T_404;
  wire [4:0] T_405;
  wire [4:0] T_406;
  wire [4:0] T_407;
  wire [4:0] T_408;
  wire [4:0] T_409;
  wire [4:0] T_410;
  wire [4:0] T_411;
  wire [4:0] T_412;
  wire [4:0] T_413;
  wire [4:0] T_414;
  wire [4:0] T_415;
  wire [4:0] T_416;
  wire [4:0] T_417;
  wire [4:0] T_418;
  wire [4:0] T_419;
  wire [53:0] GEN_113;
  wire [53:0] T_420;
  wire [21:0] T_421;
  wire [22:0] T_423;
  wire [8:0] GEN_114;
  wire [9:0] T_426;
  wire [8:0] T_427;
  wire [8:0] GEN_115;
  wire [8:0] T_428;
  wire [8:0] T_429;
  wire [1:0] T_433;
  wire [7:0] GEN_116;
  wire [7:0] T_434;
  wire [8:0] GEN_117;
  wire [9:0] T_435;
  wire [8:0] T_436;
  wire [1:0] T_437;
  wire  T_439;
  wire  T_441;
  wire  T_442;
  wire [2:0] GEN_118;
  wire [3:0] T_444;
  wire [2:0] T_445;
  wire [8:0] GEN_119;
  wire [8:0] T_446;
  wire [8:0] T_447;
  wire [8:0] T_448;
  wire [6:0] GEN_120;
  wire [6:0] T_449;
  wire [8:0] GEN_121;
  wire [8:0] T_450;
  wire [22:0] T_451;
  wire [9:0] T_452;
  wire [32:0] rec_s;
  wire  T_453;
  wire [10:0] T_454;
  wire [51:0] T_455;
  wire [10:0] GEN_122;
  wire  T_457;
  wire [51:0] GEN_123;
  wire  T_459;
  wire  T_460;
  wire [63:0] GEN_124;
  wire [63:0] T_461;
  wire  T_462;
  wire  T_464;
  wire  T_466;
  wire  T_468;
  wire  T_470;
  wire  T_472;
  wire  T_474;
  wire  T_476;
  wire  T_478;
  wire  T_480;
  wire  T_482;
  wire  T_484;
  wire  T_486;
  wire  T_488;
  wire  T_490;
  wire  T_492;
  wire  T_494;
  wire  T_496;
  wire  T_498;
  wire  T_500;
  wire  T_502;
  wire  T_504;
  wire  T_506;
  wire  T_508;
  wire  T_510;
  wire  T_512;
  wire  T_514;
  wire  T_516;
  wire  T_518;
  wire  T_520;
  wire  T_522;
  wire  T_524;
  wire  T_526;
  wire  T_528;
  wire  T_530;
  wire  T_532;
  wire  T_534;
  wire  T_536;
  wire  T_538;
  wire  T_540;
  wire  T_542;
  wire  T_544;
  wire  T_546;
  wire  T_548;
  wire  T_550;
  wire  T_552;
  wire  T_554;
  wire  T_556;
  wire  T_558;
  wire  T_560;
  wire  T_562;
  wire  T_564;
  wire  T_566;
  wire  T_568;
  wire  T_570;
  wire  T_572;
  wire  T_574;
  wire  T_576;
  wire  T_578;
  wire  T_580;
  wire  T_582;
  wire  T_584;
  wire  T_586;
  wire [1:0] T_588;
  wire [1:0] T_589;
  wire [2:0] T_590;
  wire [2:0] T_591;
  wire [2:0] T_592;
  wire [2:0] T_593;
  wire [3:0] T_594;
  wire [3:0] T_595;
  wire [3:0] T_596;
  wire [3:0] T_597;
  wire [3:0] T_598;
  wire [3:0] T_599;
  wire [3:0] T_600;
  wire [3:0] T_601;
  wire [4:0] T_602;
  wire [4:0] T_603;
  wire [4:0] T_604;
  wire [4:0] T_605;
  wire [4:0] T_606;
  wire [4:0] T_607;
  wire [4:0] T_608;
  wire [4:0] T_609;
  wire [4:0] T_610;
  wire [4:0] T_611;
  wire [4:0] T_612;
  wire [4:0] T_613;
  wire [4:0] T_614;
  wire [4:0] T_615;
  wire [4:0] T_616;
  wire [4:0] T_617;
  wire [5:0] T_618;
  wire [5:0] T_619;
  wire [5:0] T_620;
  wire [5:0] T_621;
  wire [5:0] T_622;
  wire [5:0] T_623;
  wire [5:0] T_624;
  wire [5:0] T_625;
  wire [5:0] T_626;
  wire [5:0] T_627;
  wire [5:0] T_628;
  wire [5:0] T_629;
  wire [5:0] T_630;
  wire [5:0] T_631;
  wire [5:0] T_632;
  wire [5:0] T_633;
  wire [5:0] T_634;
  wire [5:0] T_635;
  wire [5:0] T_636;
  wire [5:0] T_637;
  wire [5:0] T_638;
  wire [5:0] T_639;
  wire [5:0] T_640;
  wire [5:0] T_641;
  wire [5:0] T_642;
  wire [5:0] T_643;
  wire [5:0] T_644;
  wire [5:0] T_645;
  wire [5:0] T_646;
  wire [5:0] T_647;
  wire [5:0] T_648;
  wire [5:0] T_649;
  wire [5:0] T_650;
  wire [114:0] GEN_125;
  wire [114:0] T_651;
  wire [50:0] T_652;
  wire [51:0] T_654;
  wire [11:0] GEN_126;
  wire [12:0] T_657;
  wire [11:0] T_658;
  wire [11:0] GEN_127;
  wire [11:0] T_659;
  wire [11:0] T_660;
  wire [1:0] T_664;
  wire [10:0] GEN_128;
  wire [10:0] T_665;
  wire [11:0] GEN_129;
  wire [12:0] T_666;
  wire [11:0] T_667;
  wire [1:0] T_668;
  wire  T_670;
  wire  T_672;
  wire  T_673;
  wire [2:0] GEN_130;
  wire [3:0] T_675;
  wire [2:0] T_676;
  wire [11:0] GEN_131;
  wire [11:0] T_677;
  wire [11:0] T_678;
  wire [11:0] T_679;
  wire [9:0] GEN_132;
  wire [9:0] T_680;
  wire [11:0] GEN_133;
  wire [11:0] T_681;
  wire [51:0] T_682;
  wire [12:0] T_683;
  wire [64:0] rec_d;
  wire [31:0] GEN_134;
  wire [31:0] T_685;
  wire [64:0] T_686;
  wire [64:0] load_wb_data_recoded;
  reg [64:0] regfile [0:31];
  reg [95:0] GEN_203;
  wire [64:0] regfile_ex_rs1_data;
  wire [4:0] regfile_ex_rs1_addr;
  wire  regfile_ex_rs1_en;
  wire [64:0] regfile_ex_rs2_data;
  wire [4:0] regfile_ex_rs2_addr;
  wire  regfile_ex_rs2_en;
  wire [64:0] regfile_ex_rs3_data;
  wire [4:0] regfile_ex_rs3_addr;
  wire  regfile_ex_rs3_en;
  wire [64:0] regfile_T_689_data;
  wire [4:0] regfile_T_689_addr;
  wire  regfile_T_689_mask;
  wire  regfile_T_689_en;
  wire [64:0] regfile_T_919_data;
  wire [4:0] regfile_T_919_addr;
  wire  regfile_T_919_mask;
  wire  regfile_T_919_en;
  reg [4:0] ex_ra1;
  reg [31:0] GEN_204;
  reg [4:0] ex_ra2;
  reg [31:0] GEN_205;
  reg [4:0] ex_ra3;
  reg [31:0] GEN_206;
  wire  T_694;
  wire [4:0] T_695;
  wire [4:0] GEN_63;
  wire [4:0] GEN_64;
  wire [4:0] GEN_65;
  wire [4:0] GEN_66;
  wire [4:0] T_697;
  wire [4:0] GEN_67;
  wire [4:0] GEN_68;
  wire  T_702;
  wire  T_703;
  wire [4:0] GEN_69;
  wire [4:0] GEN_70;
  wire [4:0] GEN_71;
  wire [4:0] GEN_72;
  wire [4:0] T_705;
  wire [4:0] GEN_73;
  wire [4:0] GEN_74;
  wire [4:0] GEN_75;
  wire [4:0] GEN_76;
  wire [2:0] T_706;
  wire  T_708;
  wire [2:0] ex_rm;
  wire [64:0] cp_rs2;
  wire [64:0] cp_rs3;
  wire [4:0] req_cmd;
  wire  req_ldst;
  wire  req_wen;
  wire  req_ren1;
  wire  req_ren2;
  wire  req_ren3;
  wire  req_swap12;
  wire  req_swap23;
  wire  req_single;
  wire  req_fromint;
  wire  req_toint;
  wire  req_fastpipe;
  wire  req_fma;
  wire  req_div;
  wire  req_sqrt;
  wire  req_round;
  wire  req_wflags;
  wire [2:0] req_rm;
  wire [1:0] req_typ;
  wire [64:0] req_in1;
  wire [64:0] req_in2;
  wire [64:0] req_in3;
  wire [2:0] T_755;
  wire [64:0] T_756;
  wire [64:0] T_757;
  wire [64:0] T_758;
  wire [1:0] T_759;
  wire [1:0] T_760;
  wire  sfma_clk;
  wire  sfma_reset;
  wire  sfma_io_in_valid;
  wire [4:0] sfma_io_in_bits_cmd;
  wire  sfma_io_in_bits_ldst;
  wire  sfma_io_in_bits_wen;
  wire  sfma_io_in_bits_ren1;
  wire  sfma_io_in_bits_ren2;
  wire  sfma_io_in_bits_ren3;
  wire  sfma_io_in_bits_swap12;
  wire  sfma_io_in_bits_swap23;
  wire  sfma_io_in_bits_single;
  wire  sfma_io_in_bits_fromint;
  wire  sfma_io_in_bits_toint;
  wire  sfma_io_in_bits_fastpipe;
  wire  sfma_io_in_bits_fma;
  wire  sfma_io_in_bits_div;
  wire  sfma_io_in_bits_sqrt;
  wire  sfma_io_in_bits_round;
  wire  sfma_io_in_bits_wflags;
  wire [2:0] sfma_io_in_bits_rm;
  wire [1:0] sfma_io_in_bits_typ;
  wire [64:0] sfma_io_in_bits_in1;
  wire [64:0] sfma_io_in_bits_in2;
  wire [64:0] sfma_io_in_bits_in3;
  wire  sfma_io_out_valid;
  wire [64:0] sfma_io_out_bits_data;
  wire [4:0] sfma_io_out_bits_exc;
  wire  T_761;
  wire  T_762;
  wire  dfma_clk;
  wire  dfma_reset;
  wire  dfma_io_in_valid;
  wire [4:0] dfma_io_in_bits_cmd;
  wire  dfma_io_in_bits_ldst;
  wire  dfma_io_in_bits_wen;
  wire  dfma_io_in_bits_ren1;
  wire  dfma_io_in_bits_ren2;
  wire  dfma_io_in_bits_ren3;
  wire  dfma_io_in_bits_swap12;
  wire  dfma_io_in_bits_swap23;
  wire  dfma_io_in_bits_single;
  wire  dfma_io_in_bits_fromint;
  wire  dfma_io_in_bits_toint;
  wire  dfma_io_in_bits_fastpipe;
  wire  dfma_io_in_bits_fma;
  wire  dfma_io_in_bits_div;
  wire  dfma_io_in_bits_sqrt;
  wire  dfma_io_in_bits_round;
  wire  dfma_io_in_bits_wflags;
  wire [2:0] dfma_io_in_bits_rm;
  wire [1:0] dfma_io_in_bits_typ;
  wire [64:0] dfma_io_in_bits_in1;
  wire [64:0] dfma_io_in_bits_in2;
  wire [64:0] dfma_io_in_bits_in3;
  wire  dfma_io_out_valid;
  wire [64:0] dfma_io_out_bits_data;
  wire [4:0] dfma_io_out_bits_exc;
  wire  T_765;
  wire  T_766;
  wire  fpiu_clk;
  wire  fpiu_reset;
  wire  fpiu_io_in_valid;
  wire [4:0] fpiu_io_in_bits_cmd;
  wire  fpiu_io_in_bits_ldst;
  wire  fpiu_io_in_bits_wen;
  wire  fpiu_io_in_bits_ren1;
  wire  fpiu_io_in_bits_ren2;
  wire  fpiu_io_in_bits_ren3;
  wire  fpiu_io_in_bits_swap12;
  wire  fpiu_io_in_bits_swap23;
  wire  fpiu_io_in_bits_single;
  wire  fpiu_io_in_bits_fromint;
  wire  fpiu_io_in_bits_toint;
  wire  fpiu_io_in_bits_fastpipe;
  wire  fpiu_io_in_bits_fma;
  wire  fpiu_io_in_bits_div;
  wire  fpiu_io_in_bits_sqrt;
  wire  fpiu_io_in_bits_round;
  wire  fpiu_io_in_bits_wflags;
  wire [2:0] fpiu_io_in_bits_rm;
  wire [1:0] fpiu_io_in_bits_typ;
  wire [64:0] fpiu_io_in_bits_in1;
  wire [64:0] fpiu_io_in_bits_in2;
  wire [64:0] fpiu_io_in_bits_in3;
  wire [4:0] fpiu_io_as_double_cmd;
  wire  fpiu_io_as_double_ldst;
  wire  fpiu_io_as_double_wen;
  wire  fpiu_io_as_double_ren1;
  wire  fpiu_io_as_double_ren2;
  wire  fpiu_io_as_double_ren3;
  wire  fpiu_io_as_double_swap12;
  wire  fpiu_io_as_double_swap23;
  wire  fpiu_io_as_double_single;
  wire  fpiu_io_as_double_fromint;
  wire  fpiu_io_as_double_toint;
  wire  fpiu_io_as_double_fastpipe;
  wire  fpiu_io_as_double_fma;
  wire  fpiu_io_as_double_div;
  wire  fpiu_io_as_double_sqrt;
  wire  fpiu_io_as_double_round;
  wire  fpiu_io_as_double_wflags;
  wire [2:0] fpiu_io_as_double_rm;
  wire [1:0] fpiu_io_as_double_typ;
  wire [64:0] fpiu_io_as_double_in1;
  wire [64:0] fpiu_io_as_double_in2;
  wire [64:0] fpiu_io_as_double_in3;
  wire  fpiu_io_out_valid;
  wire  fpiu_io_out_bits_lt;
  wire [63:0] fpiu_io_out_bits_store;
  wire [63:0] fpiu_io_out_bits_toint;
  wire [4:0] fpiu_io_out_bits_exc;
  wire  T_767;
  wire  T_768;
  wire [4:0] GEN_135;
  wire [4:0] T_771;
  wire [4:0] GEN_136;
  wire  T_772;
  wire  T_773;
  wire  T_774;
  wire  T_775;
  wire  T_776;
  wire [63:0] GEN_77;
  wire  ifpu_clk;
  wire  ifpu_reset;
  wire  ifpu_io_in_valid;
  wire [4:0] ifpu_io_in_bits_cmd;
  wire  ifpu_io_in_bits_ldst;
  wire  ifpu_io_in_bits_wen;
  wire  ifpu_io_in_bits_ren1;
  wire  ifpu_io_in_bits_ren2;
  wire  ifpu_io_in_bits_ren3;
  wire  ifpu_io_in_bits_swap12;
  wire  ifpu_io_in_bits_swap23;
  wire  ifpu_io_in_bits_single;
  wire  ifpu_io_in_bits_fromint;
  wire  ifpu_io_in_bits_toint;
  wire  ifpu_io_in_bits_fastpipe;
  wire  ifpu_io_in_bits_fma;
  wire  ifpu_io_in_bits_div;
  wire  ifpu_io_in_bits_sqrt;
  wire  ifpu_io_in_bits_round;
  wire  ifpu_io_in_bits_wflags;
  wire [2:0] ifpu_io_in_bits_rm;
  wire [1:0] ifpu_io_in_bits_typ;
  wire [64:0] ifpu_io_in_bits_in1;
  wire [64:0] ifpu_io_in_bits_in2;
  wire [64:0] ifpu_io_in_bits_in3;
  wire  ifpu_io_out_valid;
  wire [64:0] ifpu_io_out_bits_data;
  wire [4:0] ifpu_io_out_bits_exc;
  wire  T_778;
  wire [64:0] T_779;
  wire  fpmu_clk;
  wire  fpmu_reset;
  wire  fpmu_io_in_valid;
  wire [4:0] fpmu_io_in_bits_cmd;
  wire  fpmu_io_in_bits_ldst;
  wire  fpmu_io_in_bits_wen;
  wire  fpmu_io_in_bits_ren1;
  wire  fpmu_io_in_bits_ren2;
  wire  fpmu_io_in_bits_ren3;
  wire  fpmu_io_in_bits_swap12;
  wire  fpmu_io_in_bits_swap23;
  wire  fpmu_io_in_bits_single;
  wire  fpmu_io_in_bits_fromint;
  wire  fpmu_io_in_bits_toint;
  wire  fpmu_io_in_bits_fastpipe;
  wire  fpmu_io_in_bits_fma;
  wire  fpmu_io_in_bits_div;
  wire  fpmu_io_in_bits_sqrt;
  wire  fpmu_io_in_bits_round;
  wire  fpmu_io_in_bits_wflags;
  wire [2:0] fpmu_io_in_bits_rm;
  wire [1:0] fpmu_io_in_bits_typ;
  wire [64:0] fpmu_io_in_bits_in1;
  wire [64:0] fpmu_io_in_bits_in2;
  wire [64:0] fpmu_io_in_bits_in3;
  wire  fpmu_io_out_valid;
  wire [64:0] fpmu_io_out_bits_data;
  wire [4:0] fpmu_io_out_bits_exc;
  wire  fpmu_io_lt;
  wire  T_780;
  reg  divSqrt_wen;
  reg [31:0] GEN_207;
  wire  divSqrt_inReady;
  reg [4:0] divSqrt_waddr;
  reg [31:0] GEN_208;
  wire [64:0] divSqrt_wdata;
  wire [4:0] divSqrt_flags;
  reg  divSqrt_in_flight;
  reg [31:0] GEN_209;
  reg  divSqrt_killed;
  reg [31:0] GEN_210;
  wire [1:0] T_793;
  wire  T_794;
  wire  T_799;
  wire  T_800;
  wire [1:0] T_803;
  wire [1:0] GEN_137;
  wire [1:0] T_804;
  wire [1:0] GEN_138;
  wire [1:0] T_805;
  wire [1:0] memLatencyMask;
  reg [1:0] wen;
  reg [31:0] GEN_211;
  reg [8:0] winfo_0;
  reg [31:0] GEN_212;
  reg [8:0] winfo_1;
  reg [31:0] GEN_213;
  wire  T_814;
  wire  T_815;
  wire  mem_wen;
  wire [1:0] T_818;
  wire [2:0] T_821;
  wire  T_822;
  wire [1:0] T_825;
  wire  T_828;
  wire [2:0] T_831;
  wire [2:0] GEN_139;
  wire [2:0] T_832;
  wire [2:0] GEN_140;
  wire [2:0] T_833;
  wire [2:0] T_834;
  wire [2:0] GEN_141;
  wire [2:0] T_835;
  wire [2:0] GEN_142;
  wire  T_837;
  wire  T_838;
  wire [2:0] T_841;
  wire [3:0] T_844;
  wire [2:0] T_848;
  wire [3:0] T_854;
  wire [3:0] GEN_143;
  wire [3:0] T_855;
  wire [3:0] GEN_144;
  wire [3:0] T_856;
  wire [3:0] T_857;
  wire [3:0] GEN_145;
  wire [3:0] T_858;
  wire [3:0] GEN_146;
  wire  T_860;
  wire  T_861;
  reg  write_port_busy;
  reg [31:0] GEN_214;
  wire  GEN_79;
  wire [1:0] T_871;
  wire [1:0] T_877;
  wire [1:0] GEN_147;
  wire [1:0] T_879;
  wire [1:0] T_880;
  wire [4:0] T_881;
  wire [5:0] T_882;
  wire [2:0] T_883;
  wire [8:0] mem_winfo;
  wire  T_884;
  wire [8:0] GEN_80;
  wire  T_885;
  wire [1:0] GEN_148;
  wire [1:0] T_889;
  wire [1:0] GEN_81;
  wire  T_891;
  wire  T_892;
  wire  T_893;
  wire [8:0] GEN_82;
  wire  T_896;
  wire  T_897;
  wire [8:0] GEN_83;
  wire [1:0] GEN_84;
  wire [8:0] GEN_85;
  wire [8:0] GEN_86;
  wire [4:0] T_898;
  wire [4:0] waddr;
  wire [2:0] T_899;
  wire [1:0] wsrc;
  wire  wcp;
  wire [64:0] T_905_0;
  wire [64:0] T_905_1;
  wire [64:0] T_905_2;
  wire [64:0] T_905_3;
  wire [64:0] GEN_0;
  wire [1:0] GEN_149;
  wire [64:0] GEN_87;
  wire [64:0] GEN_88;
  wire [64:0] GEN_89;
  wire [64:0] wdata;
  wire [4:0] T_912_0;
  wire [4:0] T_912_1;
  wire [4:0] T_912_2;
  wire [4:0] T_912_3;
  wire  T_915;
  wire  T_916;
  wire  T_917;
  wire  T_918;
  wire  T_921;
  wire [64:0] GEN_95;
  wire  GEN_96;
  wire  wb_toint_valid;
  reg [4:0] wb_toint_exc;
  reg [31:0] GEN_215;
  wire [4:0] GEN_97;
  wire  T_925;
  wire  T_927;
  wire [4:0] T_929;
  wire [4:0] T_931;
  wire [4:0] T_932;
  wire [4:0] GEN_1;
  wire [4:0] GEN_98;
  wire [4:0] GEN_99;
  wire [4:0] GEN_100;
  wire [4:0] T_935;
  wire [4:0] T_936;
  wire  T_937;
  wire  T_938;
  wire  T_940;
  wire [1:0] GEN_151;
  wire  T_942;
  wire  T_943;
  wire  units_busy;
  wire  T_944;
  wire  T_945;
  wire  T_946;
  wire  T_948;
  wire  T_951;
  wire  T_952;
  wire  T_954;
  wire  T_955;
  wire  T_956;
  wire  T_958;
  wire  T_959;
  reg  T_963;
  reg [31:0] GEN_216;
  wire  T_964;
  wire  T_971;
  wire  T_972;
  wire  T_973;
  reg  T_977;
  reg [31:0] GEN_217;
  reg [1:0] T_979;
  reg [31:0] GEN_218;
  reg [4:0] T_981;
  reg [31:0] GEN_219;
  reg [64:0] T_983;
  reg [95:0] GEN_220;
  wire  DivSqrtRecF64_984_clk;
  wire  DivSqrtRecF64_984_reset;
  wire  DivSqrtRecF64_984_io_inReady_div;
  wire  DivSqrtRecF64_984_io_inReady_sqrt;
  wire  DivSqrtRecF64_984_io_inValid;
  wire  DivSqrtRecF64_984_io_sqrtOp;
  wire [64:0] DivSqrtRecF64_984_io_a;
  wire [64:0] DivSqrtRecF64_984_io_b;
  wire [1:0] DivSqrtRecF64_984_io_roundingMode;
  wire  DivSqrtRecF64_984_io_outValid_div;
  wire  DivSqrtRecF64_984_io_outValid_sqrt;
  wire [64:0] DivSqrtRecF64_984_io_out;
  wire [4:0] DivSqrtRecF64_984_io_exceptionFlags;
  wire  T_985;
  wire  T_986;
  wire  T_990;
  wire  T_991;
  wire  T_992;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire [4:0] GEN_104;
  wire [1:0] GEN_105;
  wire  T_996;
  wire  GEN_106;
  wire [64:0] GEN_107;
  wire  GEN_108;
  wire [4:0] GEN_109;
  wire  RecFNToRecFN_99_998_clk;
  wire  RecFNToRecFN_99_998_reset;
  wire [64:0] RecFNToRecFN_99_998_io_in;
  wire [1:0] RecFNToRecFN_99_998_io_roundingMode;
  wire [32:0] RecFNToRecFN_99_998_io_out;
  wire [4:0] RecFNToRecFN_99_998_io_exceptionFlags;
  wire [64:0] T_999;
  wire [4:0] T_1001;
  wire [4:0] T_1002;
  reg [4:0] GEN_58;
  reg [31:0] GEN_221;
  FPUDecoder fp_decoder (
    .clk(fp_decoder_clk),
    .reset(fp_decoder_reset),
    .io_inst(fp_decoder_io_inst),
    .io_sigs_cmd(fp_decoder_io_sigs_cmd),
    .io_sigs_ldst(fp_decoder_io_sigs_ldst),
    .io_sigs_wen(fp_decoder_io_sigs_wen),
    .io_sigs_ren1(fp_decoder_io_sigs_ren1),
    .io_sigs_ren2(fp_decoder_io_sigs_ren2),
    .io_sigs_ren3(fp_decoder_io_sigs_ren3),
    .io_sigs_swap12(fp_decoder_io_sigs_swap12),
    .io_sigs_swap23(fp_decoder_io_sigs_swap23),
    .io_sigs_single(fp_decoder_io_sigs_single),
    .io_sigs_fromint(fp_decoder_io_sigs_fromint),
    .io_sigs_toint(fp_decoder_io_sigs_toint),
    .io_sigs_fastpipe(fp_decoder_io_sigs_fastpipe),
    .io_sigs_fma(fp_decoder_io_sigs_fma),
    .io_sigs_div(fp_decoder_io_sigs_div),
    .io_sigs_sqrt(fp_decoder_io_sigs_sqrt),
    .io_sigs_round(fp_decoder_io_sigs_round),
    .io_sigs_wflags(fp_decoder_io_sigs_wflags)
  );
  FPUFMAPipe sfma (
    .clk(sfma_clk),
    .reset(sfma_reset),
    .io_in_valid(sfma_io_in_valid),
    .io_in_bits_cmd(sfma_io_in_bits_cmd),
    .io_in_bits_ldst(sfma_io_in_bits_ldst),
    .io_in_bits_wen(sfma_io_in_bits_wen),
    .io_in_bits_ren1(sfma_io_in_bits_ren1),
    .io_in_bits_ren2(sfma_io_in_bits_ren2),
    .io_in_bits_ren3(sfma_io_in_bits_ren3),
    .io_in_bits_swap12(sfma_io_in_bits_swap12),
    .io_in_bits_swap23(sfma_io_in_bits_swap23),
    .io_in_bits_single(sfma_io_in_bits_single),
    .io_in_bits_fromint(sfma_io_in_bits_fromint),
    .io_in_bits_toint(sfma_io_in_bits_toint),
    .io_in_bits_fastpipe(sfma_io_in_bits_fastpipe),
    .io_in_bits_fma(sfma_io_in_bits_fma),
    .io_in_bits_div(sfma_io_in_bits_div),
    .io_in_bits_sqrt(sfma_io_in_bits_sqrt),
    .io_in_bits_round(sfma_io_in_bits_round),
    .io_in_bits_wflags(sfma_io_in_bits_wflags),
    .io_in_bits_rm(sfma_io_in_bits_rm),
    .io_in_bits_typ(sfma_io_in_bits_typ),
    .io_in_bits_in1(sfma_io_in_bits_in1),
    .io_in_bits_in2(sfma_io_in_bits_in2),
    .io_in_bits_in3(sfma_io_in_bits_in3),
    .io_out_valid(sfma_io_out_valid),
    .io_out_bits_data(sfma_io_out_bits_data),
    .io_out_bits_exc(sfma_io_out_bits_exc)
  );
  FPUFMAPipe_90 dfma (
    .clk(dfma_clk),
    .reset(dfma_reset),
    .io_in_valid(dfma_io_in_valid),
    .io_in_bits_cmd(dfma_io_in_bits_cmd),
    .io_in_bits_ldst(dfma_io_in_bits_ldst),
    .io_in_bits_wen(dfma_io_in_bits_wen),
    .io_in_bits_ren1(dfma_io_in_bits_ren1),
    .io_in_bits_ren2(dfma_io_in_bits_ren2),
    .io_in_bits_ren3(dfma_io_in_bits_ren3),
    .io_in_bits_swap12(dfma_io_in_bits_swap12),
    .io_in_bits_swap23(dfma_io_in_bits_swap23),
    .io_in_bits_single(dfma_io_in_bits_single),
    .io_in_bits_fromint(dfma_io_in_bits_fromint),
    .io_in_bits_toint(dfma_io_in_bits_toint),
    .io_in_bits_fastpipe(dfma_io_in_bits_fastpipe),
    .io_in_bits_fma(dfma_io_in_bits_fma),
    .io_in_bits_div(dfma_io_in_bits_div),
    .io_in_bits_sqrt(dfma_io_in_bits_sqrt),
    .io_in_bits_round(dfma_io_in_bits_round),
    .io_in_bits_wflags(dfma_io_in_bits_wflags),
    .io_in_bits_rm(dfma_io_in_bits_rm),
    .io_in_bits_typ(dfma_io_in_bits_typ),
    .io_in_bits_in1(dfma_io_in_bits_in1),
    .io_in_bits_in2(dfma_io_in_bits_in2),
    .io_in_bits_in3(dfma_io_in_bits_in3),
    .io_out_valid(dfma_io_out_valid),
    .io_out_bits_data(dfma_io_out_bits_data),
    .io_out_bits_exc(dfma_io_out_bits_exc)
  );
  FPToInt fpiu (
    .clk(fpiu_clk),
    .reset(fpiu_reset),
    .io_in_valid(fpiu_io_in_valid),
    .io_in_bits_cmd(fpiu_io_in_bits_cmd),
    .io_in_bits_ldst(fpiu_io_in_bits_ldst),
    .io_in_bits_wen(fpiu_io_in_bits_wen),
    .io_in_bits_ren1(fpiu_io_in_bits_ren1),
    .io_in_bits_ren2(fpiu_io_in_bits_ren2),
    .io_in_bits_ren3(fpiu_io_in_bits_ren3),
    .io_in_bits_swap12(fpiu_io_in_bits_swap12),
    .io_in_bits_swap23(fpiu_io_in_bits_swap23),
    .io_in_bits_single(fpiu_io_in_bits_single),
    .io_in_bits_fromint(fpiu_io_in_bits_fromint),
    .io_in_bits_toint(fpiu_io_in_bits_toint),
    .io_in_bits_fastpipe(fpiu_io_in_bits_fastpipe),
    .io_in_bits_fma(fpiu_io_in_bits_fma),
    .io_in_bits_div(fpiu_io_in_bits_div),
    .io_in_bits_sqrt(fpiu_io_in_bits_sqrt),
    .io_in_bits_round(fpiu_io_in_bits_round),
    .io_in_bits_wflags(fpiu_io_in_bits_wflags),
    .io_in_bits_rm(fpiu_io_in_bits_rm),
    .io_in_bits_typ(fpiu_io_in_bits_typ),
    .io_in_bits_in1(fpiu_io_in_bits_in1),
    .io_in_bits_in2(fpiu_io_in_bits_in2),
    .io_in_bits_in3(fpiu_io_in_bits_in3),
    .io_as_double_cmd(fpiu_io_as_double_cmd),
    .io_as_double_ldst(fpiu_io_as_double_ldst),
    .io_as_double_wen(fpiu_io_as_double_wen),
    .io_as_double_ren1(fpiu_io_as_double_ren1),
    .io_as_double_ren2(fpiu_io_as_double_ren2),
    .io_as_double_ren3(fpiu_io_as_double_ren3),
    .io_as_double_swap12(fpiu_io_as_double_swap12),
    .io_as_double_swap23(fpiu_io_as_double_swap23),
    .io_as_double_single(fpiu_io_as_double_single),
    .io_as_double_fromint(fpiu_io_as_double_fromint),
    .io_as_double_toint(fpiu_io_as_double_toint),
    .io_as_double_fastpipe(fpiu_io_as_double_fastpipe),
    .io_as_double_fma(fpiu_io_as_double_fma),
    .io_as_double_div(fpiu_io_as_double_div),
    .io_as_double_sqrt(fpiu_io_as_double_sqrt),
    .io_as_double_round(fpiu_io_as_double_round),
    .io_as_double_wflags(fpiu_io_as_double_wflags),
    .io_as_double_rm(fpiu_io_as_double_rm),
    .io_as_double_typ(fpiu_io_as_double_typ),
    .io_as_double_in1(fpiu_io_as_double_in1),
    .io_as_double_in2(fpiu_io_as_double_in2),
    .io_as_double_in3(fpiu_io_as_double_in3),
    .io_out_valid(fpiu_io_out_valid),
    .io_out_bits_lt(fpiu_io_out_bits_lt),
    .io_out_bits_store(fpiu_io_out_bits_store),
    .io_out_bits_toint(fpiu_io_out_bits_toint),
    .io_out_bits_exc(fpiu_io_out_bits_exc)
  );
  IntToFP ifpu (
    .clk(ifpu_clk),
    .reset(ifpu_reset),
    .io_in_valid(ifpu_io_in_valid),
    .io_in_bits_cmd(ifpu_io_in_bits_cmd),
    .io_in_bits_ldst(ifpu_io_in_bits_ldst),
    .io_in_bits_wen(ifpu_io_in_bits_wen),
    .io_in_bits_ren1(ifpu_io_in_bits_ren1),
    .io_in_bits_ren2(ifpu_io_in_bits_ren2),
    .io_in_bits_ren3(ifpu_io_in_bits_ren3),
    .io_in_bits_swap12(ifpu_io_in_bits_swap12),
    .io_in_bits_swap23(ifpu_io_in_bits_swap23),
    .io_in_bits_single(ifpu_io_in_bits_single),
    .io_in_bits_fromint(ifpu_io_in_bits_fromint),
    .io_in_bits_toint(ifpu_io_in_bits_toint),
    .io_in_bits_fastpipe(ifpu_io_in_bits_fastpipe),
    .io_in_bits_fma(ifpu_io_in_bits_fma),
    .io_in_bits_div(ifpu_io_in_bits_div),
    .io_in_bits_sqrt(ifpu_io_in_bits_sqrt),
    .io_in_bits_round(ifpu_io_in_bits_round),
    .io_in_bits_wflags(ifpu_io_in_bits_wflags),
    .io_in_bits_rm(ifpu_io_in_bits_rm),
    .io_in_bits_typ(ifpu_io_in_bits_typ),
    .io_in_bits_in1(ifpu_io_in_bits_in1),
    .io_in_bits_in2(ifpu_io_in_bits_in2),
    .io_in_bits_in3(ifpu_io_in_bits_in3),
    .io_out_valid(ifpu_io_out_valid),
    .io_out_bits_data(ifpu_io_out_bits_data),
    .io_out_bits_exc(ifpu_io_out_bits_exc)
  );
  FPToFP fpmu (
    .clk(fpmu_clk),
    .reset(fpmu_reset),
    .io_in_valid(fpmu_io_in_valid),
    .io_in_bits_cmd(fpmu_io_in_bits_cmd),
    .io_in_bits_ldst(fpmu_io_in_bits_ldst),
    .io_in_bits_wen(fpmu_io_in_bits_wen),
    .io_in_bits_ren1(fpmu_io_in_bits_ren1),
    .io_in_bits_ren2(fpmu_io_in_bits_ren2),
    .io_in_bits_ren3(fpmu_io_in_bits_ren3),
    .io_in_bits_swap12(fpmu_io_in_bits_swap12),
    .io_in_bits_swap23(fpmu_io_in_bits_swap23),
    .io_in_bits_single(fpmu_io_in_bits_single),
    .io_in_bits_fromint(fpmu_io_in_bits_fromint),
    .io_in_bits_toint(fpmu_io_in_bits_toint),
    .io_in_bits_fastpipe(fpmu_io_in_bits_fastpipe),
    .io_in_bits_fma(fpmu_io_in_bits_fma),
    .io_in_bits_div(fpmu_io_in_bits_div),
    .io_in_bits_sqrt(fpmu_io_in_bits_sqrt),
    .io_in_bits_round(fpmu_io_in_bits_round),
    .io_in_bits_wflags(fpmu_io_in_bits_wflags),
    .io_in_bits_rm(fpmu_io_in_bits_rm),
    .io_in_bits_typ(fpmu_io_in_bits_typ),
    .io_in_bits_in1(fpmu_io_in_bits_in1),
    .io_in_bits_in2(fpmu_io_in_bits_in2),
    .io_in_bits_in3(fpmu_io_in_bits_in3),
    .io_out_valid(fpmu_io_out_valid),
    .io_out_bits_data(fpmu_io_out_bits_data),
    .io_out_bits_exc(fpmu_io_out_bits_exc),
    .io_lt(fpmu_io_lt)
  );
  DivSqrtRecF64 DivSqrtRecF64_984 (
    .clk(DivSqrtRecF64_984_clk),
    .reset(DivSqrtRecF64_984_reset),
    .io_inReady_div(DivSqrtRecF64_984_io_inReady_div),
    .io_inReady_sqrt(DivSqrtRecF64_984_io_inReady_sqrt),
    .io_inValid(DivSqrtRecF64_984_io_inValid),
    .io_sqrtOp(DivSqrtRecF64_984_io_sqrtOp),
    .io_a(DivSqrtRecF64_984_io_a),
    .io_b(DivSqrtRecF64_984_io_b),
    .io_roundingMode(DivSqrtRecF64_984_io_roundingMode),
    .io_outValid_div(DivSqrtRecF64_984_io_outValid_div),
    .io_outValid_sqrt(DivSqrtRecF64_984_io_outValid_sqrt),
    .io_out(DivSqrtRecF64_984_io_out),
    .io_exceptionFlags(DivSqrtRecF64_984_io_exceptionFlags)
  );
  RecFNToRecFN_99 RecFNToRecFN_99_998 (
    .clk(RecFNToRecFN_99_998_clk),
    .reset(RecFNToRecFN_99_998_reset),
    .io_in(RecFNToRecFN_99_998_io_in),
    .io_roundingMode(RecFNToRecFN_99_998_io_roundingMode),
    .io_out(RecFNToRecFN_99_998_io_out),
    .io_exceptionFlags(RecFNToRecFN_99_998_io_exceptionFlags)
  );
  assign io_fcsr_flags_valid = T_927;
  assign io_fcsr_flags_bits = T_936;
  assign io_store_data = fpiu_io_out_bits_store;
  assign io_toint_data = fpiu_io_out_bits_toint;
  assign io_fcsr_rdy = T_954;
  assign io_nack_mem = T_956;
  assign io_illegal_rm = T_973;
  assign io_dec_cmd = fp_decoder_io_sigs_cmd;
  assign io_dec_ldst = fp_decoder_io_sigs_ldst;
  assign io_dec_wen = fp_decoder_io_sigs_wen;
  assign io_dec_ren1 = fp_decoder_io_sigs_ren1;
  assign io_dec_ren2 = fp_decoder_io_sigs_ren2;
  assign io_dec_ren3 = fp_decoder_io_sigs_ren3;
  assign io_dec_swap12 = fp_decoder_io_sigs_swap12;
  assign io_dec_swap23 = fp_decoder_io_sigs_swap23;
  assign io_dec_single = fp_decoder_io_sigs_single;
  assign io_dec_fromint = fp_decoder_io_sigs_fromint;
  assign io_dec_toint = fp_decoder_io_sigs_toint;
  assign io_dec_fastpipe = fp_decoder_io_sigs_fastpipe;
  assign io_dec_fma = fp_decoder_io_sigs_fma;
  assign io_dec_div = fp_decoder_io_sigs_div;
  assign io_dec_sqrt = fp_decoder_io_sigs_sqrt;
  assign io_dec_round = fp_decoder_io_sigs_round;
  assign io_dec_wflags = fp_decoder_io_sigs_wflags;
  assign io_sboard_set = T_964;
  assign io_sboard_clr = T_971;
  assign io_sboard_clra = waddr;
  assign io_cp_req_ready = T_193;
  assign io_cp_resp_valid = GEN_96;
  assign io_cp_resp_bits_data = GEN_95;
  assign io_cp_resp_bits_exc = GEN_58;
  assign req_valid = ex_reg_valid | io_cp_req_valid;
  assign GEN_2 = io_valid ? io_inst : ex_reg_inst;
  assign T_193 = ex_reg_valid == 1'h0;
  assign ex_cp_valid = io_cp_req_valid & T_193;
  assign T_195 = io_killx == 1'h0;
  assign T_196 = ex_reg_valid & T_195;
  assign T_197 = T_196 | ex_cp_valid;
  assign GEN_3 = ex_reg_valid ? ex_reg_inst : mem_reg_inst;
  assign T_200 = io_killm | io_nack_mem;
  assign T_202 = mem_cp_valid == 1'h0;
  assign killm = T_200 & T_202;
  assign T_204 = killm == 1'h0;
  assign T_205 = T_204 | mem_cp_valid;
  assign T_206 = mem_reg_valid & T_205;
  assign fp_decoder_clk = clk;
  assign fp_decoder_reset = reset;
  assign fp_decoder_io_inst = io_inst;
  assign cp_ctrl_cmd = io_cp_req_bits_cmd;
  assign cp_ctrl_ldst = io_cp_req_bits_ldst;
  assign cp_ctrl_wen = io_cp_req_bits_wen;
  assign cp_ctrl_ren1 = io_cp_req_bits_ren1;
  assign cp_ctrl_ren2 = io_cp_req_bits_ren2;
  assign cp_ctrl_ren3 = io_cp_req_bits_ren3;
  assign cp_ctrl_swap12 = io_cp_req_bits_swap12;
  assign cp_ctrl_swap23 = io_cp_req_bits_swap23;
  assign cp_ctrl_single = io_cp_req_bits_single;
  assign cp_ctrl_fromint = io_cp_req_bits_fromint;
  assign cp_ctrl_toint = io_cp_req_bits_toint;
  assign cp_ctrl_fastpipe = io_cp_req_bits_fastpipe;
  assign cp_ctrl_fma = io_cp_req_bits_fma;
  assign cp_ctrl_div = io_cp_req_bits_div;
  assign cp_ctrl_sqrt = io_cp_req_bits_sqrt;
  assign cp_ctrl_round = io_cp_req_bits_round;
  assign cp_ctrl_wflags = io_cp_req_bits_wflags;
  assign GEN_4 = io_valid ? fp_decoder_io_sigs_cmd : T_246_cmd;
  assign GEN_5 = io_valid ? fp_decoder_io_sigs_ldst : T_246_ldst;
  assign GEN_6 = io_valid ? fp_decoder_io_sigs_wen : T_246_wen;
  assign GEN_7 = io_valid ? fp_decoder_io_sigs_ren1 : T_246_ren1;
  assign GEN_8 = io_valid ? fp_decoder_io_sigs_ren2 : T_246_ren2;
  assign GEN_9 = io_valid ? fp_decoder_io_sigs_ren3 : T_246_ren3;
  assign GEN_10 = io_valid ? fp_decoder_io_sigs_swap12 : T_246_swap12;
  assign GEN_11 = io_valid ? fp_decoder_io_sigs_swap23 : T_246_swap23;
  assign GEN_12 = io_valid ? fp_decoder_io_sigs_single : T_246_single;
  assign GEN_13 = io_valid ? fp_decoder_io_sigs_fromint : T_246_fromint;
  assign GEN_14 = io_valid ? fp_decoder_io_sigs_toint : T_246_toint;
  assign GEN_15 = io_valid ? fp_decoder_io_sigs_fastpipe : T_246_fastpipe;
  assign GEN_16 = io_valid ? fp_decoder_io_sigs_fma : T_246_fma;
  assign GEN_17 = io_valid ? fp_decoder_io_sigs_div : T_246_div;
  assign GEN_18 = io_valid ? fp_decoder_io_sigs_sqrt : T_246_sqrt;
  assign GEN_19 = io_valid ? fp_decoder_io_sigs_round : T_246_round;
  assign GEN_20 = io_valid ? fp_decoder_io_sigs_wflags : T_246_wflags;
  assign ex_ctrl_cmd = ex_reg_valid ? T_246_cmd : cp_ctrl_cmd;
  assign ex_ctrl_ldst = ex_reg_valid ? T_246_ldst : cp_ctrl_ldst;
  assign ex_ctrl_wen = ex_reg_valid ? T_246_wen : cp_ctrl_wen;
  assign ex_ctrl_ren1 = ex_reg_valid ? T_246_ren1 : cp_ctrl_ren1;
  assign ex_ctrl_ren2 = ex_reg_valid ? T_246_ren2 : cp_ctrl_ren2;
  assign ex_ctrl_ren3 = ex_reg_valid ? T_246_ren3 : cp_ctrl_ren3;
  assign ex_ctrl_swap12 = ex_reg_valid ? T_246_swap12 : cp_ctrl_swap12;
  assign ex_ctrl_swap23 = ex_reg_valid ? T_246_swap23 : cp_ctrl_swap23;
  assign ex_ctrl_single = ex_reg_valid ? T_246_single : cp_ctrl_single;
  assign ex_ctrl_fromint = ex_reg_valid ? T_246_fromint : cp_ctrl_fromint;
  assign ex_ctrl_toint = ex_reg_valid ? T_246_toint : cp_ctrl_toint;
  assign ex_ctrl_fastpipe = ex_reg_valid ? T_246_fastpipe : cp_ctrl_fastpipe;
  assign ex_ctrl_fma = ex_reg_valid ? T_246_fma : cp_ctrl_fma;
  assign ex_ctrl_div = ex_reg_valid ? T_246_div : cp_ctrl_div;
  assign ex_ctrl_sqrt = ex_reg_valid ? T_246_sqrt : cp_ctrl_sqrt;
  assign ex_ctrl_round = ex_reg_valid ? T_246_round : cp_ctrl_round;
  assign ex_ctrl_wflags = ex_reg_valid ? T_246_wflags : cp_ctrl_wflags;
  assign GEN_21 = req_valid ? ex_ctrl_cmd : mem_ctrl_cmd;
  assign GEN_22 = req_valid ? ex_ctrl_ldst : mem_ctrl_ldst;
  assign GEN_23 = req_valid ? ex_ctrl_wen : mem_ctrl_wen;
  assign GEN_24 = req_valid ? ex_ctrl_ren1 : mem_ctrl_ren1;
  assign GEN_25 = req_valid ? ex_ctrl_ren2 : mem_ctrl_ren2;
  assign GEN_26 = req_valid ? ex_ctrl_ren3 : mem_ctrl_ren3;
  assign GEN_27 = req_valid ? ex_ctrl_swap12 : mem_ctrl_swap12;
  assign GEN_28 = req_valid ? ex_ctrl_swap23 : mem_ctrl_swap23;
  assign GEN_29 = req_valid ? ex_ctrl_single : mem_ctrl_single;
  assign GEN_30 = req_valid ? ex_ctrl_fromint : mem_ctrl_fromint;
  assign GEN_31 = req_valid ? ex_ctrl_toint : mem_ctrl_toint;
  assign GEN_32 = req_valid ? ex_ctrl_fastpipe : mem_ctrl_fastpipe;
  assign GEN_33 = req_valid ? ex_ctrl_fma : mem_ctrl_fma;
  assign GEN_34 = req_valid ? ex_ctrl_div : mem_ctrl_div;
  assign GEN_35 = req_valid ? ex_ctrl_sqrt : mem_ctrl_sqrt;
  assign GEN_36 = req_valid ? ex_ctrl_round : mem_ctrl_round;
  assign GEN_37 = req_valid ? ex_ctrl_wflags : mem_ctrl_wflags;
  assign GEN_38 = mem_reg_valid ? mem_ctrl_cmd : wb_ctrl_cmd;
  assign GEN_39 = mem_reg_valid ? mem_ctrl_ldst : wb_ctrl_ldst;
  assign GEN_40 = mem_reg_valid ? mem_ctrl_wen : wb_ctrl_wen;
  assign GEN_41 = mem_reg_valid ? mem_ctrl_ren1 : wb_ctrl_ren1;
  assign GEN_42 = mem_reg_valid ? mem_ctrl_ren2 : wb_ctrl_ren2;
  assign GEN_43 = mem_reg_valid ? mem_ctrl_ren3 : wb_ctrl_ren3;
  assign GEN_44 = mem_reg_valid ? mem_ctrl_swap12 : wb_ctrl_swap12;
  assign GEN_45 = mem_reg_valid ? mem_ctrl_swap23 : wb_ctrl_swap23;
  assign GEN_46 = mem_reg_valid ? mem_ctrl_single : wb_ctrl_single;
  assign GEN_47 = mem_reg_valid ? mem_ctrl_fromint : wb_ctrl_fromint;
  assign GEN_48 = mem_reg_valid ? mem_ctrl_toint : wb_ctrl_toint;
  assign GEN_49 = mem_reg_valid ? mem_ctrl_fastpipe : wb_ctrl_fastpipe;
  assign GEN_50 = mem_reg_valid ? mem_ctrl_fma : wb_ctrl_fma;
  assign GEN_51 = mem_reg_valid ? mem_ctrl_div : wb_ctrl_div;
  assign GEN_52 = mem_reg_valid ? mem_ctrl_sqrt : wb_ctrl_sqrt;
  assign GEN_53 = mem_reg_valid ? mem_ctrl_round : wb_ctrl_round;
  assign GEN_54 = mem_reg_valid ? mem_ctrl_wflags : wb_ctrl_wflags;
  assign T_315 = io_dmem_resp_type == 3'h2;
  assign T_316 = io_dmem_resp_type == 3'h6;
  assign T_317 = T_315 | T_316;
  assign GEN_55 = io_dmem_resp_val ? T_317 : load_wb_single;
  assign GEN_56 = io_dmem_resp_val ? io_dmem_resp_data : load_wb_data;
  assign GEN_57 = io_dmem_resp_val ? io_dmem_resp_tag : load_wb_tag;
  assign T_318 = load_wb_data[31];
  assign T_319 = load_wb_data[30:23];
  assign T_320 = load_wb_data[22:0];
  assign GEN_110 = {{7'd0}, 1'h0};
  assign T_322 = T_319 == GEN_110;
  assign GEN_111 = {{22'd0}, 1'h0};
  assign T_324 = T_320 == GEN_111;
  assign T_325 = T_322 & T_324;
  assign GEN_112 = {{9'd0}, T_320};
  assign T_326 = GEN_112 << 9;
  assign T_327 = T_326[31];
  assign T_329 = T_326[30];
  assign T_331 = T_326[29];
  assign T_333 = T_326[28];
  assign T_335 = T_326[27];
  assign T_337 = T_326[26];
  assign T_339 = T_326[25];
  assign T_341 = T_326[24];
  assign T_343 = T_326[23];
  assign T_345 = T_326[22];
  assign T_347 = T_326[21];
  assign T_349 = T_326[20];
  assign T_351 = T_326[19];
  assign T_353 = T_326[18];
  assign T_355 = T_326[17];
  assign T_357 = T_326[16];
  assign T_359 = T_326[15];
  assign T_361 = T_326[14];
  assign T_363 = T_326[13];
  assign T_365 = T_326[12];
  assign T_367 = T_326[11];
  assign T_369 = T_326[10];
  assign T_371 = T_326[9];
  assign T_373 = T_326[8];
  assign T_375 = T_326[7];
  assign T_377 = T_326[6];
  assign T_379 = T_326[5];
  assign T_381 = T_326[4];
  assign T_383 = T_326[3];
  assign T_385 = T_326[2];
  assign T_387 = T_326[1];
  assign T_389 = T_385 ? 2'h2 : {{1'd0}, T_387};
  assign T_390 = T_383 ? 2'h3 : T_389;
  assign T_391 = T_381 ? 3'h4 : {{1'd0}, T_390};
  assign T_392 = T_379 ? 3'h5 : T_391;
  assign T_393 = T_377 ? 3'h6 : T_392;
  assign T_394 = T_375 ? 3'h7 : T_393;
  assign T_395 = T_373 ? 4'h8 : {{1'd0}, T_394};
  assign T_396 = T_371 ? 4'h9 : T_395;
  assign T_397 = T_369 ? 4'ha : T_396;
  assign T_398 = T_367 ? 4'hb : T_397;
  assign T_399 = T_365 ? 4'hc : T_398;
  assign T_400 = T_363 ? 4'hd : T_399;
  assign T_401 = T_361 ? 4'he : T_400;
  assign T_402 = T_359 ? 4'hf : T_401;
  assign T_403 = T_357 ? 5'h10 : {{1'd0}, T_402};
  assign T_404 = T_355 ? 5'h11 : T_403;
  assign T_405 = T_353 ? 5'h12 : T_404;
  assign T_406 = T_351 ? 5'h13 : T_405;
  assign T_407 = T_349 ? 5'h14 : T_406;
  assign T_408 = T_347 ? 5'h15 : T_407;
  assign T_409 = T_345 ? 5'h16 : T_408;
  assign T_410 = T_343 ? 5'h17 : T_409;
  assign T_411 = T_341 ? 5'h18 : T_410;
  assign T_412 = T_339 ? 5'h19 : T_411;
  assign T_413 = T_337 ? 5'h1a : T_412;
  assign T_414 = T_335 ? 5'h1b : T_413;
  assign T_415 = T_333 ? 5'h1c : T_414;
  assign T_416 = T_331 ? 5'h1d : T_415;
  assign T_417 = T_329 ? 5'h1e : T_416;
  assign T_418 = T_327 ? 5'h1f : T_417;
  assign T_419 = ~ T_418;
  assign GEN_113 = {{31'd0}, T_320};
  assign T_420 = GEN_113 << T_419;
  assign T_421 = T_420[21:0];
  assign T_423 = {T_421,1'h0};
  assign GEN_114 = {{8'd0}, 1'h1};
  assign T_426 = 9'h0 - GEN_114;
  assign T_427 = T_426[8:0];
  assign GEN_115 = {{4'd0}, T_419};
  assign T_428 = GEN_115 ^ T_427;
  assign T_429 = T_322 ? T_428 : {{1'd0}, T_319};
  assign T_433 = T_322 ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_116 = {{6'd0}, T_433};
  assign T_434 = 8'h80 | GEN_116;
  assign GEN_117 = {{1'd0}, T_434};
  assign T_435 = T_429 + GEN_117;
  assign T_436 = T_435[8:0];
  assign T_437 = T_436[8:7];
  assign T_439 = T_437 == 2'h3;
  assign T_441 = T_324 == 1'h0;
  assign T_442 = T_439 & T_441;
  assign GEN_118 = {{2'd0}, T_325};
  assign T_444 = 3'h0 - GEN_118;
  assign T_445 = T_444[2:0];
  assign GEN_119 = {{6'd0}, T_445};
  assign T_446 = GEN_119 << 6;
  assign T_447 = ~ T_446;
  assign T_448 = T_436 & T_447;
  assign GEN_120 = {{6'd0}, T_442};
  assign T_449 = GEN_120 << 6;
  assign GEN_121 = {{2'd0}, T_449};
  assign T_450 = T_448 | GEN_121;
  assign T_451 = T_322 ? T_423 : T_320;
  assign T_452 = {T_318,T_450};
  assign rec_s = {T_452,T_451};
  assign T_453 = load_wb_data[63];
  assign T_454 = load_wb_data[62:52];
  assign T_455 = load_wb_data[51:0];
  assign GEN_122 = {{10'd0}, 1'h0};
  assign T_457 = T_454 == GEN_122;
  assign GEN_123 = {{51'd0}, 1'h0};
  assign T_459 = T_455 == GEN_123;
  assign T_460 = T_457 & T_459;
  assign GEN_124 = {{12'd0}, T_455};
  assign T_461 = GEN_124 << 12;
  assign T_462 = T_461[63];
  assign T_464 = T_461[62];
  assign T_466 = T_461[61];
  assign T_468 = T_461[60];
  assign T_470 = T_461[59];
  assign T_472 = T_461[58];
  assign T_474 = T_461[57];
  assign T_476 = T_461[56];
  assign T_478 = T_461[55];
  assign T_480 = T_461[54];
  assign T_482 = T_461[53];
  assign T_484 = T_461[52];
  assign T_486 = T_461[51];
  assign T_488 = T_461[50];
  assign T_490 = T_461[49];
  assign T_492 = T_461[48];
  assign T_494 = T_461[47];
  assign T_496 = T_461[46];
  assign T_498 = T_461[45];
  assign T_500 = T_461[44];
  assign T_502 = T_461[43];
  assign T_504 = T_461[42];
  assign T_506 = T_461[41];
  assign T_508 = T_461[40];
  assign T_510 = T_461[39];
  assign T_512 = T_461[38];
  assign T_514 = T_461[37];
  assign T_516 = T_461[36];
  assign T_518 = T_461[35];
  assign T_520 = T_461[34];
  assign T_522 = T_461[33];
  assign T_524 = T_461[32];
  assign T_526 = T_461[31];
  assign T_528 = T_461[30];
  assign T_530 = T_461[29];
  assign T_532 = T_461[28];
  assign T_534 = T_461[27];
  assign T_536 = T_461[26];
  assign T_538 = T_461[25];
  assign T_540 = T_461[24];
  assign T_542 = T_461[23];
  assign T_544 = T_461[22];
  assign T_546 = T_461[21];
  assign T_548 = T_461[20];
  assign T_550 = T_461[19];
  assign T_552 = T_461[18];
  assign T_554 = T_461[17];
  assign T_556 = T_461[16];
  assign T_558 = T_461[15];
  assign T_560 = T_461[14];
  assign T_562 = T_461[13];
  assign T_564 = T_461[12];
  assign T_566 = T_461[11];
  assign T_568 = T_461[10];
  assign T_570 = T_461[9];
  assign T_572 = T_461[8];
  assign T_574 = T_461[7];
  assign T_576 = T_461[6];
  assign T_578 = T_461[5];
  assign T_580 = T_461[4];
  assign T_582 = T_461[3];
  assign T_584 = T_461[2];
  assign T_586 = T_461[1];
  assign T_588 = T_584 ? 2'h2 : {{1'd0}, T_586};
  assign T_589 = T_582 ? 2'h3 : T_588;
  assign T_590 = T_580 ? 3'h4 : {{1'd0}, T_589};
  assign T_591 = T_578 ? 3'h5 : T_590;
  assign T_592 = T_576 ? 3'h6 : T_591;
  assign T_593 = T_574 ? 3'h7 : T_592;
  assign T_594 = T_572 ? 4'h8 : {{1'd0}, T_593};
  assign T_595 = T_570 ? 4'h9 : T_594;
  assign T_596 = T_568 ? 4'ha : T_595;
  assign T_597 = T_566 ? 4'hb : T_596;
  assign T_598 = T_564 ? 4'hc : T_597;
  assign T_599 = T_562 ? 4'hd : T_598;
  assign T_600 = T_560 ? 4'he : T_599;
  assign T_601 = T_558 ? 4'hf : T_600;
  assign T_602 = T_556 ? 5'h10 : {{1'd0}, T_601};
  assign T_603 = T_554 ? 5'h11 : T_602;
  assign T_604 = T_552 ? 5'h12 : T_603;
  assign T_605 = T_550 ? 5'h13 : T_604;
  assign T_606 = T_548 ? 5'h14 : T_605;
  assign T_607 = T_546 ? 5'h15 : T_606;
  assign T_608 = T_544 ? 5'h16 : T_607;
  assign T_609 = T_542 ? 5'h17 : T_608;
  assign T_610 = T_540 ? 5'h18 : T_609;
  assign T_611 = T_538 ? 5'h19 : T_610;
  assign T_612 = T_536 ? 5'h1a : T_611;
  assign T_613 = T_534 ? 5'h1b : T_612;
  assign T_614 = T_532 ? 5'h1c : T_613;
  assign T_615 = T_530 ? 5'h1d : T_614;
  assign T_616 = T_528 ? 5'h1e : T_615;
  assign T_617 = T_526 ? 5'h1f : T_616;
  assign T_618 = T_524 ? 6'h20 : {{1'd0}, T_617};
  assign T_619 = T_522 ? 6'h21 : T_618;
  assign T_620 = T_520 ? 6'h22 : T_619;
  assign T_621 = T_518 ? 6'h23 : T_620;
  assign T_622 = T_516 ? 6'h24 : T_621;
  assign T_623 = T_514 ? 6'h25 : T_622;
  assign T_624 = T_512 ? 6'h26 : T_623;
  assign T_625 = T_510 ? 6'h27 : T_624;
  assign T_626 = T_508 ? 6'h28 : T_625;
  assign T_627 = T_506 ? 6'h29 : T_626;
  assign T_628 = T_504 ? 6'h2a : T_627;
  assign T_629 = T_502 ? 6'h2b : T_628;
  assign T_630 = T_500 ? 6'h2c : T_629;
  assign T_631 = T_498 ? 6'h2d : T_630;
  assign T_632 = T_496 ? 6'h2e : T_631;
  assign T_633 = T_494 ? 6'h2f : T_632;
  assign T_634 = T_492 ? 6'h30 : T_633;
  assign T_635 = T_490 ? 6'h31 : T_634;
  assign T_636 = T_488 ? 6'h32 : T_635;
  assign T_637 = T_486 ? 6'h33 : T_636;
  assign T_638 = T_484 ? 6'h34 : T_637;
  assign T_639 = T_482 ? 6'h35 : T_638;
  assign T_640 = T_480 ? 6'h36 : T_639;
  assign T_641 = T_478 ? 6'h37 : T_640;
  assign T_642 = T_476 ? 6'h38 : T_641;
  assign T_643 = T_474 ? 6'h39 : T_642;
  assign T_644 = T_472 ? 6'h3a : T_643;
  assign T_645 = T_470 ? 6'h3b : T_644;
  assign T_646 = T_468 ? 6'h3c : T_645;
  assign T_647 = T_466 ? 6'h3d : T_646;
  assign T_648 = T_464 ? 6'h3e : T_647;
  assign T_649 = T_462 ? 6'h3f : T_648;
  assign T_650 = ~ T_649;
  assign GEN_125 = {{63'd0}, T_455};
  assign T_651 = GEN_125 << T_650;
  assign T_652 = T_651[50:0];
  assign T_654 = {T_652,1'h0};
  assign GEN_126 = {{11'd0}, 1'h1};
  assign T_657 = 12'h0 - GEN_126;
  assign T_658 = T_657[11:0];
  assign GEN_127 = {{6'd0}, T_650};
  assign T_659 = GEN_127 ^ T_658;
  assign T_660 = T_457 ? T_659 : {{1'd0}, T_454};
  assign T_664 = T_457 ? 2'h2 : {{1'd0}, 1'h1};
  assign GEN_128 = {{9'd0}, T_664};
  assign T_665 = 11'h400 | GEN_128;
  assign GEN_129 = {{1'd0}, T_665};
  assign T_666 = T_660 + GEN_129;
  assign T_667 = T_666[11:0];
  assign T_668 = T_667[11:10];
  assign T_670 = T_668 == 2'h3;
  assign T_672 = T_459 == 1'h0;
  assign T_673 = T_670 & T_672;
  assign GEN_130 = {{2'd0}, T_460};
  assign T_675 = 3'h0 - GEN_130;
  assign T_676 = T_675[2:0];
  assign GEN_131 = {{9'd0}, T_676};
  assign T_677 = GEN_131 << 9;
  assign T_678 = ~ T_677;
  assign T_679 = T_667 & T_678;
  assign GEN_132 = {{9'd0}, T_673};
  assign T_680 = GEN_132 << 9;
  assign GEN_133 = {{2'd0}, T_680};
  assign T_681 = T_679 | GEN_133;
  assign T_682 = T_457 ? T_654 : T_455;
  assign T_683 = {T_453,T_681};
  assign rec_d = {T_683,T_682};
  assign GEN_134 = $signed(32'hffffffff);
  assign T_685 = $unsigned(GEN_134);
  assign T_686 = {T_685,rec_s};
  assign load_wb_data_recoded = load_wb_single ? T_686 : rec_d;
  assign regfile_ex_rs1_addr = ex_ra1;
  assign regfile_ex_rs1_en = 1'h1;
  `ifdef SYNTHESIS
  assign regfile_ex_rs1_data = regfile[regfile_ex_rs1_addr];
  `else
  assign regfile_ex_rs1_data = regfile_ex_rs1_addr >= 6'h20 ? $random : regfile[regfile_ex_rs1_addr];
  `endif
  assign regfile_ex_rs2_addr = ex_ra2;
  assign regfile_ex_rs2_en = 1'h1;
  `ifdef SYNTHESIS
  assign regfile_ex_rs2_data = regfile[regfile_ex_rs2_addr];
  `else
  assign regfile_ex_rs2_data = regfile_ex_rs2_addr >= 6'h20 ? $random : regfile[regfile_ex_rs2_addr];
  `endif
  assign regfile_ex_rs3_addr = ex_ra3;
  assign regfile_ex_rs3_en = 1'h1;
  `ifdef SYNTHESIS
  assign regfile_ex_rs3_data = regfile[regfile_ex_rs3_addr];
  `else
  assign regfile_ex_rs3_data = regfile_ex_rs3_addr >= 6'h20 ? $random : regfile[regfile_ex_rs3_addr];
  `endif
  assign regfile_T_689_data = load_wb_data_recoded;
  assign regfile_T_689_addr = load_wb_tag;
  assign regfile_T_689_mask = load_wb;
  assign regfile_T_689_en = load_wb;
  assign regfile_T_919_data = wdata;
  assign regfile_T_919_addr = waddr;
  assign regfile_T_919_mask = T_918;
  assign regfile_T_919_en = T_918;
  assign T_694 = fp_decoder_io_sigs_swap12 == 1'h0;
  assign T_695 = io_inst[19:15];
  assign GEN_63 = T_694 ? T_695 : ex_ra1;
  assign GEN_64 = fp_decoder_io_sigs_swap12 ? T_695 : ex_ra2;
  assign GEN_65 = fp_decoder_io_sigs_ren1 ? GEN_63 : ex_ra1;
  assign GEN_66 = fp_decoder_io_sigs_ren1 ? GEN_64 : ex_ra2;
  assign T_697 = io_inst[24:20];
  assign GEN_67 = fp_decoder_io_sigs_swap12 ? T_697 : GEN_65;
  assign GEN_68 = fp_decoder_io_sigs_swap23 ? T_697 : ex_ra3;
  assign T_702 = fp_decoder_io_sigs_swap23 == 1'h0;
  assign T_703 = T_694 & T_702;
  assign GEN_69 = T_703 ? T_697 : GEN_66;
  assign GEN_70 = fp_decoder_io_sigs_ren2 ? GEN_67 : GEN_65;
  assign GEN_71 = fp_decoder_io_sigs_ren2 ? GEN_68 : ex_ra3;
  assign GEN_72 = fp_decoder_io_sigs_ren2 ? GEN_69 : GEN_66;
  assign T_705 = io_inst[31:27];
  assign GEN_73 = fp_decoder_io_sigs_ren3 ? T_705 : GEN_71;
  assign GEN_74 = io_valid ? GEN_70 : ex_ra1;
  assign GEN_75 = io_valid ? GEN_72 : ex_ra2;
  assign GEN_76 = io_valid ? GEN_73 : ex_ra3;
  assign T_706 = ex_reg_inst[14:12];
  assign T_708 = T_706 == 3'h7;
  assign ex_rm = T_708 ? io_fcsr_rm : T_706;
  assign cp_rs2 = io_cp_req_bits_swap23 ? io_cp_req_bits_in3 : io_cp_req_bits_in2;
  assign cp_rs3 = io_cp_req_bits_swap23 ? io_cp_req_bits_in2 : io_cp_req_bits_in3;
  assign req_cmd = ex_ctrl_cmd;
  assign req_ldst = ex_ctrl_ldst;
  assign req_wen = ex_ctrl_wen;
  assign req_ren1 = ex_ctrl_ren1;
  assign req_ren2 = ex_ctrl_ren2;
  assign req_ren3 = ex_ctrl_ren3;
  assign req_swap12 = ex_ctrl_swap12;
  assign req_swap23 = ex_ctrl_swap23;
  assign req_single = ex_ctrl_single;
  assign req_fromint = ex_ctrl_fromint;
  assign req_toint = ex_ctrl_toint;
  assign req_fastpipe = ex_ctrl_fastpipe;
  assign req_fma = ex_ctrl_fma;
  assign req_div = ex_ctrl_div;
  assign req_sqrt = ex_ctrl_sqrt;
  assign req_round = ex_ctrl_round;
  assign req_wflags = ex_ctrl_wflags;
  assign req_rm = T_755;
  assign req_typ = T_760;
  assign req_in1 = T_756;
  assign req_in2 = T_757;
  assign req_in3 = T_758;
  assign T_755 = ex_reg_valid ? ex_rm : io_cp_req_bits_rm;
  assign T_756 = ex_reg_valid ? regfile_ex_rs1_data : io_cp_req_bits_in1;
  assign T_757 = ex_reg_valid ? regfile_ex_rs2_data : cp_rs2;
  assign T_758 = ex_reg_valid ? regfile_ex_rs3_data : cp_rs3;
  assign T_759 = ex_reg_inst[21:20];
  assign T_760 = ex_reg_valid ? T_759 : io_cp_req_bits_typ;
  assign sfma_clk = clk;
  assign sfma_reset = reset;
  assign sfma_io_in_valid = T_762;
  assign sfma_io_in_bits_cmd = req_cmd;
  assign sfma_io_in_bits_ldst = req_ldst;
  assign sfma_io_in_bits_wen = req_wen;
  assign sfma_io_in_bits_ren1 = req_ren1;
  assign sfma_io_in_bits_ren2 = req_ren2;
  assign sfma_io_in_bits_ren3 = req_ren3;
  assign sfma_io_in_bits_swap12 = req_swap12;
  assign sfma_io_in_bits_swap23 = req_swap23;
  assign sfma_io_in_bits_single = req_single;
  assign sfma_io_in_bits_fromint = req_fromint;
  assign sfma_io_in_bits_toint = req_toint;
  assign sfma_io_in_bits_fastpipe = req_fastpipe;
  assign sfma_io_in_bits_fma = req_fma;
  assign sfma_io_in_bits_div = req_div;
  assign sfma_io_in_bits_sqrt = req_sqrt;
  assign sfma_io_in_bits_round = req_round;
  assign sfma_io_in_bits_wflags = req_wflags;
  assign sfma_io_in_bits_rm = req_rm;
  assign sfma_io_in_bits_typ = req_typ;
  assign sfma_io_in_bits_in1 = req_in1;
  assign sfma_io_in_bits_in2 = req_in2;
  assign sfma_io_in_bits_in3 = req_in3;
  assign T_761 = req_valid & ex_ctrl_fma;
  assign T_762 = T_761 & ex_ctrl_single;
  assign dfma_clk = clk;
  assign dfma_reset = reset;
  assign dfma_io_in_valid = T_766;
  assign dfma_io_in_bits_cmd = req_cmd;
  assign dfma_io_in_bits_ldst = req_ldst;
  assign dfma_io_in_bits_wen = req_wen;
  assign dfma_io_in_bits_ren1 = req_ren1;
  assign dfma_io_in_bits_ren2 = req_ren2;
  assign dfma_io_in_bits_ren3 = req_ren3;
  assign dfma_io_in_bits_swap12 = req_swap12;
  assign dfma_io_in_bits_swap23 = req_swap23;
  assign dfma_io_in_bits_single = req_single;
  assign dfma_io_in_bits_fromint = req_fromint;
  assign dfma_io_in_bits_toint = req_toint;
  assign dfma_io_in_bits_fastpipe = req_fastpipe;
  assign dfma_io_in_bits_fma = req_fma;
  assign dfma_io_in_bits_div = req_div;
  assign dfma_io_in_bits_sqrt = req_sqrt;
  assign dfma_io_in_bits_round = req_round;
  assign dfma_io_in_bits_wflags = req_wflags;
  assign dfma_io_in_bits_rm = req_rm;
  assign dfma_io_in_bits_typ = req_typ;
  assign dfma_io_in_bits_in1 = req_in1;
  assign dfma_io_in_bits_in2 = req_in2;
  assign dfma_io_in_bits_in3 = req_in3;
  assign T_765 = ex_ctrl_single == 1'h0;
  assign T_766 = T_761 & T_765;
  assign fpiu_clk = clk;
  assign fpiu_reset = reset;
  assign fpiu_io_in_valid = T_774;
  assign fpiu_io_in_bits_cmd = req_cmd;
  assign fpiu_io_in_bits_ldst = req_ldst;
  assign fpiu_io_in_bits_wen = req_wen;
  assign fpiu_io_in_bits_ren1 = req_ren1;
  assign fpiu_io_in_bits_ren2 = req_ren2;
  assign fpiu_io_in_bits_ren3 = req_ren3;
  assign fpiu_io_in_bits_swap12 = req_swap12;
  assign fpiu_io_in_bits_swap23 = req_swap23;
  assign fpiu_io_in_bits_single = req_single;
  assign fpiu_io_in_bits_fromint = req_fromint;
  assign fpiu_io_in_bits_toint = req_toint;
  assign fpiu_io_in_bits_fastpipe = req_fastpipe;
  assign fpiu_io_in_bits_fma = req_fma;
  assign fpiu_io_in_bits_div = req_div;
  assign fpiu_io_in_bits_sqrt = req_sqrt;
  assign fpiu_io_in_bits_round = req_round;
  assign fpiu_io_in_bits_wflags = req_wflags;
  assign fpiu_io_in_bits_rm = req_rm;
  assign fpiu_io_in_bits_typ = req_typ;
  assign fpiu_io_in_bits_in1 = req_in1;
  assign fpiu_io_in_bits_in2 = req_in2;
  assign fpiu_io_in_bits_in3 = req_in3;
  assign T_767 = ex_ctrl_toint | ex_ctrl_div;
  assign T_768 = T_767 | ex_ctrl_sqrt;
  assign GEN_135 = {{1'd0}, 4'hd};
  assign T_771 = ex_ctrl_cmd & GEN_135;
  assign GEN_136 = {{2'd0}, 3'h5};
  assign T_772 = GEN_136 == T_771;
  assign T_773 = T_768 | T_772;
  assign T_774 = req_valid & T_773;
  assign T_775 = fpiu_io_out_valid & mem_cp_valid;
  assign T_776 = T_775 & mem_ctrl_toint;
  assign GEN_77 = T_776 ? fpiu_io_out_bits_toint : {{63'd0}, 1'h0};
  assign ifpu_clk = clk;
  assign ifpu_reset = reset;
  assign ifpu_io_in_valid = T_778;
  assign ifpu_io_in_bits_cmd = req_cmd;
  assign ifpu_io_in_bits_ldst = req_ldst;
  assign ifpu_io_in_bits_wen = req_wen;
  assign ifpu_io_in_bits_ren1 = req_ren1;
  assign ifpu_io_in_bits_ren2 = req_ren2;
  assign ifpu_io_in_bits_ren3 = req_ren3;
  assign ifpu_io_in_bits_swap12 = req_swap12;
  assign ifpu_io_in_bits_swap23 = req_swap23;
  assign ifpu_io_in_bits_single = req_single;
  assign ifpu_io_in_bits_fromint = req_fromint;
  assign ifpu_io_in_bits_toint = req_toint;
  assign ifpu_io_in_bits_fastpipe = req_fastpipe;
  assign ifpu_io_in_bits_fma = req_fma;
  assign ifpu_io_in_bits_div = req_div;
  assign ifpu_io_in_bits_sqrt = req_sqrt;
  assign ifpu_io_in_bits_round = req_round;
  assign ifpu_io_in_bits_wflags = req_wflags;
  assign ifpu_io_in_bits_rm = req_rm;
  assign ifpu_io_in_bits_typ = req_typ;
  assign ifpu_io_in_bits_in1 = T_779;
  assign ifpu_io_in_bits_in2 = req_in2;
  assign ifpu_io_in_bits_in3 = req_in3;
  assign T_778 = req_valid & ex_ctrl_fromint;
  assign T_779 = ex_reg_valid ? {{1'd0}, io_fromint_data} : io_cp_req_bits_in1;
  assign fpmu_clk = clk;
  assign fpmu_reset = reset;
  assign fpmu_io_in_valid = T_780;
  assign fpmu_io_in_bits_cmd = req_cmd;
  assign fpmu_io_in_bits_ldst = req_ldst;
  assign fpmu_io_in_bits_wen = req_wen;
  assign fpmu_io_in_bits_ren1 = req_ren1;
  assign fpmu_io_in_bits_ren2 = req_ren2;
  assign fpmu_io_in_bits_ren3 = req_ren3;
  assign fpmu_io_in_bits_swap12 = req_swap12;
  assign fpmu_io_in_bits_swap23 = req_swap23;
  assign fpmu_io_in_bits_single = req_single;
  assign fpmu_io_in_bits_fromint = req_fromint;
  assign fpmu_io_in_bits_toint = req_toint;
  assign fpmu_io_in_bits_fastpipe = req_fastpipe;
  assign fpmu_io_in_bits_fma = req_fma;
  assign fpmu_io_in_bits_div = req_div;
  assign fpmu_io_in_bits_sqrt = req_sqrt;
  assign fpmu_io_in_bits_round = req_round;
  assign fpmu_io_in_bits_wflags = req_wflags;
  assign fpmu_io_in_bits_rm = req_rm;
  assign fpmu_io_in_bits_typ = req_typ;
  assign fpmu_io_in_bits_in1 = req_in1;
  assign fpmu_io_in_bits_in2 = req_in2;
  assign fpmu_io_in_bits_in3 = req_in3;
  assign fpmu_io_lt = fpiu_io_out_bits_lt;
  assign T_780 = req_valid & ex_ctrl_fastpipe;
  assign divSqrt_inReady = T_985;
  assign divSqrt_wdata = T_999;
  assign divSqrt_flags = T_1002;
  assign T_793 = mem_ctrl_fromint ? 2'h2 : {{1'd0}, 1'h0};
  assign T_794 = mem_ctrl_fma & mem_ctrl_single;
  assign T_799 = mem_ctrl_single == 1'h0;
  assign T_800 = mem_ctrl_fma & T_799;
  assign T_803 = T_800 ? 2'h2 : {{1'd0}, 1'h0};
  assign GEN_137 = {{1'd0}, mem_ctrl_fastpipe};
  assign T_804 = GEN_137 | T_793;
  assign GEN_138 = {{1'd0}, T_794};
  assign T_805 = T_804 | GEN_138;
  assign memLatencyMask = T_805 | T_803;
  assign T_814 = mem_ctrl_fma | mem_ctrl_fastpipe;
  assign T_815 = T_814 | mem_ctrl_fromint;
  assign mem_wen = mem_reg_valid & T_815;
  assign T_818 = ex_ctrl_fastpipe ? 2'h2 : {{1'd0}, 1'h0};
  assign T_821 = ex_ctrl_fromint ? 3'h4 : {{2'd0}, 1'h0};
  assign T_822 = ex_ctrl_fma & ex_ctrl_single;
  assign T_825 = T_822 ? 2'h2 : {{1'd0}, 1'h0};
  assign T_828 = ex_ctrl_fma & T_765;
  assign T_831 = T_828 ? 3'h4 : {{2'd0}, 1'h0};
  assign GEN_139 = {{1'd0}, T_818};
  assign T_832 = GEN_139 | T_821;
  assign GEN_140 = {{1'd0}, T_825};
  assign T_833 = T_832 | GEN_140;
  assign T_834 = T_833 | T_831;
  assign GEN_141 = {{1'd0}, memLatencyMask};
  assign T_835 = GEN_141 & T_834;
  assign GEN_142 = {{2'd0}, 1'h0};
  assign T_837 = T_835 != GEN_142;
  assign T_838 = mem_wen & T_837;
  assign T_841 = ex_ctrl_fastpipe ? 3'h4 : {{2'd0}, 1'h0};
  assign T_844 = ex_ctrl_fromint ? 4'h8 : {{3'd0}, 1'h0};
  assign T_848 = T_822 ? 3'h4 : {{2'd0}, 1'h0};
  assign T_854 = T_828 ? 4'h8 : {{3'd0}, 1'h0};
  assign GEN_143 = {{1'd0}, T_841};
  assign T_855 = GEN_143 | T_844;
  assign GEN_144 = {{1'd0}, T_848};
  assign T_856 = T_855 | GEN_144;
  assign T_857 = T_856 | T_854;
  assign GEN_145 = {{2'd0}, wen};
  assign T_858 = GEN_145 & T_857;
  assign GEN_146 = {{3'd0}, 1'h0};
  assign T_860 = T_858 != GEN_146;
  assign T_861 = T_838 | T_860;
  assign GEN_79 = req_valid ? T_861 : write_port_busy;
  assign T_871 = T_794 ? 2'h2 : {{1'd0}, 1'h0};
  assign T_877 = T_800 ? 2'h3 : {{1'd0}, 1'h0};
  assign GEN_147 = {{1'd0}, mem_ctrl_fromint};
  assign T_879 = GEN_147 | T_871;
  assign T_880 = T_879 | T_877;
  assign T_881 = mem_reg_inst[11:7];
  assign T_882 = {mem_ctrl_single,T_881};
  assign T_883 = {mem_cp_valid,T_880};
  assign mem_winfo = {T_883,T_882};
  assign T_884 = wen[1];
  assign GEN_80 = T_884 ? winfo_1 : winfo_0;
  assign T_885 = wen[1:1];
  assign GEN_148 = {{1'd0}, T_885};
  assign T_889 = GEN_148 | memLatencyMask;
  assign GEN_81 = T_204 ? T_889 : {{1'd0}, T_885};
  assign T_891 = write_port_busy == 1'h0;
  assign T_892 = memLatencyMask[0];
  assign T_893 = T_891 & T_892;
  assign GEN_82 = T_893 ? mem_winfo : GEN_80;
  assign T_896 = memLatencyMask[1];
  assign T_897 = T_891 & T_896;
  assign GEN_83 = T_897 ? mem_winfo : winfo_1;
  assign GEN_84 = mem_wen ? GEN_81 : {{1'd0}, T_885};
  assign GEN_85 = mem_wen ? GEN_82 : GEN_80;
  assign GEN_86 = mem_wen ? GEN_83 : winfo_1;
  assign T_898 = winfo_0[4:0];
  assign waddr = divSqrt_wen ? divSqrt_waddr : T_898;
  assign T_899 = winfo_0[8:6];
  assign wsrc = T_899[1:0];
  assign wcp = winfo_0[8];
  assign T_905_0 = fpmu_io_out_bits_data;
  assign T_905_1 = ifpu_io_out_bits_data;
  assign T_905_2 = sfma_io_out_bits_data;
  assign T_905_3 = dfma_io_out_bits_data;
  assign GEN_0 = GEN_89;
  assign GEN_149 = {{1'd0}, 1'h1};
  assign GEN_87 = GEN_149 == wsrc ? T_905_1 : T_905_0;
  assign GEN_88 = 2'h2 == wsrc ? T_905_2 : GEN_87;
  assign GEN_89 = 2'h3 == wsrc ? T_905_3 : GEN_88;
  assign wdata = divSqrt_wen ? divSqrt_wdata : GEN_0;
  assign T_912_0 = fpmu_io_out_bits_exc;
  assign T_912_1 = ifpu_io_out_bits_exc;
  assign T_912_2 = sfma_io_out_bits_exc;
  assign T_912_3 = dfma_io_out_bits_exc;
  assign T_915 = wcp == 1'h0;
  assign T_916 = wen[0];
  assign T_917 = T_915 & T_916;
  assign T_918 = T_917 | divSqrt_wen;
  assign T_921 = wcp & T_916;
  assign GEN_95 = T_921 ? wdata : {{1'd0}, GEN_77};
  assign GEN_96 = T_921 ? 1'h1 : T_776;
  assign wb_toint_valid = wb_reg_valid & wb_ctrl_toint;
  assign GEN_97 = mem_ctrl_toint ? fpiu_io_out_bits_exc : wb_toint_exc;
  assign T_925 = wb_toint_valid | divSqrt_wen;
  assign T_927 = T_925 | T_916;
  assign T_929 = wb_toint_valid ? wb_toint_exc : {{4'd0}, 1'h0};
  assign T_931 = divSqrt_wen ? divSqrt_flags : {{4'd0}, 1'h0};
  assign T_932 = T_929 | T_931;
  assign GEN_1 = GEN_100;
  assign GEN_98 = GEN_149 == wsrc ? T_912_1 : T_912_0;
  assign GEN_99 = 2'h2 == wsrc ? T_912_2 : GEN_98;
  assign GEN_100 = 2'h3 == wsrc ? T_912_3 : GEN_99;
  assign T_935 = T_916 ? GEN_1 : {{4'd0}, 1'h0};
  assign T_936 = T_932 | T_935;
  assign T_937 = mem_ctrl_div | mem_ctrl_sqrt;
  assign T_938 = mem_reg_valid & T_937;
  assign T_940 = divSqrt_inReady == 1'h0;
  assign GEN_151 = {{1'd0}, 1'h0};
  assign T_942 = wen != GEN_151;
  assign T_943 = T_940 | T_942;
  assign units_busy = T_938 & T_943;
  assign T_944 = ex_reg_valid & ex_ctrl_wflags;
  assign T_945 = mem_reg_valid & mem_ctrl_wflags;
  assign T_946 = T_944 | T_945;
  assign T_948 = T_946 | wb_toint_valid;
  assign T_951 = T_948 | T_942;
  assign T_952 = T_951 | divSqrt_in_flight;
  assign T_954 = T_952 == 1'h0;
  assign T_955 = units_busy | write_port_busy;
  assign T_956 = T_955 | divSqrt_in_flight;
  assign T_958 = wb_cp_valid == 1'h0;
  assign T_959 = wb_reg_valid & T_958;
  assign T_964 = T_959 & T_963;
  assign T_971 = T_958 & divSqrt_wen;
  assign T_972 = ex_rm[2];
  assign T_973 = T_972 & ex_ctrl_round;
  assign DivSqrtRecF64_984_clk = clk;
  assign DivSqrtRecF64_984_reset = reset;
  assign DivSqrtRecF64_984_io_inValid = T_991;
  assign DivSqrtRecF64_984_io_sqrtOp = mem_ctrl_sqrt;
  assign DivSqrtRecF64_984_io_a = fpiu_io_as_double_in1;
  assign DivSqrtRecF64_984_io_b = fpiu_io_as_double_in2;
  assign DivSqrtRecF64_984_io_roundingMode = fpiu_io_as_double_rm[1:0];
  assign T_985 = DivSqrtRecF64_984_io_sqrtOp ? DivSqrtRecF64_984_io_inReady_sqrt : DivSqrtRecF64_984_io_inReady_div;
  assign T_986 = DivSqrtRecF64_984_io_outValid_div | DivSqrtRecF64_984_io_outValid_sqrt;
  assign T_990 = divSqrt_in_flight == 1'h0;
  assign T_991 = T_938 & T_990;
  assign T_992 = DivSqrtRecF64_984_io_inValid & divSqrt_inReady;
  assign GEN_101 = T_992 ? 1'h1 : divSqrt_in_flight;
  assign GEN_102 = T_992 ? killm : divSqrt_killed;
  assign GEN_103 = T_992 ? mem_ctrl_single : T_977;
  assign GEN_104 = T_992 ? T_881 : divSqrt_waddr;
  assign GEN_105 = T_992 ? DivSqrtRecF64_984_io_roundingMode : T_979;
  assign T_996 = divSqrt_killed == 1'h0;
  assign GEN_106 = T_986 ? T_996 : 1'h0;
  assign GEN_107 = T_986 ? DivSqrtRecF64_984_io_out : T_983;
  assign GEN_108 = T_986 ? 1'h0 : GEN_101;
  assign GEN_109 = T_986 ? DivSqrtRecF64_984_io_exceptionFlags : T_981;
  assign RecFNToRecFN_99_998_clk = clk;
  assign RecFNToRecFN_99_998_reset = reset;
  assign RecFNToRecFN_99_998_io_in = T_983;
  assign RecFNToRecFN_99_998_io_roundingMode = T_979;
  assign T_999 = T_977 ? {{32'd0}, RecFNToRecFN_99_998_io_out} : T_983;
  assign T_1001 = T_977 ? RecFNToRecFN_99_998_io_exceptionFlags : {{4'd0}, 1'h0};
  assign T_1002 = T_981 | T_1001;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_59 = {1{$random}};
  ex_reg_valid = GEN_59[0:0];
  GEN_60 = {1{$random}};
  ex_reg_inst = GEN_60[31:0];
  GEN_61 = {1{$random}};
  mem_reg_valid = GEN_61[0:0];
  GEN_62 = {1{$random}};
  mem_reg_inst = GEN_62[31:0];
  GEN_78 = {1{$random}};
  mem_cp_valid = GEN_78[0:0];
  GEN_90 = {1{$random}};
  wb_reg_valid = GEN_90[0:0];
  GEN_91 = {1{$random}};
  wb_cp_valid = GEN_91[0:0];
  GEN_92 = {1{$random}};
  T_246_cmd = GEN_92[4:0];
  GEN_93 = {1{$random}};
  T_246_ldst = GEN_93[0:0];
  GEN_94 = {1{$random}};
  T_246_wen = GEN_94[0:0];
  GEN_150 = {1{$random}};
  T_246_ren1 = GEN_150[0:0];
  GEN_152 = {1{$random}};
  T_246_ren2 = GEN_152[0:0];
  GEN_153 = {1{$random}};
  T_246_ren3 = GEN_153[0:0];
  GEN_154 = {1{$random}};
  T_246_swap12 = GEN_154[0:0];
  GEN_155 = {1{$random}};
  T_246_swap23 = GEN_155[0:0];
  GEN_156 = {1{$random}};
  T_246_single = GEN_156[0:0];
  GEN_157 = {1{$random}};
  T_246_fromint = GEN_157[0:0];
  GEN_158 = {1{$random}};
  T_246_toint = GEN_158[0:0];
  GEN_159 = {1{$random}};
  T_246_fastpipe = GEN_159[0:0];
  GEN_160 = {1{$random}};
  T_246_fma = GEN_160[0:0];
  GEN_161 = {1{$random}};
  T_246_div = GEN_161[0:0];
  GEN_162 = {1{$random}};
  T_246_sqrt = GEN_162[0:0];
  GEN_163 = {1{$random}};
  T_246_round = GEN_163[0:0];
  GEN_164 = {1{$random}};
  T_246_wflags = GEN_164[0:0];
  GEN_165 = {1{$random}};
  mem_ctrl_cmd = GEN_165[4:0];
  GEN_166 = {1{$random}};
  mem_ctrl_ldst = GEN_166[0:0];
  GEN_167 = {1{$random}};
  mem_ctrl_wen = GEN_167[0:0];
  GEN_168 = {1{$random}};
  mem_ctrl_ren1 = GEN_168[0:0];
  GEN_169 = {1{$random}};
  mem_ctrl_ren2 = GEN_169[0:0];
  GEN_170 = {1{$random}};
  mem_ctrl_ren3 = GEN_170[0:0];
  GEN_171 = {1{$random}};
  mem_ctrl_swap12 = GEN_171[0:0];
  GEN_172 = {1{$random}};
  mem_ctrl_swap23 = GEN_172[0:0];
  GEN_173 = {1{$random}};
  mem_ctrl_single = GEN_173[0:0];
  GEN_174 = {1{$random}};
  mem_ctrl_fromint = GEN_174[0:0];
  GEN_175 = {1{$random}};
  mem_ctrl_toint = GEN_175[0:0];
  GEN_176 = {1{$random}};
  mem_ctrl_fastpipe = GEN_176[0:0];
  GEN_177 = {1{$random}};
  mem_ctrl_fma = GEN_177[0:0];
  GEN_178 = {1{$random}};
  mem_ctrl_div = GEN_178[0:0];
  GEN_179 = {1{$random}};
  mem_ctrl_sqrt = GEN_179[0:0];
  GEN_180 = {1{$random}};
  mem_ctrl_round = GEN_180[0:0];
  GEN_181 = {1{$random}};
  mem_ctrl_wflags = GEN_181[0:0];
  GEN_182 = {1{$random}};
  wb_ctrl_cmd = GEN_182[4:0];
  GEN_183 = {1{$random}};
  wb_ctrl_ldst = GEN_183[0:0];
  GEN_184 = {1{$random}};
  wb_ctrl_wen = GEN_184[0:0];
  GEN_185 = {1{$random}};
  wb_ctrl_ren1 = GEN_185[0:0];
  GEN_186 = {1{$random}};
  wb_ctrl_ren2 = GEN_186[0:0];
  GEN_187 = {1{$random}};
  wb_ctrl_ren3 = GEN_187[0:0];
  GEN_188 = {1{$random}};
  wb_ctrl_swap12 = GEN_188[0:0];
  GEN_189 = {1{$random}};
  wb_ctrl_swap23 = GEN_189[0:0];
  GEN_190 = {1{$random}};
  wb_ctrl_single = GEN_190[0:0];
  GEN_191 = {1{$random}};
  wb_ctrl_fromint = GEN_191[0:0];
  GEN_192 = {1{$random}};
  wb_ctrl_toint = GEN_192[0:0];
  GEN_193 = {1{$random}};
  wb_ctrl_fastpipe = GEN_193[0:0];
  GEN_194 = {1{$random}};
  wb_ctrl_fma = GEN_194[0:0];
  GEN_195 = {1{$random}};
  wb_ctrl_div = GEN_195[0:0];
  GEN_196 = {1{$random}};
  wb_ctrl_sqrt = GEN_196[0:0];
  GEN_197 = {1{$random}};
  wb_ctrl_round = GEN_197[0:0];
  GEN_198 = {1{$random}};
  wb_ctrl_wflags = GEN_198[0:0];
  GEN_199 = {1{$random}};
  load_wb = GEN_199[0:0];
  GEN_200 = {1{$random}};
  load_wb_single = GEN_200[0:0];
  GEN_201 = {2{$random}};
  load_wb_data = GEN_201[63:0];
  GEN_202 = {1{$random}};
  load_wb_tag = GEN_202[4:0];
  GEN_203 = {3{$random}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = GEN_203[64:0];
  GEN_204 = {1{$random}};
  ex_ra1 = GEN_204[4:0];
  GEN_205 = {1{$random}};
  ex_ra2 = GEN_205[4:0];
  GEN_206 = {1{$random}};
  ex_ra3 = GEN_206[4:0];
  GEN_207 = {1{$random}};
  divSqrt_wen = GEN_207[0:0];
  GEN_208 = {1{$random}};
  divSqrt_waddr = GEN_208[4:0];
  GEN_209 = {1{$random}};
  divSqrt_in_flight = GEN_209[0:0];
  GEN_210 = {1{$random}};
  divSqrt_killed = GEN_210[0:0];
  GEN_211 = {1{$random}};
  wen = GEN_211[1:0];
  GEN_212 = {1{$random}};
  winfo_0 = GEN_212[8:0];
  GEN_213 = {1{$random}};
  winfo_1 = GEN_213[8:0];
  GEN_214 = {1{$random}};
  write_port_busy = GEN_214[0:0];
  GEN_215 = {1{$random}};
  wb_toint_exc = GEN_215[4:0];
  GEN_216 = {1{$random}};
  T_963 = GEN_216[0:0];
  GEN_217 = {1{$random}};
  T_977 = GEN_217[0:0];
  GEN_218 = {1{$random}};
  T_979 = GEN_218[1:0];
  GEN_219 = {1{$random}};
  T_981 = GEN_219[4:0];
  GEN_220 = {3{$random}};
  T_983 = GEN_220[64:0];
  GEN_221 = {1{$random}};
  GEN_58 = GEN_221[4:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      ex_reg_valid <= 1'h0;
    end else begin
      ex_reg_valid <= io_valid;
    end
    if(1'h0) begin
    end else begin
      ex_reg_inst <= GEN_2;
    end
    if(reset) begin
      mem_reg_valid <= 1'h0;
    end else begin
      mem_reg_valid <= T_197;
    end
    if(1'h0) begin
    end else begin
      mem_reg_inst <= GEN_3;
    end
    if(reset) begin
      mem_cp_valid <= 1'h0;
    end else begin
      mem_cp_valid <= ex_cp_valid;
    end
    if(reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= T_206;
    end
    if(reset) begin
      wb_cp_valid <= 1'h0;
    end else begin
      wb_cp_valid <= mem_cp_valid;
    end
    if(1'h0) begin
    end else begin
      T_246_cmd <= GEN_4;
    end
    if(1'h0) begin
    end else begin
      T_246_ldst <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      T_246_wen <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      T_246_ren1 <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      T_246_ren2 <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      T_246_ren3 <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      T_246_swap12 <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      T_246_swap23 <= GEN_11;
    end
    if(1'h0) begin
    end else begin
      T_246_single <= GEN_12;
    end
    if(1'h0) begin
    end else begin
      T_246_fromint <= GEN_13;
    end
    if(1'h0) begin
    end else begin
      T_246_toint <= GEN_14;
    end
    if(1'h0) begin
    end else begin
      T_246_fastpipe <= GEN_15;
    end
    if(1'h0) begin
    end else begin
      T_246_fma <= GEN_16;
    end
    if(1'h0) begin
    end else begin
      T_246_div <= GEN_17;
    end
    if(1'h0) begin
    end else begin
      T_246_sqrt <= GEN_18;
    end
    if(1'h0) begin
    end else begin
      T_246_round <= GEN_19;
    end
    if(1'h0) begin
    end else begin
      T_246_wflags <= GEN_20;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_cmd <= GEN_21;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_ldst <= GEN_22;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_wen <= GEN_23;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_ren1 <= GEN_24;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_ren2 <= GEN_25;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_ren3 <= GEN_26;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_swap12 <= GEN_27;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_swap23 <= GEN_28;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_single <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fromint <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_toint <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fastpipe <= GEN_32;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_fma <= GEN_33;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_div <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_sqrt <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_round <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      mem_ctrl_wflags <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_cmd <= GEN_38;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_ldst <= GEN_39;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_wen <= GEN_40;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_ren1 <= GEN_41;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_ren2 <= GEN_42;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_ren3 <= GEN_43;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_swap12 <= GEN_44;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_swap23 <= GEN_45;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_single <= GEN_46;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fromint <= GEN_47;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_toint <= GEN_48;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fastpipe <= GEN_49;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_fma <= GEN_50;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_div <= GEN_51;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_sqrt <= GEN_52;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_round <= GEN_53;
    end
    if(1'h0) begin
    end else begin
      wb_ctrl_wflags <= GEN_54;
    end
    if(1'h0) begin
    end else begin
      load_wb <= io_dmem_resp_val;
    end
    if(1'h0) begin
    end else begin
      load_wb_single <= GEN_55;
    end
    if(1'h0) begin
    end else begin
      load_wb_data <= GEN_56;
    end
    if(1'h0) begin
    end else begin
      load_wb_tag <= GEN_57;
    end
    if(regfile_T_689_en & regfile_T_689_mask) begin
      regfile[regfile_T_689_addr] <= regfile_T_689_data;
    end
    if(regfile_T_919_en & regfile_T_919_mask) begin
      regfile[regfile_T_919_addr] <= regfile_T_919_data;
    end
    if(1'h0) begin
    end else begin
      ex_ra1 <= GEN_74;
    end
    if(1'h0) begin
    end else begin
      ex_ra2 <= GEN_75;
    end
    if(1'h0) begin
    end else begin
      ex_ra3 <= GEN_76;
    end
    if(1'h0) begin
    end else begin
      divSqrt_wen <= GEN_106;
    end
    if(1'h0) begin
    end else begin
      divSqrt_waddr <= GEN_104;
    end
    if(reset) begin
      divSqrt_in_flight <= 1'h0;
    end else begin
      divSqrt_in_flight <= GEN_108;
    end
    if(1'h0) begin
    end else begin
      divSqrt_killed <= GEN_102;
    end
    if(reset) begin
      wen <= 2'h0;
    end else begin
      wen <= GEN_84;
    end
    if(1'h0) begin
    end else begin
      winfo_0 <= GEN_85;
    end
    if(1'h0) begin
    end else begin
      winfo_1 <= GEN_86;
    end
    if(1'h0) begin
    end else begin
      write_port_busy <= GEN_79;
    end
    if(1'h0) begin
    end else begin
      wb_toint_exc <= GEN_97;
    end
    if(1'h0) begin
    end else begin
      T_963 <= T_937;
    end
    if(1'h0) begin
    end else begin
      T_977 <= GEN_103;
    end
    if(1'h0) begin
    end else begin
      T_979 <= GEN_105;
    end
    if(1'h0) begin
    end else begin
      T_981 <= GEN_109;
    end
    if(1'h0) begin
    end else begin
      T_983 <= GEN_107;
    end
  end
endmodule
module ClientUncachedTileLinkIOArbiter_101(
  input   clk,
  input   reset,
  output  io_in_0_acquire_ready,
  input   io_in_0_acquire_valid,
  input  [25:0] io_in_0_acquire_bits_addr_block,
  input  [1:0] io_in_0_acquire_bits_client_xact_id,
  input  [2:0] io_in_0_acquire_bits_addr_beat,
  input   io_in_0_acquire_bits_is_builtin_type,
  input  [2:0] io_in_0_acquire_bits_a_type,
  input  [11:0] io_in_0_acquire_bits_union,
  input  [63:0] io_in_0_acquire_bits_data,
  input   io_in_0_grant_ready,
  output  io_in_0_grant_valid,
  output [2:0] io_in_0_grant_bits_addr_beat,
  output [1:0] io_in_0_grant_bits_client_xact_id,
  output [2:0] io_in_0_grant_bits_manager_xact_id,
  output  io_in_0_grant_bits_is_builtin_type,
  output [3:0] io_in_0_grant_bits_g_type,
  output [63:0] io_in_0_grant_bits_data,
  input   io_out_acquire_ready,
  output  io_out_acquire_valid,
  output [25:0] io_out_acquire_bits_addr_block,
  output [1:0] io_out_acquire_bits_client_xact_id,
  output [2:0] io_out_acquire_bits_addr_beat,
  output  io_out_acquire_bits_is_builtin_type,
  output [2:0] io_out_acquire_bits_a_type,
  output [11:0] io_out_acquire_bits_union,
  output [63:0] io_out_acquire_bits_data,
  output  io_out_grant_ready,
  input   io_out_grant_valid,
  input  [2:0] io_out_grant_bits_addr_beat,
  input  [1:0] io_out_grant_bits_client_xact_id,
  input  [2:0] io_out_grant_bits_manager_xact_id,
  input   io_out_grant_bits_is_builtin_type,
  input  [3:0] io_out_grant_bits_g_type,
  input  [63:0] io_out_grant_bits_data
);
  assign io_in_0_acquire_ready = io_out_acquire_ready;
  assign io_in_0_grant_valid = io_out_grant_valid;
  assign io_in_0_grant_bits_addr_beat = io_out_grant_bits_addr_beat;
  assign io_in_0_grant_bits_client_xact_id = io_out_grant_bits_client_xact_id;
  assign io_in_0_grant_bits_manager_xact_id = io_out_grant_bits_manager_xact_id;
  assign io_in_0_grant_bits_is_builtin_type = io_out_grant_bits_is_builtin_type;
  assign io_in_0_grant_bits_g_type = io_out_grant_bits_g_type;
  assign io_in_0_grant_bits_data = io_out_grant_bits_data;
  assign io_out_acquire_valid = io_in_0_acquire_valid;
  assign io_out_acquire_bits_addr_block = io_in_0_acquire_bits_addr_block;
  assign io_out_acquire_bits_client_xact_id = io_in_0_acquire_bits_client_xact_id;
  assign io_out_acquire_bits_addr_beat = io_in_0_acquire_bits_addr_beat;
  assign io_out_acquire_bits_is_builtin_type = io_in_0_acquire_bits_is_builtin_type;
  assign io_out_acquire_bits_a_type = io_in_0_acquire_bits_a_type;
  assign io_out_acquire_bits_union = io_in_0_acquire_bits_union;
  assign io_out_acquire_bits_data = io_in_0_acquire_bits_data;
  assign io_out_grant_ready = io_in_0_grant_ready;
endmodule
module RRArbiter(
  input   clk,
  input   reset,
  output  io_in_0_ready,
  input   io_in_0_valid,
  input  [26:0] io_in_0_bits_addr,
  input  [1:0] io_in_0_bits_prv,
  input   io_in_0_bits_store,
  input   io_in_0_bits_fetch,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input  [26:0] io_in_1_bits_addr,
  input  [1:0] io_in_1_bits_prv,
  input   io_in_1_bits_store,
  input   io_in_1_bits_fetch,
  input   io_out_ready,
  output  io_out_valid,
  output [26:0] io_out_bits_addr,
  output [1:0] io_out_bits_prv,
  output  io_out_bits_store,
  output  io_out_bits_fetch,
  output  io_chosen
);
  wire  T_143;
  wire  GEN_0;
  wire  GEN_5;
  wire [26:0] GEN_1;
  wire [26:0] GEN_6;
  wire [1:0] GEN_2;
  wire [1:0] GEN_7;
  wire  GEN_3;
  wire  GEN_8;
  wire  GEN_4;
  wire  GEN_9;
  wire  T_169;
  reg  T_170;
  reg [31:0] GEN_13;
  wire  GEN_10;
  wire  T_173;
  wire  T_175;
  wire  T_178;
  wire  T_182;
  wire  T_184;
  wire  T_188;
  wire  T_189;
  wire  T_190;
  wire  GEN_11;
  wire  GEN_12;
  assign io_in_0_ready = T_189;
  assign io_in_1_ready = T_190;
  assign io_out_valid = GEN_0;
  assign io_out_bits_addr = GEN_1;
  assign io_out_bits_prv = GEN_2;
  assign io_out_bits_store = GEN_3;
  assign io_out_bits_fetch = GEN_4;
  assign io_chosen = T_143;
  assign T_143 = GEN_12;
  assign GEN_0 = GEN_5;
  assign GEN_5 = io_chosen ? io_in_1_valid : io_in_0_valid;
  assign GEN_1 = GEN_6;
  assign GEN_6 = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr;
  assign GEN_2 = GEN_7;
  assign GEN_7 = io_chosen ? io_in_1_bits_prv : io_in_0_bits_prv;
  assign GEN_3 = GEN_8;
  assign GEN_8 = io_chosen ? io_in_1_bits_store : io_in_0_bits_store;
  assign GEN_4 = GEN_9;
  assign GEN_9 = io_chosen ? io_in_1_bits_fetch : io_in_0_bits_fetch;
  assign T_169 = io_out_ready & io_out_valid;
  assign GEN_10 = T_169 ? io_chosen : T_170;
  assign T_173 = 1'h1 > T_170;
  assign T_175 = io_in_1_valid & T_173;
  assign T_178 = T_175 | io_in_0_valid;
  assign T_182 = T_175 == 1'h0;
  assign T_184 = T_178 == 1'h0;
  assign T_188 = T_173 | T_184;
  assign T_189 = T_182 & io_out_ready;
  assign T_190 = T_188 & io_out_ready;
  assign GEN_11 = io_in_0_valid ? 1'h0 : 1'h1;
  assign GEN_12 = T_175 ? 1'h1 : GEN_11;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_13 = {1{$random}};
  T_170 = GEN_13[0:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      T_170 <= GEN_10;
    end
  end
endmodule
module PTW(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [26:0] io_requestor_0_req_bits_addr,
  input  [1:0] io_requestor_0_req_bits_prv,
  input   io_requestor_0_req_bits_store,
  input   io_requestor_0_req_bits_fetch,
  output  io_requestor_0_resp_valid,
  output [19:0] io_requestor_0_resp_bits_pte_ppn,
  output [2:0] io_requestor_0_resp_bits_pte_reserved_for_software,
  output  io_requestor_0_resp_bits_pte_d,
  output  io_requestor_0_resp_bits_pte_r,
  output [3:0] io_requestor_0_resp_bits_pte_typ,
  output  io_requestor_0_resp_bits_pte_v,
  output  io_requestor_0_status_debug,
  output [1:0] io_requestor_0_status_prv,
  output  io_requestor_0_status_sd,
  output [30:0] io_requestor_0_status_zero3,
  output  io_requestor_0_status_sd_rv32,
  output [1:0] io_requestor_0_status_zero2,
  output [4:0] io_requestor_0_status_vm,
  output [4:0] io_requestor_0_status_zero1,
  output  io_requestor_0_status_pum,
  output  io_requestor_0_status_mprv,
  output [1:0] io_requestor_0_status_xs,
  output [1:0] io_requestor_0_status_fs,
  output [1:0] io_requestor_0_status_mpp,
  output [1:0] io_requestor_0_status_hpp,
  output  io_requestor_0_status_spp,
  output  io_requestor_0_status_mpie,
  output  io_requestor_0_status_hpie,
  output  io_requestor_0_status_spie,
  output  io_requestor_0_status_upie,
  output  io_requestor_0_status_mie,
  output  io_requestor_0_status_hie,
  output  io_requestor_0_status_sie,
  output  io_requestor_0_status_uie,
  output  io_requestor_0_invalidate,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [26:0] io_requestor_1_req_bits_addr,
  input  [1:0] io_requestor_1_req_bits_prv,
  input   io_requestor_1_req_bits_store,
  input   io_requestor_1_req_bits_fetch,
  output  io_requestor_1_resp_valid,
  output [19:0] io_requestor_1_resp_bits_pte_ppn,
  output [2:0] io_requestor_1_resp_bits_pte_reserved_for_software,
  output  io_requestor_1_resp_bits_pte_d,
  output  io_requestor_1_resp_bits_pte_r,
  output [3:0] io_requestor_1_resp_bits_pte_typ,
  output  io_requestor_1_resp_bits_pte_v,
  output  io_requestor_1_status_debug,
  output [1:0] io_requestor_1_status_prv,
  output  io_requestor_1_status_sd,
  output [30:0] io_requestor_1_status_zero3,
  output  io_requestor_1_status_sd_rv32,
  output [1:0] io_requestor_1_status_zero2,
  output [4:0] io_requestor_1_status_vm,
  output [4:0] io_requestor_1_status_zero1,
  output  io_requestor_1_status_pum,
  output  io_requestor_1_status_mprv,
  output [1:0] io_requestor_1_status_xs,
  output [1:0] io_requestor_1_status_fs,
  output [1:0] io_requestor_1_status_mpp,
  output [1:0] io_requestor_1_status_hpp,
  output  io_requestor_1_status_spp,
  output  io_requestor_1_status_mpie,
  output  io_requestor_1_status_hpie,
  output  io_requestor_1_status_spie,
  output  io_requestor_1_status_upie,
  output  io_requestor_1_status_mie,
  output  io_requestor_1_status_hie,
  output  io_requestor_1_status_sie,
  output  io_requestor_1_status_uie,
  output  io_requestor_1_invalidate,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [8:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [8:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered,
  input  [19:0] io_dpath_ptbr,
  input   io_dpath_invalidate,
  input   io_dpath_status_debug,
  input  [1:0] io_dpath_status_prv,
  input   io_dpath_status_sd,
  input  [30:0] io_dpath_status_zero3,
  input   io_dpath_status_sd_rv32,
  input  [1:0] io_dpath_status_zero2,
  input  [4:0] io_dpath_status_vm,
  input  [4:0] io_dpath_status_zero1,
  input   io_dpath_status_pum,
  input   io_dpath_status_mprv,
  input  [1:0] io_dpath_status_xs,
  input  [1:0] io_dpath_status_fs,
  input  [1:0] io_dpath_status_mpp,
  input  [1:0] io_dpath_status_hpp,
  input   io_dpath_status_spp,
  input   io_dpath_status_mpie,
  input   io_dpath_status_hpie,
  input   io_dpath_status_spie,
  input   io_dpath_status_upie,
  input   io_dpath_status_mie,
  input   io_dpath_status_hie,
  input   io_dpath_status_sie,
  input   io_dpath_status_uie
);
  reg [2:0] state;
  reg [31:0] GEN_20;
  reg [1:0] count;
  reg [31:0] GEN_21;
  reg [26:0] r_req_addr;
  reg [31:0] GEN_22;
  reg [1:0] r_req_prv;
  reg [31:0] GEN_23;
  reg  r_req_store;
  reg [31:0] GEN_24;
  reg  r_req_fetch;
  reg [31:0] GEN_25;
  reg  r_req_dest;
  reg [31:0] GEN_26;
  reg [19:0] r_pte_ppn;
  reg [31:0] GEN_27;
  reg [2:0] r_pte_reserved_for_software;
  reg [31:0] GEN_28;
  reg  r_pte_d;
  reg [31:0] GEN_41;
  reg  r_pte_r;
  reg [31:0] GEN_42;
  reg [3:0] r_pte_typ;
  reg [31:0] GEN_73;
  reg  r_pte_v;
  reg [31:0] GEN_75;
  wire [8:0] T_1845;
  wire [17:0] T_1847;
  wire [8:0] T_1848;
  wire [8:0] T_1850;
  wire [8:0] T_1856_0;
  wire [8:0] T_1856_1;
  wire [8:0] T_1856_2;
  wire  arb_clk;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [26:0] arb_io_in_0_bits_addr;
  wire [1:0] arb_io_in_0_bits_prv;
  wire  arb_io_in_0_bits_store;
  wire  arb_io_in_0_bits_fetch;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [26:0] arb_io_in_1_bits_addr;
  wire [1:0] arb_io_in_1_bits_prv;
  wire  arb_io_in_1_bits_store;
  wire  arb_io_in_1_bits_fetch;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [26:0] arb_io_out_bits_addr;
  wire [1:0] arb_io_out_bits_prv;
  wire  arb_io_out_bits_store;
  wire  arb_io_out_bits_fetch;
  wire  arb_io_chosen;
  wire  T_1863;
  wire [19:0] pte_ppn;
  wire [2:0] pte_reserved_for_software;
  wire  pte_d;
  wire  pte_r;
  wire [3:0] pte_typ;
  wire  pte_v;
  wire  T_1884;
  wire [3:0] T_1885;
  wire  T_1886;
  wire  T_1887;
  wire [2:0] T_1888;
  wire [19:0] T_1889;
  wire [8:0] GEN_0;
  wire [1:0] GEN_69;
  wire [8:0] GEN_4;
  wire [8:0] GEN_5;
  wire [28:0] T_1890;
  wire [31:0] GEN_70;
  wire [31:0] pte_addr;
  wire  T_1891;
  wire [26:0] GEN_6;
  wire [1:0] GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire  GEN_10;
  wire [19:0] GEN_11;
  reg [2:0] T_1893;
  reg [31:0] GEN_80;
  reg  T_1900_0;
  reg [31:0] GEN_81;
  reg  T_1900_1;
  reg [31:0] GEN_82;
  reg  T_1900_2;
  reg [31:0] GEN_83;
  wire [1:0] T_1902;
  wire [2:0] T_1903;
  reg [31:0] T_1906 [0:2];
  reg [31:0] GEN_84;
  wire [31:0] T_1906_T_1911_data;
  wire [1:0] T_1906_T_1911_addr;
  wire  T_1906_T_1911_en;
  wire [31:0] T_1906_T_1914_data;
  wire [1:0] T_1906_T_1914_addr;
  wire  T_1906_T_1914_en;
  wire [31:0] T_1906_T_1917_data;
  wire [1:0] T_1906_T_1917_addr;
  wire  T_1906_T_1917_en;
  wire [31:0] T_1906_T_1959_data;
  wire [1:0] T_1906_T_1959_addr;
  wire  T_1906_T_1959_mask;
  wire  T_1906_T_1959_en;
  reg [19:0] T_1909 [0:2];
  reg [31:0] GEN_85;
  wire [19:0] T_1909_T_1999_data;
  wire [1:0] T_1909_T_1999_addr;
  wire  T_1909_T_1999_en;
  wire [19:0] T_1909_T_2001_data;
  wire [1:0] T_1909_T_2001_addr;
  wire  T_1909_T_2001_en;
  wire [19:0] T_1909_T_2003_data;
  wire [1:0] T_1909_T_2003_addr;
  wire  T_1909_T_2003_en;
  wire [19:0] T_1909_T_1960_data;
  wire [1:0] T_1909_T_1960_addr;
  wire  T_1909_T_1960_mask;
  wire  T_1909_T_1960_en;
  wire  T_1912;
  wire  T_1915;
  wire  T_1918;
  wire  T_1924_0;
  wire  T_1924_1;
  wire  T_1924_2;
  wire [1:0] T_1926;
  wire [2:0] T_1927;
  wire [2:0] T_1928;
  wire [2:0] GEN_71;
  wire  pte_cache_hit;
  wire [3:0] GEN_72;
  wire  T_1931;
  wire  T_1932;
  wire  T_1933;
  wire  T_1935;
  wire  T_1936;
  wire [2:0] T_1937;
  wire  T_1939;
  wire [2:0] T_1941;
  wire  T_1942;
  wire [1:0] T_1943;
  wire [2:0] T_1944;
  wire  T_1945;
  wire [2:0] T_1946;
  wire [1:0] T_1947;
  wire  T_1949;
  wire  T_1950;
  wire [1:0] T_1955;
  wire [1:0] T_1956;
  wire [1:0] T_1957;
  wire  GEN_1;
  wire [1:0] GEN_74;
  wire  GEN_12;
  wire  GEN_13;
  wire  GEN_14;
  wire  GEN_16;
  wire  GEN_17;
  wire  GEN_18;
  wire  T_1961;
  wire  T_1962;
  wire  T_1963;
  wire [1:0] T_1964;
  wire [1:0] GEN_76;
  wire [1:0] T_1967;
  wire  T_1968;
  wire [1:0] T_1969;
  wire  T_1971;
  wire [3:0] GEN_77;
  wire [3:0] T_1973;
  wire [2:0] T_1974;
  wire [2:0] T_1975;
  wire [2:0] T_1976;
  wire [2:0] T_1978;
  wire [2:0] T_1979;
  wire [1:0] T_1980;
  wire  T_1981;
  wire [5:0] GEN_78;
  wire [5:0] T_1983;
  wire [2:0] T_1984;
  wire [2:0] T_1985;
  wire [2:0] T_1986;
  wire [2:0] T_1988;
  wire [2:0] T_1989;
  wire [2:0] GEN_29;
  wire  T_1991;
  wire  GEN_30;
  wire  GEN_31;
  wire  GEN_32;
  wire  T_1995;
  wire  T_1996;
  wire [19:0] T_2005;
  wire [19:0] T_2007;
  wire [19:0] T_2009;
  wire [19:0] T_2011;
  wire [19:0] T_2012;
  wire [19:0] pte_cache_data;
  wire  T_2013;
  wire [3:0] GEN_79;
  wire  T_2015;
  wire  T_2016;
  wire  T_2017;
  wire  T_2018;
  wire  T_2020;
  wire  T_2021;
  wire  T_2022;
  wire  T_2023;
  wire  T_2027;
  wire  T_2028;
  wire  T_2033;
  wire  T_2034;
  wire  T_2036;
  wire  T_2044;
  wire  T_2051;
  wire  T_2052;
  wire  perm_ok;
  wire  T_2054;
  wire  T_2056;
  wire  T_2057;
  wire  T_2058;
  wire  set_dirty_bit;
  wire  T_2059;
  wire  T_2060;
  wire  T_2062;
  wire  T_2063;
  wire [19:0] GEN_33;
  wire [2:0] GEN_34;
  wire  GEN_35;
  wire  GEN_36;
  wire [3:0] GEN_37;
  wire  GEN_38;
  wire [19:0] T_2079_ppn;
  wire [2:0] T_2079_reserved_for_software;
  wire  T_2079_d;
  wire  T_2079_r;
  wire [3:0] T_2079_typ;
  wire  T_2079_v;
  wire [29:0] T_2087;
  wire  T_2088;
  wire [3:0] T_2089;
  wire  T_2090;
  wire  T_2091;
  wire [2:0] T_2092;
  wire [19:0] T_2093;
  wire [19:0] pte_wdata_ppn;
  wire [2:0] pte_wdata_reserved_for_software;
  wire  pte_wdata_d;
  wire  pte_wdata_r;
  wire [3:0] pte_wdata_typ;
  wire  pte_wdata_v;
  wire  T_2102;
  wire  T_2103;
  wire [4:0] T_2106;
  wire [4:0] T_2107;
  wire [5:0] T_2108;
  wire [22:0] T_2109;
  wire [23:0] T_2110;
  wire [29:0] T_2111;
  wire [27:0] r_resp_ppn;
  wire [9:0] T_2114;
  wire [17:0] T_2115;
  wire [27:0] T_2116;
  wire [18:0] T_2117;
  wire [27:0] T_2119;
  wire [27:0] T_2125_0;
  wire [27:0] T_2125_1;
  wire [27:0] T_2125_2;
  wire  resp_val;
  wire  T_2128;
  wire  T_2129;
  wire [27:0] GEN_2;
  wire [27:0] GEN_39;
  wire [27:0] GEN_40;
  wire  T_2132;
  wire [27:0] GEN_3;
  wire  T_2133;
  wire [2:0] GEN_43;
  wire [2:0] GEN_44;
  wire [1:0] GEN_45;
  wire  T_2135;
  wire  T_2137;
  wire  T_2138;
  wire [2:0] T_2141;
  wire [1:0] T_2142;
  wire  GEN_46;
  wire [2:0] GEN_47;
  wire [1:0] GEN_48;
  wire [19:0] GEN_49;
  wire  T_2144;
  wire  T_2145;
  wire [2:0] GEN_50;
  wire  GEN_51;
  wire [2:0] GEN_52;
  wire [1:0] GEN_53;
  wire [19:0] GEN_54;
  wire  T_2146;
  wire [2:0] GEN_55;
  wire  T_2150;
  wire [2:0] GEN_56;
  wire  T_2156;
  wire [2:0] GEN_57;
  wire [1:0] GEN_58;
  wire [2:0] GEN_59;
  wire [1:0] GEN_60;
  wire [2:0] GEN_61;
  wire [1:0] GEN_62;
  wire  T_2160;
  wire [2:0] GEN_63;
  wire [2:0] GEN_64;
  wire  T_2161;
  wire [2:0] GEN_65;
  wire [2:0] GEN_66;
  wire [2:0] GEN_67;
  wire  T_2162;
  wire [2:0] GEN_68;
  reg [8:0] GEN_15;
  reg [31:0] GEN_86;
  reg [63:0] GEN_19;
  reg [63:0] GEN_87;
  RRArbiter arb (
    .clk(arb_clk),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_prv(arb_io_in_0_bits_prv),
    .io_in_0_bits_store(arb_io_in_0_bits_store),
    .io_in_0_bits_fetch(arb_io_in_0_bits_fetch),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_prv(arb_io_in_1_bits_prv),
    .io_in_1_bits_store(arb_io_in_1_bits_store),
    .io_in_1_bits_fetch(arb_io_in_1_bits_fetch),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_prv(arb_io_out_bits_prv),
    .io_out_bits_store(arb_io_out_bits_store),
    .io_out_bits_fetch(arb_io_out_bits_fetch),
    .io_chosen(arb_io_chosen)
  );
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_0_resp_valid = T_2129;
  assign io_requestor_0_resp_bits_pte_ppn = GEN_2[19:0];
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign io_requestor_0_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign io_requestor_0_status_debug = io_dpath_status_debug;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_pum = io_dpath_status_pum;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_mpp = io_dpath_status_mpp;
  assign io_requestor_0_status_hpp = io_dpath_status_hpp;
  assign io_requestor_0_status_spp = io_dpath_status_spp;
  assign io_requestor_0_status_mpie = io_dpath_status_mpie;
  assign io_requestor_0_status_hpie = io_dpath_status_hpie;
  assign io_requestor_0_status_spie = io_dpath_status_spie;
  assign io_requestor_0_status_upie = io_dpath_status_upie;
  assign io_requestor_0_status_mie = io_dpath_status_mie;
  assign io_requestor_0_status_hie = io_dpath_status_hie;
  assign io_requestor_0_status_sie = io_dpath_status_sie;
  assign io_requestor_0_status_uie = io_dpath_status_uie;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  assign io_requestor_1_resp_valid = T_2132;
  assign io_requestor_1_resp_bits_pte_ppn = GEN_3[19:0];
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_typ = r_pte_typ;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_status_debug = io_dpath_status_debug;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_pum = io_dpath_status_pum;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_mpp = io_dpath_status_mpp;
  assign io_requestor_1_status_hpp = io_dpath_status_hpp;
  assign io_requestor_1_status_spp = io_dpath_status_spp;
  assign io_requestor_1_status_mpie = io_dpath_status_mpie;
  assign io_requestor_1_status_hpie = io_dpath_status_hpie;
  assign io_requestor_1_status_spie = io_dpath_status_spie;
  assign io_requestor_1_status_upie = io_dpath_status_upie;
  assign io_requestor_1_status_mie = io_dpath_status_mie;
  assign io_requestor_1_status_hie = io_dpath_status_hie;
  assign io_requestor_1_status_sie = io_dpath_status_sie;
  assign io_requestor_1_status_uie = io_dpath_status_uie;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_mem_req_valid = GEN_51;
  assign io_mem_req_bits_addr = {{8'd0}, pte_addr};
  assign io_mem_req_bits_tag = GEN_15;
  assign io_mem_req_bits_cmd = T_2106;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_data = GEN_19;
  assign io_mem_s1_kill = 1'h0;
  assign io_mem_s1_data = {{34'd0}, T_2111};
  assign io_mem_invalidate_lr = 1'h0;
  assign T_1845 = r_req_addr[26:18];
  assign T_1847 = r_req_addr[26:9];
  assign T_1848 = T_1847[8:0];
  assign T_1850 = r_req_addr[8:0];
  assign T_1856_0 = T_1845;
  assign T_1856_1 = T_1848;
  assign T_1856_2 = T_1850;
  assign arb_clk = clk;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_requestor_0_req_valid;
  assign arb_io_in_0_bits_addr = io_requestor_0_req_bits_addr;
  assign arb_io_in_0_bits_prv = io_requestor_0_req_bits_prv;
  assign arb_io_in_0_bits_store = io_requestor_0_req_bits_store;
  assign arb_io_in_0_bits_fetch = io_requestor_0_req_bits_fetch;
  assign arb_io_in_1_valid = io_requestor_1_req_valid;
  assign arb_io_in_1_bits_addr = io_requestor_1_req_bits_addr;
  assign arb_io_in_1_bits_prv = io_requestor_1_req_bits_prv;
  assign arb_io_in_1_bits_store = io_requestor_1_req_bits_store;
  assign arb_io_in_1_bits_fetch = io_requestor_1_req_bits_fetch;
  assign arb_io_out_ready = T_1863;
  assign T_1863 = state == 3'h0;
  assign pte_ppn = T_1889;
  assign pte_reserved_for_software = T_1888;
  assign pte_d = T_1887;
  assign pte_r = T_1886;
  assign pte_typ = T_1885;
  assign pte_v = T_1884;
  assign T_1884 = io_mem_resp_bits_data[0];
  assign T_1885 = io_mem_resp_bits_data[4:1];
  assign T_1886 = io_mem_resp_bits_data[5];
  assign T_1887 = io_mem_resp_bits_data[6];
  assign T_1888 = io_mem_resp_bits_data[9:7];
  assign T_1889 = io_mem_resp_bits_data[29:10];
  assign GEN_0 = GEN_5;
  assign GEN_69 = {{1'd0}, 1'h1};
  assign GEN_4 = GEN_69 == count ? T_1856_1 : T_1856_0;
  assign GEN_5 = 2'h2 == count ? T_1856_2 : GEN_4;
  assign T_1890 = {r_pte_ppn,GEN_0};
  assign GEN_70 = {{3'd0}, T_1890};
  assign pte_addr = GEN_70 << 3;
  assign T_1891 = arb_io_out_ready & arb_io_out_valid;
  assign GEN_6 = T_1891 ? arb_io_out_bits_addr : r_req_addr;
  assign GEN_7 = T_1891 ? arb_io_out_bits_prv : r_req_prv;
  assign GEN_8 = T_1891 ? arb_io_out_bits_store : r_req_store;
  assign GEN_9 = T_1891 ? arb_io_out_bits_fetch : r_req_fetch;
  assign GEN_10 = T_1891 ? arb_io_chosen : r_req_dest;
  assign GEN_11 = T_1891 ? io_dpath_ptbr : r_pte_ppn;
  assign T_1902 = {T_1900_2,T_1900_1};
  assign T_1903 = {T_1902,T_1900_0};
  assign T_1906_T_1911_addr = {{1'd0}, 1'h0};
  assign T_1906_T_1911_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1906_T_1911_data = T_1906[T_1906_T_1911_addr];
  `else
  assign T_1906_T_1911_data = T_1906_T_1911_addr >= 2'h3 ? $random : T_1906[T_1906_T_1911_addr];
  `endif
  assign T_1906_T_1914_addr = {{1'd0}, 1'h1};
  assign T_1906_T_1914_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1906_T_1914_data = T_1906[T_1906_T_1914_addr];
  `else
  assign T_1906_T_1914_data = T_1906_T_1914_addr >= 2'h3 ? $random : T_1906[T_1906_T_1914_addr];
  `endif
  assign T_1906_T_1917_addr = 2'h2;
  assign T_1906_T_1917_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1906_T_1917_data = T_1906[T_1906_T_1917_addr];
  `else
  assign T_1906_T_1917_data = T_1906_T_1917_addr >= 2'h3 ? $random : T_1906[T_1906_T_1917_addr];
  `endif
  assign T_1906_T_1959_data = pte_addr;
  assign T_1906_T_1959_addr = T_1957;
  assign T_1906_T_1959_mask = T_1936;
  assign T_1906_T_1959_en = T_1936;
  assign T_1909_T_1999_addr = {{1'd0}, 1'h0};
  assign T_1909_T_1999_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1909_T_1999_data = T_1909[T_1909_T_1999_addr];
  `else
  assign T_1909_T_1999_data = T_1909_T_1999_addr >= 2'h3 ? $random : T_1909[T_1909_T_1999_addr];
  `endif
  assign T_1909_T_2001_addr = {{1'd0}, 1'h1};
  assign T_1909_T_2001_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1909_T_2001_data = T_1909[T_1909_T_2001_addr];
  `else
  assign T_1909_T_2001_data = T_1909_T_2001_addr >= 2'h3 ? $random : T_1909[T_1909_T_2001_addr];
  `endif
  assign T_1909_T_2003_addr = 2'h2;
  assign T_1909_T_2003_en = 1'h1;
  `ifdef SYNTHESIS
  assign T_1909_T_2003_data = T_1909[T_1909_T_2003_addr];
  `else
  assign T_1909_T_2003_data = T_1909_T_2003_addr >= 2'h3 ? $random : T_1909[T_1909_T_2003_addr];
  `endif
  assign T_1909_T_1960_data = pte_ppn;
  assign T_1909_T_1960_addr = T_1957;
  assign T_1909_T_1960_mask = T_1936;
  assign T_1909_T_1960_en = T_1936;
  assign T_1912 = T_1906_T_1911_data == pte_addr;
  assign T_1915 = T_1906_T_1914_data == pte_addr;
  assign T_1918 = T_1906_T_1917_data == pte_addr;
  assign T_1924_0 = T_1912;
  assign T_1924_1 = T_1915;
  assign T_1924_2 = T_1918;
  assign T_1926 = {T_1924_2,T_1924_1};
  assign T_1927 = {T_1926,T_1924_0};
  assign T_1928 = T_1927 & T_1903;
  assign GEN_71 = {{2'd0}, 1'h0};
  assign pte_cache_hit = T_1928 != GEN_71;
  assign GEN_72 = {{2'd0}, 2'h2};
  assign T_1931 = pte_typ < GEN_72;
  assign T_1932 = pte_v & T_1931;
  assign T_1933 = io_mem_resp_valid & T_1932;
  assign T_1935 = pte_cache_hit == 1'h0;
  assign T_1936 = T_1933 & T_1935;
  assign T_1937 = ~ T_1903;
  assign T_1939 = T_1937 == GEN_71;
  assign T_1941 = T_1893 >> 1'h1;
  assign T_1942 = T_1941[0];
  assign T_1943 = {1'h1,T_1942};
  assign T_1944 = T_1893 >> T_1943;
  assign T_1945 = T_1944[0];
  assign T_1946 = {T_1943,T_1945};
  assign T_1947 = T_1946[1:0];
  assign T_1949 = T_1937[0];
  assign T_1950 = T_1937[1];
  assign T_1955 = T_1950 ? {{1'd0}, 1'h1} : 2'h2;
  assign T_1956 = T_1949 ? {{1'd0}, 1'h0} : T_1955;
  assign T_1957 = T_1939 ? T_1947 : T_1956;
  assign GEN_1 = 1'h1;
  assign GEN_74 = {{1'd0}, 1'h0};
  assign GEN_12 = GEN_74 == T_1957 ? GEN_1 : T_1900_0;
  assign GEN_13 = GEN_69 == T_1957 ? GEN_1 : T_1900_1;
  assign GEN_14 = 2'h2 == T_1957 ? GEN_1 : T_1900_2;
  assign GEN_16 = T_1936 ? GEN_12 : T_1900_0;
  assign GEN_17 = T_1936 ? GEN_13 : T_1900_1;
  assign GEN_18 = T_1936 ? GEN_14 : T_1900_2;
  assign T_1961 = state == 3'h1;
  assign T_1962 = pte_cache_hit & T_1961;
  assign T_1963 = T_1928[2];
  assign T_1964 = T_1928[1:0];
  assign GEN_76 = {{1'd0}, T_1963};
  assign T_1967 = GEN_76 | T_1964;
  assign T_1968 = T_1967[1];
  assign T_1969 = {T_1963,T_1968};
  assign T_1971 = T_1969[1];
  assign GEN_77 = {{1'd0}, 3'h1};
  assign T_1973 = GEN_77 << 1'h1;
  assign T_1974 = T_1973[2:0];
  assign T_1975 = ~ T_1974;
  assign T_1976 = T_1893 & T_1975;
  assign T_1978 = T_1971 ? {{2'd0}, 1'h0} : T_1974;
  assign T_1979 = T_1976 | T_1978;
  assign T_1980 = {1'h1,T_1971};
  assign T_1981 = T_1969[0];
  assign GEN_78 = {{3'd0}, 3'h1};
  assign T_1983 = GEN_78 << T_1980;
  assign T_1984 = T_1983[2:0];
  assign T_1985 = ~ T_1984;
  assign T_1986 = T_1979 & T_1985;
  assign T_1988 = T_1981 ? {{2'd0}, 1'h0} : T_1984;
  assign T_1989 = T_1986 | T_1988;
  assign GEN_29 = T_1962 ? T_1989 : T_1893;
  assign T_1991 = reset | io_dpath_invalidate;
  assign GEN_30 = T_1991 ? 1'h0 : GEN_16;
  assign GEN_31 = T_1991 ? 1'h0 : GEN_17;
  assign GEN_32 = T_1991 ? 1'h0 : GEN_18;
  assign T_1995 = T_1928[0];
  assign T_1996 = T_1928[1];
  assign T_2005 = T_1995 ? T_1909_T_1999_data : {{19'd0}, 1'h0};
  assign T_2007 = T_1996 ? T_1909_T_2001_data : {{19'd0}, 1'h0};
  assign T_2009 = T_1963 ? T_1909_T_2003_data : {{19'd0}, 1'h0};
  assign T_2011 = T_2005 | T_2007;
  assign T_2012 = T_2011 | T_2009;
  assign pte_cache_data = T_2012;
  assign T_2013 = r_req_prv[0];
  assign GEN_79 = {{1'd0}, 3'h4};
  assign T_2015 = pte_typ >= GEN_79;
  assign T_2016 = pte_v & T_2015;
  assign T_2017 = pte_typ[1];
  assign T_2018 = T_2016 & T_2017;
  assign T_2020 = pte_typ >= GEN_72;
  assign T_2021 = pte_v & T_2020;
  assign T_2022 = pte_typ[0];
  assign T_2023 = T_2021 & T_2022;
  assign T_2027 = r_req_store ? T_2023 : T_2021;
  assign T_2028 = r_req_fetch ? T_2018 : T_2027;
  assign T_2033 = pte_typ < 4'h8;
  assign T_2034 = T_2021 & T_2033;
  assign T_2036 = T_2034 & T_2017;
  assign T_2044 = T_2034 & T_2022;
  assign T_2051 = r_req_store ? T_2044 : T_2034;
  assign T_2052 = r_req_fetch ? T_2036 : T_2051;
  assign perm_ok = T_2013 ? T_2028 : T_2052;
  assign T_2054 = pte_r == 1'h0;
  assign T_2056 = pte_d == 1'h0;
  assign T_2057 = r_req_store & T_2056;
  assign T_2058 = T_2054 | T_2057;
  assign set_dirty_bit = perm_ok & T_2058;
  assign T_2059 = state == 3'h2;
  assign T_2060 = io_mem_resp_valid & T_2059;
  assign T_2062 = set_dirty_bit == 1'h0;
  assign T_2063 = T_2060 & T_2062;
  assign GEN_33 = T_2063 ? pte_ppn : GEN_11;
  assign GEN_34 = T_2063 ? pte_reserved_for_software : r_pte_reserved_for_software;
  assign GEN_35 = T_2063 ? pte_d : r_pte_d;
  assign GEN_36 = T_2063 ? pte_r : r_pte_r;
  assign GEN_37 = T_2063 ? pte_typ : r_pte_typ;
  assign GEN_38 = T_2063 ? pte_v : r_pte_v;
  assign T_2079_ppn = T_2093;
  assign T_2079_reserved_for_software = T_2092;
  assign T_2079_d = T_2091;
  assign T_2079_r = T_2090;
  assign T_2079_typ = T_2089;
  assign T_2079_v = T_2088;
  assign T_2087 = {{29'd0}, 1'h0};
  assign T_2088 = T_2087[0];
  assign T_2089 = T_2087[4:1];
  assign T_2090 = T_2087[5];
  assign T_2091 = T_2087[6];
  assign T_2092 = T_2087[9:7];
  assign T_2093 = T_2087[29:10];
  assign pte_wdata_ppn = T_2079_ppn;
  assign pte_wdata_reserved_for_software = T_2079_reserved_for_software;
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_r = 1'h1;
  assign pte_wdata_typ = T_2079_typ;
  assign pte_wdata_v = T_2079_v;
  assign T_2102 = state == 3'h3;
  assign T_2103 = T_1961 | T_2102;
  assign T_2106 = T_2102 ? 5'ha : 5'h0;
  assign T_2107 = {pte_wdata_r,pte_wdata_typ};
  assign T_2108 = {T_2107,pte_wdata_v};
  assign T_2109 = {pte_wdata_ppn,pte_wdata_reserved_for_software};
  assign T_2110 = {T_2109,pte_wdata_d};
  assign T_2111 = {T_2110,T_2108};
  assign r_resp_ppn = io_mem_req_bits_addr[39:12];
  assign T_2114 = r_resp_ppn[27:18];
  assign T_2115 = r_req_addr[17:0];
  assign T_2116 = {T_2114,T_2115};
  assign T_2117 = r_resp_ppn[27:9];
  assign T_2119 = {T_2117,T_1850};
  assign T_2125_0 = T_2116;
  assign T_2125_1 = T_2119;
  assign T_2125_2 = r_resp_ppn;
  assign resp_val = state == 3'h5;
  assign T_2128 = r_req_dest == 1'h0;
  assign T_2129 = resp_val & T_2128;
  assign GEN_2 = GEN_40;
  assign GEN_39 = GEN_69 == count ? T_2125_1 : T_2125_0;
  assign GEN_40 = 2'h2 == count ? T_2125_2 : GEN_39;
  assign T_2132 = resp_val & r_req_dest;
  assign GEN_3 = GEN_40;
  assign T_2133 = 3'h0 == state;
  assign GEN_43 = arb_io_out_valid ? 3'h1 : state;
  assign GEN_44 = T_2133 ? GEN_43 : state;
  assign GEN_45 = T_2133 ? {{1'd0}, 1'h0} : count;
  assign T_2135 = 3'h1 == state;
  assign T_2137 = count < 2'h2;
  assign T_2138 = pte_cache_hit & T_2137;
  assign T_2141 = count + GEN_69;
  assign T_2142 = T_2141[1:0];
  assign GEN_46 = T_2138 ? 1'h0 : T_2103;
  assign GEN_47 = T_2138 ? 3'h1 : GEN_44;
  assign GEN_48 = T_2138 ? T_2142 : GEN_45;
  assign GEN_49 = T_2138 ? pte_cache_data : GEN_33;
  assign T_2144 = T_2138 == 1'h0;
  assign T_2145 = T_2144 & io_mem_req_ready;
  assign GEN_50 = T_2145 ? 3'h2 : GEN_47;
  assign GEN_51 = T_2135 ? GEN_46 : T_2103;
  assign GEN_52 = T_2135 ? GEN_50 : GEN_44;
  assign GEN_53 = T_2135 ? GEN_48 : GEN_45;
  assign GEN_54 = T_2135 ? GEN_49 : GEN_33;
  assign T_2146 = 3'h2 == state;
  assign GEN_55 = io_mem_s2_nack ? 3'h1 : GEN_52;
  assign T_2150 = T_2021 & set_dirty_bit;
  assign GEN_56 = T_2150 ? 3'h3 : 3'h5;
  assign T_2156 = T_1932 & T_2137;
  assign GEN_57 = T_2156 ? 3'h1 : GEN_56;
  assign GEN_58 = T_2156 ? T_2142 : GEN_53;
  assign GEN_59 = io_mem_resp_valid ? GEN_57 : GEN_55;
  assign GEN_60 = io_mem_resp_valid ? GEN_58 : GEN_53;
  assign GEN_61 = T_2146 ? GEN_59 : GEN_52;
  assign GEN_62 = T_2146 ? GEN_60 : GEN_53;
  assign T_2160 = 3'h3 == state;
  assign GEN_63 = io_mem_req_ready ? 3'h4 : GEN_61;
  assign GEN_64 = T_2160 ? GEN_63 : GEN_61;
  assign T_2161 = 3'h4 == state;
  assign GEN_65 = io_mem_s2_nack ? 3'h3 : GEN_64;
  assign GEN_66 = io_mem_resp_valid ? 3'h1 : GEN_65;
  assign GEN_67 = T_2161 ? GEN_66 : GEN_64;
  assign T_2162 = 3'h5 == state;
  assign GEN_68 = T_2162 ? 3'h0 : GEN_67;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_20 = {1{$random}};
  state = GEN_20[2:0];
  GEN_21 = {1{$random}};
  count = GEN_21[1:0];
  GEN_22 = {1{$random}};
  r_req_addr = GEN_22[26:0];
  GEN_23 = {1{$random}};
  r_req_prv = GEN_23[1:0];
  GEN_24 = {1{$random}};
  r_req_store = GEN_24[0:0];
  GEN_25 = {1{$random}};
  r_req_fetch = GEN_25[0:0];
  GEN_26 = {1{$random}};
  r_req_dest = GEN_26[0:0];
  GEN_27 = {1{$random}};
  r_pte_ppn = GEN_27[19:0];
  GEN_28 = {1{$random}};
  r_pte_reserved_for_software = GEN_28[2:0];
  GEN_41 = {1{$random}};
  r_pte_d = GEN_41[0:0];
  GEN_42 = {1{$random}};
  r_pte_r = GEN_42[0:0];
  GEN_73 = {1{$random}};
  r_pte_typ = GEN_73[3:0];
  GEN_75 = {1{$random}};
  r_pte_v = GEN_75[0:0];
  GEN_80 = {1{$random}};
  T_1893 = GEN_80[2:0];
  GEN_81 = {1{$random}};
  T_1900_0 = GEN_81[0:0];
  GEN_82 = {1{$random}};
  T_1900_1 = GEN_82[0:0];
  GEN_83 = {1{$random}};
  T_1900_2 = GEN_83[0:0];
  GEN_84 = {1{$random}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    T_1906[initvar] = GEN_84[31:0];
  GEN_85 = {1{$random}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    T_1909[initvar] = GEN_85[19:0];
  GEN_86 = {1{$random}};
  GEN_15 = GEN_86[8:0];
  GEN_87 = {2{$random}};
  GEN_19 = GEN_87[63:0];
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      state <= 3'h0;
    end else begin
      state <= GEN_68;
    end
    if(1'h0) begin
    end else begin
      count <= GEN_62;
    end
    if(1'h0) begin
    end else begin
      r_req_addr <= GEN_6;
    end
    if(1'h0) begin
    end else begin
      r_req_prv <= GEN_7;
    end
    if(1'h0) begin
    end else begin
      r_req_store <= GEN_8;
    end
    if(1'h0) begin
    end else begin
      r_req_fetch <= GEN_9;
    end
    if(1'h0) begin
    end else begin
      r_req_dest <= GEN_10;
    end
    if(1'h0) begin
    end else begin
      r_pte_ppn <= GEN_54;
    end
    if(1'h0) begin
    end else begin
      r_pte_reserved_for_software <= GEN_34;
    end
    if(1'h0) begin
    end else begin
      r_pte_d <= GEN_35;
    end
    if(1'h0) begin
    end else begin
      r_pte_r <= GEN_36;
    end
    if(1'h0) begin
    end else begin
      r_pte_typ <= GEN_37;
    end
    if(1'h0) begin
    end else begin
      r_pte_v <= GEN_38;
    end
    if(1'h0) begin
    end else begin
      T_1893 <= GEN_29;
    end
    if(1'h0) begin
    end else begin
      T_1900_0 <= GEN_30;
    end
    if(1'h0) begin
    end else begin
      T_1900_1 <= GEN_31;
    end
    if(1'h0) begin
    end else begin
      T_1900_2 <= GEN_32;
    end
    if(T_1906_T_1959_en & T_1906_T_1959_mask) begin
      T_1906[T_1906_T_1959_addr] <= T_1906_T_1959_data;
    end
    if(T_1909_T_1960_en & T_1909_T_1960_mask) begin
      T_1909[T_1909_T_1960_addr] <= T_1909_T_1960_data;
    end
  end
endmodule
module HellaCacheArbiter(
  input   clk,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [39:0] io_requestor_0_req_bits_addr,
  input  [8:0] io_requestor_0_req_bits_tag,
  input  [4:0] io_requestor_0_req_bits_cmd,
  input  [2:0] io_requestor_0_req_bits_typ,
  input   io_requestor_0_req_bits_phys,
  input  [63:0] io_requestor_0_req_bits_data,
  input   io_requestor_0_s1_kill,
  input  [63:0] io_requestor_0_s1_data,
  output  io_requestor_0_s2_nack,
  output  io_requestor_0_resp_valid,
  output [39:0] io_requestor_0_resp_bits_addr,
  output [8:0] io_requestor_0_resp_bits_tag,
  output [4:0] io_requestor_0_resp_bits_cmd,
  output [2:0] io_requestor_0_resp_bits_typ,
  output [63:0] io_requestor_0_resp_bits_data,
  output  io_requestor_0_resp_bits_replay,
  output  io_requestor_0_resp_bits_has_data,
  output [63:0] io_requestor_0_resp_bits_data_word_bypass,
  output [63:0] io_requestor_0_resp_bits_store_data,
  output  io_requestor_0_replay_next,
  output  io_requestor_0_xcpt_ma_ld,
  output  io_requestor_0_xcpt_ma_st,
  output  io_requestor_0_xcpt_pf_ld,
  output  io_requestor_0_xcpt_pf_st,
  input   io_requestor_0_invalidate_lr,
  output  io_requestor_0_ordered,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [39:0] io_requestor_1_req_bits_addr,
  input  [8:0] io_requestor_1_req_bits_tag,
  input  [4:0] io_requestor_1_req_bits_cmd,
  input  [2:0] io_requestor_1_req_bits_typ,
  input   io_requestor_1_req_bits_phys,
  input  [63:0] io_requestor_1_req_bits_data,
  input   io_requestor_1_s1_kill,
  input  [63:0] io_requestor_1_s1_data,
  output  io_requestor_1_s2_nack,
  output  io_requestor_1_resp_valid,
  output [39:0] io_requestor_1_resp_bits_addr,
  output [8:0] io_requestor_1_resp_bits_tag,
  output [4:0] io_requestor_1_resp_bits_cmd,
  output [2:0] io_requestor_1_resp_bits_typ,
  output [63:0] io_requestor_1_resp_bits_data,
  output  io_requestor_1_resp_bits_replay,
  output  io_requestor_1_resp_bits_has_data,
  output [63:0] io_requestor_1_resp_bits_data_word_bypass,
  output [63:0] io_requestor_1_resp_bits_store_data,
  output  io_requestor_1_replay_next,
  output  io_requestor_1_xcpt_ma_ld,
  output  io_requestor_1_xcpt_ma_st,
  output  io_requestor_1_xcpt_pf_ld,
  output  io_requestor_1_xcpt_pf_st,
  input   io_requestor_1_invalidate_lr,
  output  io_requestor_1_ordered,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [8:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,
  input  [39:0] io_mem_resp_bits_addr,
  input  [8:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,
  input  [63:0] io_mem_resp_bits_data,
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered
);
  reg  s1_id;
  reg [31:0] GEN_9;
  reg  s2_id;
  reg [31:0] GEN_10;
  wire  T_7160;
  wire  T_7161;
  wire  T_7163;
  wire  T_7164;
  wire [9:0] T_7166;
  wire [9:0] T_7169;
  wire [4:0] GEN_0;
  wire [2:0] GEN_1;
  wire [39:0] GEN_2;
  wire  GEN_3;
  wire [9:0] GEN_4;
  wire  GEN_5;
  wire  T_7172;
  wire  GEN_6;
  wire [63:0] GEN_7;
  wire  T_7173;
  wire  T_7175;
  wire  T_7176;
  wire  T_7178;
  wire  T_7179;
  wire [7:0] T_7180;
  wire  T_7184;
  wire  T_7187;
  reg [63:0] GEN_8;
  reg [63:0] GEN_11;
  assign io_requestor_0_req_ready = io_mem_req_ready;
  assign io_requestor_0_s2_nack = T_7179;
  assign io_requestor_0_resp_valid = T_7176;
  assign io_requestor_0_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_0_resp_bits_tag = {{1'd0}, T_7180};
  assign io_requestor_0_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_0_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_0_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_0_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_0_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_0_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_0_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_0_replay_next = io_mem_replay_next;
  assign io_requestor_0_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_0_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_0_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_0_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_0_ordered = io_mem_ordered;
  assign io_requestor_1_req_ready = T_7164;
  assign io_requestor_1_s2_nack = T_7187;
  assign io_requestor_1_resp_valid = T_7184;
  assign io_requestor_1_resp_bits_addr = io_mem_resp_bits_addr;
  assign io_requestor_1_resp_bits_tag = {{1'd0}, T_7180};
  assign io_requestor_1_resp_bits_cmd = io_mem_resp_bits_cmd;
  assign io_requestor_1_resp_bits_typ = io_mem_resp_bits_typ;
  assign io_requestor_1_resp_bits_data = io_mem_resp_bits_data;
  assign io_requestor_1_resp_bits_replay = io_mem_resp_bits_replay;
  assign io_requestor_1_resp_bits_has_data = io_mem_resp_bits_has_data;
  assign io_requestor_1_resp_bits_data_word_bypass = io_mem_resp_bits_data_word_bypass;
  assign io_requestor_1_resp_bits_store_data = io_mem_resp_bits_store_data;
  assign io_requestor_1_replay_next = io_mem_replay_next;
  assign io_requestor_1_xcpt_ma_ld = io_mem_xcpt_ma_ld;
  assign io_requestor_1_xcpt_ma_st = io_mem_xcpt_ma_st;
  assign io_requestor_1_xcpt_pf_ld = io_mem_xcpt_pf_ld;
  assign io_requestor_1_xcpt_pf_st = io_mem_xcpt_pf_st;
  assign io_requestor_1_ordered = io_mem_ordered;
  assign io_mem_req_valid = T_7161;
  assign io_mem_req_bits_addr = GEN_2;
  assign io_mem_req_bits_tag = GEN_4[8:0];
  assign io_mem_req_bits_cmd = GEN_0;
  assign io_mem_req_bits_typ = GEN_1;
  assign io_mem_req_bits_phys = GEN_3;
  assign io_mem_req_bits_data = GEN_8;
  assign io_mem_s1_kill = GEN_6;
  assign io_mem_s1_data = GEN_7;
  assign io_mem_invalidate_lr = T_7160;
  assign T_7160 = io_requestor_0_invalidate_lr | io_requestor_1_invalidate_lr;
  assign T_7161 = io_requestor_0_req_valid | io_requestor_1_req_valid;
  assign T_7163 = io_requestor_0_req_valid == 1'h0;
  assign T_7164 = io_requestor_0_req_ready & T_7163;
  assign T_7166 = {io_requestor_1_req_bits_tag,1'h1};
  assign T_7169 = {io_requestor_0_req_bits_tag,1'h0};
  assign GEN_0 = io_requestor_0_req_valid ? io_requestor_0_req_bits_cmd : io_requestor_1_req_bits_cmd;
  assign GEN_1 = io_requestor_0_req_valid ? io_requestor_0_req_bits_typ : io_requestor_1_req_bits_typ;
  assign GEN_2 = io_requestor_0_req_valid ? io_requestor_0_req_bits_addr : io_requestor_1_req_bits_addr;
  assign GEN_3 = io_requestor_0_req_valid ? io_requestor_0_req_bits_phys : io_requestor_1_req_bits_phys;
  assign GEN_4 = io_requestor_0_req_valid ? T_7169 : T_7166;
  assign GEN_5 = io_requestor_0_req_valid ? 1'h0 : 1'h1;
  assign T_7172 = s1_id == 1'h0;
  assign GEN_6 = T_7172 ? io_requestor_0_s1_kill : io_requestor_1_s1_kill;
  assign GEN_7 = T_7172 ? io_requestor_0_s1_data : io_requestor_1_s1_data;
  assign T_7173 = io_mem_resp_bits_tag[0];
  assign T_7175 = T_7173 == 1'h0;
  assign T_7176 = io_mem_resp_valid & T_7175;
  assign T_7178 = s2_id == 1'h0;
  assign T_7179 = io_mem_s2_nack & T_7178;
  assign T_7180 = io_mem_resp_bits_tag[8:1];
  assign T_7184 = io_mem_resp_valid & T_7173;
  assign T_7187 = io_mem_s2_nack & s2_id;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_9 = {1{$random}};
  s1_id = GEN_9[0:0];
  GEN_10 = {1{$random}};
  s2_id = GEN_10[0:0];
  GEN_11 = {2{$random}};
  GEN_8 = GEN_11[63:0];
  end
`endif
  always @(posedge clk) begin
    if(1'h0) begin
    end else begin
      s1_id <= GEN_5;
    end
    if(1'h0) begin
    end else begin
      s2_id <= s1_id;
    end
  end
endmodule
module RocketTile(
  input   clk,
  input   reset,
  input   io_cached_0_acquire_ready,
  output  io_cached_0_acquire_valid,
  output [25:0] io_cached_0_acquire_bits_addr_block,
  output [1:0] io_cached_0_acquire_bits_client_xact_id,
  output [2:0] io_cached_0_acquire_bits_addr_beat,
  output  io_cached_0_acquire_bits_is_builtin_type,
  output [2:0] io_cached_0_acquire_bits_a_type,
  output [11:0] io_cached_0_acquire_bits_union,
  output [63:0] io_cached_0_acquire_bits_data,
  output  io_cached_0_probe_ready,
  input   io_cached_0_probe_valid,
  input  [25:0] io_cached_0_probe_bits_addr_block,
  input  [1:0] io_cached_0_probe_bits_p_type,
  input   io_cached_0_release_ready,
  output  io_cached_0_release_valid,
  output [2:0] io_cached_0_release_bits_addr_beat,
  output [25:0] io_cached_0_release_bits_addr_block,
  output [1:0] io_cached_0_release_bits_client_xact_id,
  output  io_cached_0_release_bits_voluntary,
  output [2:0] io_cached_0_release_bits_r_type,
  output [63:0] io_cached_0_release_bits_data,
  output  io_cached_0_grant_ready,
  input   io_cached_0_grant_valid,
  input  [2:0] io_cached_0_grant_bits_addr_beat,
  input  [1:0] io_cached_0_grant_bits_client_xact_id,
  input  [2:0] io_cached_0_grant_bits_manager_xact_id,
  input   io_cached_0_grant_bits_is_builtin_type,
  input  [3:0] io_cached_0_grant_bits_g_type,
  input  [63:0] io_cached_0_grant_bits_data,
  input   io_cached_0_grant_bits_manager_id,
  input   io_cached_0_finish_ready,
  output  io_cached_0_finish_valid,
  output [2:0] io_cached_0_finish_bits_manager_xact_id,
  output  io_cached_0_finish_bits_manager_id,
  input   io_uncached_0_acquire_ready,
  output  io_uncached_0_acquire_valid,
  output [25:0] io_uncached_0_acquire_bits_addr_block,
  output [1:0] io_uncached_0_acquire_bits_client_xact_id,
  output [2:0] io_uncached_0_acquire_bits_addr_beat,
  output  io_uncached_0_acquire_bits_is_builtin_type,
  output [2:0] io_uncached_0_acquire_bits_a_type,
  output [11:0] io_uncached_0_acquire_bits_union,
  output [63:0] io_uncached_0_acquire_bits_data,
  output  io_uncached_0_grant_ready,
  input   io_uncached_0_grant_valid,
  input  [2:0] io_uncached_0_grant_bits_addr_beat,
  input  [1:0] io_uncached_0_grant_bits_client_xact_id,
  input  [2:0] io_uncached_0_grant_bits_manager_xact_id,
  input   io_uncached_0_grant_bits_is_builtin_type,
  input  [3:0] io_uncached_0_grant_bits_g_type,
  input  [63:0] io_uncached_0_grant_bits_data,
  input   io_prci_reset,
  input   io_prci_id,
  input   io_prci_interrupts_mtip,
  input   io_prci_interrupts_meip,
  input   io_prci_interrupts_seip,
  input   io_prci_interrupts_debug,
  input   io_prci_interrupts_msip,
  input   io_dma_req_ready,
  output  io_dma_req_valid,
  output [1:0] io_dma_req_bits_xact_id,
  output  io_dma_req_bits_client_id,
  output [2:0] io_dma_req_bits_cmd,
  output [31:0] io_dma_req_bits_source,
  output [31:0] io_dma_req_bits_dest,
  output [31:0] io_dma_req_bits_length,
  output [1:0] io_dma_req_bits_size,
  output  io_dma_resp_ready,
  input   io_dma_resp_valid,
  input  [1:0] io_dma_resp_bits_xact_id,
  input   io_dma_resp_bits_client_id,
  input  [1:0] io_dma_resp_bits_status
);
  wire  core_clk;
  wire  core_reset;
  wire  core_io_prci_reset;
  wire  core_io_prci_id;
  wire  core_io_prci_interrupts_mtip;
  wire  core_io_prci_interrupts_meip;
  wire  core_io_prci_interrupts_seip;
  wire  core_io_prci_interrupts_debug;
  wire  core_io_prci_interrupts_msip;
  wire  core_io_imem_req_valid;
  wire [39:0] core_io_imem_req_bits_pc;
  wire  core_io_imem_resp_ready;
  wire  core_io_imem_resp_valid;
  wire [39:0] core_io_imem_resp_bits_pc;
  wire [31:0] core_io_imem_resp_bits_data_0;
  wire  core_io_imem_resp_bits_mask;
  wire  core_io_imem_resp_bits_xcpt_if;
  wire  core_io_imem_btb_resp_valid;
  wire  core_io_imem_btb_resp_bits_taken;
  wire  core_io_imem_btb_resp_bits_mask;
  wire  core_io_imem_btb_resp_bits_bridx;
  wire [38:0] core_io_imem_btb_resp_bits_target;
  wire [5:0] core_io_imem_btb_resp_bits_entry;
  wire [6:0] core_io_imem_btb_resp_bits_bht_history;
  wire [1:0] core_io_imem_btb_resp_bits_bht_value;
  wire  core_io_imem_btb_update_valid;
  wire  core_io_imem_btb_update_bits_prediction_valid;
  wire  core_io_imem_btb_update_bits_prediction_bits_taken;
  wire  core_io_imem_btb_update_bits_prediction_bits_mask;
  wire  core_io_imem_btb_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_btb_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_btb_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_btb_update_bits_pc;
  wire [38:0] core_io_imem_btb_update_bits_target;
  wire  core_io_imem_btb_update_bits_taken;
  wire  core_io_imem_btb_update_bits_isJump;
  wire  core_io_imem_btb_update_bits_isReturn;
  wire [38:0] core_io_imem_btb_update_bits_br_pc;
  wire  core_io_imem_bht_update_valid;
  wire  core_io_imem_bht_update_bits_prediction_valid;
  wire  core_io_imem_bht_update_bits_prediction_bits_taken;
  wire  core_io_imem_bht_update_bits_prediction_bits_mask;
  wire  core_io_imem_bht_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_bht_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_bht_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] core_io_imem_bht_update_bits_pc;
  wire  core_io_imem_bht_update_bits_taken;
  wire  core_io_imem_bht_update_bits_mispredict;
  wire  core_io_imem_ras_update_valid;
  wire  core_io_imem_ras_update_bits_isCall;
  wire  core_io_imem_ras_update_bits_isReturn;
  wire [38:0] core_io_imem_ras_update_bits_returnAddr;
  wire  core_io_imem_ras_update_bits_prediction_valid;
  wire  core_io_imem_ras_update_bits_prediction_bits_taken;
  wire  core_io_imem_ras_update_bits_prediction_bits_mask;
  wire  core_io_imem_ras_update_bits_prediction_bits_bridx;
  wire [38:0] core_io_imem_ras_update_bits_prediction_bits_target;
  wire [5:0] core_io_imem_ras_update_bits_prediction_bits_entry;
  wire [6:0] core_io_imem_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] core_io_imem_ras_update_bits_prediction_bits_bht_value;
  wire  core_io_imem_flush_icache;
  wire  core_io_imem_flush_tlb;
  wire [39:0] core_io_imem_npc;
  wire  core_io_dmem_req_ready;
  wire  core_io_dmem_req_valid;
  wire [39:0] core_io_dmem_req_bits_addr;
  wire [8:0] core_io_dmem_req_bits_tag;
  wire [4:0] core_io_dmem_req_bits_cmd;
  wire [2:0] core_io_dmem_req_bits_typ;
  wire  core_io_dmem_req_bits_phys;
  wire [63:0] core_io_dmem_req_bits_data;
  wire  core_io_dmem_s1_kill;
  wire [63:0] core_io_dmem_s1_data;
  wire  core_io_dmem_s2_nack;
  wire  core_io_dmem_resp_valid;
  wire [39:0] core_io_dmem_resp_bits_addr;
  wire [8:0] core_io_dmem_resp_bits_tag;
  wire [4:0] core_io_dmem_resp_bits_cmd;
  wire [2:0] core_io_dmem_resp_bits_typ;
  wire [63:0] core_io_dmem_resp_bits_data;
  wire  core_io_dmem_resp_bits_replay;
  wire  core_io_dmem_resp_bits_has_data;
  wire [63:0] core_io_dmem_resp_bits_data_word_bypass;
  wire [63:0] core_io_dmem_resp_bits_store_data;
  wire  core_io_dmem_replay_next;
  wire  core_io_dmem_xcpt_ma_ld;
  wire  core_io_dmem_xcpt_ma_st;
  wire  core_io_dmem_xcpt_pf_ld;
  wire  core_io_dmem_xcpt_pf_st;
  wire  core_io_dmem_invalidate_lr;
  wire  core_io_dmem_ordered;
  wire [19:0] core_io_ptw_ptbr;
  wire  core_io_ptw_invalidate;
  wire  core_io_ptw_status_debug;
  wire [1:0] core_io_ptw_status_prv;
  wire  core_io_ptw_status_sd;
  wire [30:0] core_io_ptw_status_zero3;
  wire  core_io_ptw_status_sd_rv32;
  wire [1:0] core_io_ptw_status_zero2;
  wire [4:0] core_io_ptw_status_vm;
  wire [4:0] core_io_ptw_status_zero1;
  wire  core_io_ptw_status_pum;
  wire  core_io_ptw_status_mprv;
  wire [1:0] core_io_ptw_status_xs;
  wire [1:0] core_io_ptw_status_fs;
  wire [1:0] core_io_ptw_status_mpp;
  wire [1:0] core_io_ptw_status_hpp;
  wire  core_io_ptw_status_spp;
  wire  core_io_ptw_status_mpie;
  wire  core_io_ptw_status_hpie;
  wire  core_io_ptw_status_spie;
  wire  core_io_ptw_status_upie;
  wire  core_io_ptw_status_mie;
  wire  core_io_ptw_status_hie;
  wire  core_io_ptw_status_sie;
  wire  core_io_ptw_status_uie;
  wire [31:0] core_io_fpu_inst;
  wire [63:0] core_io_fpu_fromint_data;
  wire [2:0] core_io_fpu_fcsr_rm;
  wire  core_io_fpu_fcsr_flags_valid;
  wire [4:0] core_io_fpu_fcsr_flags_bits;
  wire [63:0] core_io_fpu_store_data;
  wire [63:0] core_io_fpu_toint_data;
  wire  core_io_fpu_dmem_resp_val;
  wire [2:0] core_io_fpu_dmem_resp_type;
  wire [4:0] core_io_fpu_dmem_resp_tag;
  wire [63:0] core_io_fpu_dmem_resp_data;
  wire  core_io_fpu_valid;
  wire  core_io_fpu_fcsr_rdy;
  wire  core_io_fpu_nack_mem;
  wire  core_io_fpu_illegal_rm;
  wire  core_io_fpu_killx;
  wire  core_io_fpu_killm;
  wire [4:0] core_io_fpu_dec_cmd;
  wire  core_io_fpu_dec_ldst;
  wire  core_io_fpu_dec_wen;
  wire  core_io_fpu_dec_ren1;
  wire  core_io_fpu_dec_ren2;
  wire  core_io_fpu_dec_ren3;
  wire  core_io_fpu_dec_swap12;
  wire  core_io_fpu_dec_swap23;
  wire  core_io_fpu_dec_single;
  wire  core_io_fpu_dec_fromint;
  wire  core_io_fpu_dec_toint;
  wire  core_io_fpu_dec_fastpipe;
  wire  core_io_fpu_dec_fma;
  wire  core_io_fpu_dec_div;
  wire  core_io_fpu_dec_sqrt;
  wire  core_io_fpu_dec_round;
  wire  core_io_fpu_dec_wflags;
  wire  core_io_fpu_sboard_set;
  wire  core_io_fpu_sboard_clr;
  wire [4:0] core_io_fpu_sboard_clra;
  wire  core_io_fpu_cp_req_ready;
  wire  core_io_fpu_cp_req_valid;
  wire [4:0] core_io_fpu_cp_req_bits_cmd;
  wire  core_io_fpu_cp_req_bits_ldst;
  wire  core_io_fpu_cp_req_bits_wen;
  wire  core_io_fpu_cp_req_bits_ren1;
  wire  core_io_fpu_cp_req_bits_ren2;
  wire  core_io_fpu_cp_req_bits_ren3;
  wire  core_io_fpu_cp_req_bits_swap12;
  wire  core_io_fpu_cp_req_bits_swap23;
  wire  core_io_fpu_cp_req_bits_single;
  wire  core_io_fpu_cp_req_bits_fromint;
  wire  core_io_fpu_cp_req_bits_toint;
  wire  core_io_fpu_cp_req_bits_fastpipe;
  wire  core_io_fpu_cp_req_bits_fma;
  wire  core_io_fpu_cp_req_bits_div;
  wire  core_io_fpu_cp_req_bits_sqrt;
  wire  core_io_fpu_cp_req_bits_round;
  wire  core_io_fpu_cp_req_bits_wflags;
  wire [2:0] core_io_fpu_cp_req_bits_rm;
  wire [1:0] core_io_fpu_cp_req_bits_typ;
  wire [64:0] core_io_fpu_cp_req_bits_in1;
  wire [64:0] core_io_fpu_cp_req_bits_in2;
  wire [64:0] core_io_fpu_cp_req_bits_in3;
  wire  core_io_fpu_cp_resp_ready;
  wire  core_io_fpu_cp_resp_valid;
  wire [64:0] core_io_fpu_cp_resp_bits_data;
  wire [4:0] core_io_fpu_cp_resp_bits_exc;
  wire  core_io_rocc_cmd_ready;
  wire  core_io_rocc_cmd_valid;
  wire [6:0] core_io_rocc_cmd_bits_inst_funct;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rs1;
  wire  core_io_rocc_cmd_bits_inst_xd;
  wire  core_io_rocc_cmd_bits_inst_xs1;
  wire  core_io_rocc_cmd_bits_inst_xs2;
  wire [4:0] core_io_rocc_cmd_bits_inst_rd;
  wire [6:0] core_io_rocc_cmd_bits_inst_opcode;
  wire [63:0] core_io_rocc_cmd_bits_rs1;
  wire [63:0] core_io_rocc_cmd_bits_rs2;
  wire  core_io_rocc_resp_ready;
  wire  core_io_rocc_resp_valid;
  wire [4:0] core_io_rocc_resp_bits_rd;
  wire [63:0] core_io_rocc_resp_bits_data;
  wire  core_io_rocc_mem_req_ready;
  wire  core_io_rocc_mem_req_valid;
  wire [39:0] core_io_rocc_mem_req_bits_addr;
  wire [8:0] core_io_rocc_mem_req_bits_tag;
  wire [4:0] core_io_rocc_mem_req_bits_cmd;
  wire [2:0] core_io_rocc_mem_req_bits_typ;
  wire  core_io_rocc_mem_req_bits_phys;
  wire [63:0] core_io_rocc_mem_req_bits_data;
  wire  core_io_rocc_mem_s1_kill;
  wire [63:0] core_io_rocc_mem_s1_data;
  wire  core_io_rocc_mem_s2_nack;
  wire  core_io_rocc_mem_resp_valid;
  wire [39:0] core_io_rocc_mem_resp_bits_addr;
  wire [8:0] core_io_rocc_mem_resp_bits_tag;
  wire [4:0] core_io_rocc_mem_resp_bits_cmd;
  wire [2:0] core_io_rocc_mem_resp_bits_typ;
  wire [63:0] core_io_rocc_mem_resp_bits_data;
  wire  core_io_rocc_mem_resp_bits_replay;
  wire  core_io_rocc_mem_resp_bits_has_data;
  wire [63:0] core_io_rocc_mem_resp_bits_data_word_bypass;
  wire [63:0] core_io_rocc_mem_resp_bits_store_data;
  wire  core_io_rocc_mem_replay_next;
  wire  core_io_rocc_mem_xcpt_ma_ld;
  wire  core_io_rocc_mem_xcpt_ma_st;
  wire  core_io_rocc_mem_xcpt_pf_ld;
  wire  core_io_rocc_mem_xcpt_pf_st;
  wire  core_io_rocc_mem_invalidate_lr;
  wire  core_io_rocc_mem_ordered;
  wire  core_io_rocc_busy;
  wire  core_io_rocc_status_debug;
  wire [1:0] core_io_rocc_status_prv;
  wire  core_io_rocc_status_sd;
  wire [30:0] core_io_rocc_status_zero3;
  wire  core_io_rocc_status_sd_rv32;
  wire [1:0] core_io_rocc_status_zero2;
  wire [4:0] core_io_rocc_status_vm;
  wire [4:0] core_io_rocc_status_zero1;
  wire  core_io_rocc_status_pum;
  wire  core_io_rocc_status_mprv;
  wire [1:0] core_io_rocc_status_xs;
  wire [1:0] core_io_rocc_status_fs;
  wire [1:0] core_io_rocc_status_mpp;
  wire [1:0] core_io_rocc_status_hpp;
  wire  core_io_rocc_status_spp;
  wire  core_io_rocc_status_mpie;
  wire  core_io_rocc_status_hpie;
  wire  core_io_rocc_status_spie;
  wire  core_io_rocc_status_upie;
  wire  core_io_rocc_status_mie;
  wire  core_io_rocc_status_hie;
  wire  core_io_rocc_status_sie;
  wire  core_io_rocc_status_uie;
  wire  core_io_rocc_interrupt;
  wire  core_io_rocc_autl_acquire_ready;
  wire  core_io_rocc_autl_acquire_valid;
  wire [25:0] core_io_rocc_autl_acquire_bits_addr_block;
  wire [1:0] core_io_rocc_autl_acquire_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_acquire_bits_addr_beat;
  wire  core_io_rocc_autl_acquire_bits_is_builtin_type;
  wire [2:0] core_io_rocc_autl_acquire_bits_a_type;
  wire [11:0] core_io_rocc_autl_acquire_bits_union;
  wire [63:0] core_io_rocc_autl_acquire_bits_data;
  wire  core_io_rocc_autl_grant_ready;
  wire  core_io_rocc_autl_grant_valid;
  wire [2:0] core_io_rocc_autl_grant_bits_addr_beat;
  wire [1:0] core_io_rocc_autl_grant_bits_client_xact_id;
  wire [2:0] core_io_rocc_autl_grant_bits_manager_xact_id;
  wire  core_io_rocc_autl_grant_bits_is_builtin_type;
  wire [3:0] core_io_rocc_autl_grant_bits_g_type;
  wire [63:0] core_io_rocc_autl_grant_bits_data;
  wire  core_io_rocc_fpu_req_ready;
  wire  core_io_rocc_fpu_req_valid;
  wire [4:0] core_io_rocc_fpu_req_bits_cmd;
  wire  core_io_rocc_fpu_req_bits_ldst;
  wire  core_io_rocc_fpu_req_bits_wen;
  wire  core_io_rocc_fpu_req_bits_ren1;
  wire  core_io_rocc_fpu_req_bits_ren2;
  wire  core_io_rocc_fpu_req_bits_ren3;
  wire  core_io_rocc_fpu_req_bits_swap12;
  wire  core_io_rocc_fpu_req_bits_swap23;
  wire  core_io_rocc_fpu_req_bits_single;
  wire  core_io_rocc_fpu_req_bits_fromint;
  wire  core_io_rocc_fpu_req_bits_toint;
  wire  core_io_rocc_fpu_req_bits_fastpipe;
  wire  core_io_rocc_fpu_req_bits_fma;
  wire  core_io_rocc_fpu_req_bits_div;
  wire  core_io_rocc_fpu_req_bits_sqrt;
  wire  core_io_rocc_fpu_req_bits_round;
  wire  core_io_rocc_fpu_req_bits_wflags;
  wire [2:0] core_io_rocc_fpu_req_bits_rm;
  wire [1:0] core_io_rocc_fpu_req_bits_typ;
  wire [64:0] core_io_rocc_fpu_req_bits_in1;
  wire [64:0] core_io_rocc_fpu_req_bits_in2;
  wire [64:0] core_io_rocc_fpu_req_bits_in3;
  wire  core_io_rocc_fpu_resp_ready;
  wire  core_io_rocc_fpu_resp_valid;
  wire [64:0] core_io_rocc_fpu_resp_bits_data;
  wire [4:0] core_io_rocc_fpu_resp_bits_exc;
  wire  core_io_rocc_exception;
  wire [11:0] core_io_rocc_csr_waddr;
  wire [63:0] core_io_rocc_csr_wdata;
  wire  core_io_rocc_csr_wen;
  wire  core_io_rocc_host_id;
  wire  icache_clk;
  wire  icache_reset;
  wire  icache_io_cpu_req_valid;
  wire [39:0] icache_io_cpu_req_bits_pc;
  wire  icache_io_cpu_resp_ready;
  wire  icache_io_cpu_resp_valid;
  wire [39:0] icache_io_cpu_resp_bits_pc;
  wire [31:0] icache_io_cpu_resp_bits_data_0;
  wire  icache_io_cpu_resp_bits_mask;
  wire  icache_io_cpu_resp_bits_xcpt_if;
  wire  icache_io_cpu_btb_resp_valid;
  wire  icache_io_cpu_btb_resp_bits_taken;
  wire  icache_io_cpu_btb_resp_bits_mask;
  wire  icache_io_cpu_btb_resp_bits_bridx;
  wire [38:0] icache_io_cpu_btb_resp_bits_target;
  wire [5:0] icache_io_cpu_btb_resp_bits_entry;
  wire [6:0] icache_io_cpu_btb_resp_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_resp_bits_bht_value;
  wire  icache_io_cpu_btb_update_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_valid;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_btb_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_btb_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_btb_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_btb_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_btb_update_bits_pc;
  wire [38:0] icache_io_cpu_btb_update_bits_target;
  wire  icache_io_cpu_btb_update_bits_taken;
  wire  icache_io_cpu_btb_update_bits_isJump;
  wire  icache_io_cpu_btb_update_bits_isReturn;
  wire [38:0] icache_io_cpu_btb_update_bits_br_pc;
  wire  icache_io_cpu_bht_update_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_valid;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_bht_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_bht_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_bht_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_bht_update_bits_prediction_bits_bht_value;
  wire [38:0] icache_io_cpu_bht_update_bits_pc;
  wire  icache_io_cpu_bht_update_bits_taken;
  wire  icache_io_cpu_bht_update_bits_mispredict;
  wire  icache_io_cpu_ras_update_valid;
  wire  icache_io_cpu_ras_update_bits_isCall;
  wire  icache_io_cpu_ras_update_bits_isReturn;
  wire [38:0] icache_io_cpu_ras_update_bits_returnAddr;
  wire  icache_io_cpu_ras_update_bits_prediction_valid;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_taken;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_mask;
  wire  icache_io_cpu_ras_update_bits_prediction_bits_bridx;
  wire [38:0] icache_io_cpu_ras_update_bits_prediction_bits_target;
  wire [5:0] icache_io_cpu_ras_update_bits_prediction_bits_entry;
  wire [6:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_history;
  wire [1:0] icache_io_cpu_ras_update_bits_prediction_bits_bht_value;
  wire  icache_io_cpu_flush_icache;
  wire  icache_io_cpu_flush_tlb;
  wire [39:0] icache_io_cpu_npc;
  wire  icache_io_ptw_req_ready;
  wire  icache_io_ptw_req_valid;
  wire [26:0] icache_io_ptw_req_bits_addr;
  wire [1:0] icache_io_ptw_req_bits_prv;
  wire  icache_io_ptw_req_bits_store;
  wire  icache_io_ptw_req_bits_fetch;
  wire  icache_io_ptw_resp_valid;
  wire [19:0] icache_io_ptw_resp_bits_pte_ppn;
  wire [2:0] icache_io_ptw_resp_bits_pte_reserved_for_software;
  wire  icache_io_ptw_resp_bits_pte_d;
  wire  icache_io_ptw_resp_bits_pte_r;
  wire [3:0] icache_io_ptw_resp_bits_pte_typ;
  wire  icache_io_ptw_resp_bits_pte_v;
  wire  icache_io_ptw_status_debug;
  wire [1:0] icache_io_ptw_status_prv;
  wire  icache_io_ptw_status_sd;
  wire [30:0] icache_io_ptw_status_zero3;
  wire  icache_io_ptw_status_sd_rv32;
  wire [1:0] icache_io_ptw_status_zero2;
  wire [4:0] icache_io_ptw_status_vm;
  wire [4:0] icache_io_ptw_status_zero1;
  wire  icache_io_ptw_status_pum;
  wire  icache_io_ptw_status_mprv;
  wire [1:0] icache_io_ptw_status_xs;
  wire [1:0] icache_io_ptw_status_fs;
  wire [1:0] icache_io_ptw_status_mpp;
  wire [1:0] icache_io_ptw_status_hpp;
  wire  icache_io_ptw_status_spp;
  wire  icache_io_ptw_status_mpie;
  wire  icache_io_ptw_status_hpie;
  wire  icache_io_ptw_status_spie;
  wire  icache_io_ptw_status_upie;
  wire  icache_io_ptw_status_mie;
  wire  icache_io_ptw_status_hie;
  wire  icache_io_ptw_status_sie;
  wire  icache_io_ptw_status_uie;
  wire  icache_io_ptw_invalidate;
  wire  icache_io_mem_acquire_ready;
  wire  icache_io_mem_acquire_valid;
  wire [25:0] icache_io_mem_acquire_bits_addr_block;
  wire [1:0] icache_io_mem_acquire_bits_client_xact_id;
  wire [2:0] icache_io_mem_acquire_bits_addr_beat;
  wire  icache_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] icache_io_mem_acquire_bits_a_type;
  wire [11:0] icache_io_mem_acquire_bits_union;
  wire [63:0] icache_io_mem_acquire_bits_data;
  wire  icache_io_mem_grant_ready;
  wire  icache_io_mem_grant_valid;
  wire [2:0] icache_io_mem_grant_bits_addr_beat;
  wire [1:0] icache_io_mem_grant_bits_client_xact_id;
  wire [2:0] icache_io_mem_grant_bits_manager_xact_id;
  wire  icache_io_mem_grant_bits_is_builtin_type;
  wire [3:0] icache_io_mem_grant_bits_g_type;
  wire [63:0] icache_io_mem_grant_bits_data;
  wire  HellaCache_3557_clk;
  wire  HellaCache_3557_reset;
  wire  HellaCache_3557_io_cpu_req_ready;
  wire  HellaCache_3557_io_cpu_req_valid;
  wire [39:0] HellaCache_3557_io_cpu_req_bits_addr;
  wire [8:0] HellaCache_3557_io_cpu_req_bits_tag;
  wire [4:0] HellaCache_3557_io_cpu_req_bits_cmd;
  wire [2:0] HellaCache_3557_io_cpu_req_bits_typ;
  wire  HellaCache_3557_io_cpu_req_bits_phys;
  wire [63:0] HellaCache_3557_io_cpu_req_bits_data;
  wire  HellaCache_3557_io_cpu_s1_kill;
  wire [63:0] HellaCache_3557_io_cpu_s1_data;
  wire  HellaCache_3557_io_cpu_s2_nack;
  wire  HellaCache_3557_io_cpu_resp_valid;
  wire [39:0] HellaCache_3557_io_cpu_resp_bits_addr;
  wire [8:0] HellaCache_3557_io_cpu_resp_bits_tag;
  wire [4:0] HellaCache_3557_io_cpu_resp_bits_cmd;
  wire [2:0] HellaCache_3557_io_cpu_resp_bits_typ;
  wire [63:0] HellaCache_3557_io_cpu_resp_bits_data;
  wire  HellaCache_3557_io_cpu_resp_bits_replay;
  wire  HellaCache_3557_io_cpu_resp_bits_has_data;
  wire [63:0] HellaCache_3557_io_cpu_resp_bits_data_word_bypass;
  wire [63:0] HellaCache_3557_io_cpu_resp_bits_store_data;
  wire  HellaCache_3557_io_cpu_replay_next;
  wire  HellaCache_3557_io_cpu_xcpt_ma_ld;
  wire  HellaCache_3557_io_cpu_xcpt_ma_st;
  wire  HellaCache_3557_io_cpu_xcpt_pf_ld;
  wire  HellaCache_3557_io_cpu_xcpt_pf_st;
  wire  HellaCache_3557_io_cpu_invalidate_lr;
  wire  HellaCache_3557_io_cpu_ordered;
  wire  HellaCache_3557_io_ptw_req_ready;
  wire  HellaCache_3557_io_ptw_req_valid;
  wire [26:0] HellaCache_3557_io_ptw_req_bits_addr;
  wire [1:0] HellaCache_3557_io_ptw_req_bits_prv;
  wire  HellaCache_3557_io_ptw_req_bits_store;
  wire  HellaCache_3557_io_ptw_req_bits_fetch;
  wire  HellaCache_3557_io_ptw_resp_valid;
  wire [19:0] HellaCache_3557_io_ptw_resp_bits_pte_ppn;
  wire [2:0] HellaCache_3557_io_ptw_resp_bits_pte_reserved_for_software;
  wire  HellaCache_3557_io_ptw_resp_bits_pte_d;
  wire  HellaCache_3557_io_ptw_resp_bits_pte_r;
  wire [3:0] HellaCache_3557_io_ptw_resp_bits_pte_typ;
  wire  HellaCache_3557_io_ptw_resp_bits_pte_v;
  wire  HellaCache_3557_io_ptw_status_debug;
  wire [1:0] HellaCache_3557_io_ptw_status_prv;
  wire  HellaCache_3557_io_ptw_status_sd;
  wire [30:0] HellaCache_3557_io_ptw_status_zero3;
  wire  HellaCache_3557_io_ptw_status_sd_rv32;
  wire [1:0] HellaCache_3557_io_ptw_status_zero2;
  wire [4:0] HellaCache_3557_io_ptw_status_vm;
  wire [4:0] HellaCache_3557_io_ptw_status_zero1;
  wire  HellaCache_3557_io_ptw_status_pum;
  wire  HellaCache_3557_io_ptw_status_mprv;
  wire [1:0] HellaCache_3557_io_ptw_status_xs;
  wire [1:0] HellaCache_3557_io_ptw_status_fs;
  wire [1:0] HellaCache_3557_io_ptw_status_mpp;
  wire [1:0] HellaCache_3557_io_ptw_status_hpp;
  wire  HellaCache_3557_io_ptw_status_spp;
  wire  HellaCache_3557_io_ptw_status_mpie;
  wire  HellaCache_3557_io_ptw_status_hpie;
  wire  HellaCache_3557_io_ptw_status_spie;
  wire  HellaCache_3557_io_ptw_status_upie;
  wire  HellaCache_3557_io_ptw_status_mie;
  wire  HellaCache_3557_io_ptw_status_hie;
  wire  HellaCache_3557_io_ptw_status_sie;
  wire  HellaCache_3557_io_ptw_status_uie;
  wire  HellaCache_3557_io_ptw_invalidate;
  wire  HellaCache_3557_io_mem_acquire_ready;
  wire  HellaCache_3557_io_mem_acquire_valid;
  wire [25:0] HellaCache_3557_io_mem_acquire_bits_addr_block;
  wire [1:0] HellaCache_3557_io_mem_acquire_bits_client_xact_id;
  wire [2:0] HellaCache_3557_io_mem_acquire_bits_addr_beat;
  wire  HellaCache_3557_io_mem_acquire_bits_is_builtin_type;
  wire [2:0] HellaCache_3557_io_mem_acquire_bits_a_type;
  wire [11:0] HellaCache_3557_io_mem_acquire_bits_union;
  wire [63:0] HellaCache_3557_io_mem_acquire_bits_data;
  wire  HellaCache_3557_io_mem_probe_ready;
  wire  HellaCache_3557_io_mem_probe_valid;
  wire [25:0] HellaCache_3557_io_mem_probe_bits_addr_block;
  wire [1:0] HellaCache_3557_io_mem_probe_bits_p_type;
  wire  HellaCache_3557_io_mem_release_ready;
  wire  HellaCache_3557_io_mem_release_valid;
  wire [2:0] HellaCache_3557_io_mem_release_bits_addr_beat;
  wire [25:0] HellaCache_3557_io_mem_release_bits_addr_block;
  wire [1:0] HellaCache_3557_io_mem_release_bits_client_xact_id;
  wire  HellaCache_3557_io_mem_release_bits_voluntary;
  wire [2:0] HellaCache_3557_io_mem_release_bits_r_type;
  wire [63:0] HellaCache_3557_io_mem_release_bits_data;
  wire  HellaCache_3557_io_mem_grant_ready;
  wire  HellaCache_3557_io_mem_grant_valid;
  wire [2:0] HellaCache_3557_io_mem_grant_bits_addr_beat;
  wire [1:0] HellaCache_3557_io_mem_grant_bits_client_xact_id;
  wire [2:0] HellaCache_3557_io_mem_grant_bits_manager_xact_id;
  wire  HellaCache_3557_io_mem_grant_bits_is_builtin_type;
  wire [3:0] HellaCache_3557_io_mem_grant_bits_g_type;
  wire [63:0] HellaCache_3557_io_mem_grant_bits_data;
  wire  HellaCache_3557_io_mem_grant_bits_manager_id;
  wire  HellaCache_3557_io_mem_finish_ready;
  wire  HellaCache_3557_io_mem_finish_valid;
  wire [2:0] HellaCache_3557_io_mem_finish_bits_manager_xact_id;
  wire  HellaCache_3557_io_mem_finish_bits_manager_id;
  wire  FPU_3558_clk;
  wire  FPU_3558_reset;
  wire [31:0] FPU_3558_io_inst;
  wire [63:0] FPU_3558_io_fromint_data;
  wire [2:0] FPU_3558_io_fcsr_rm;
  wire  FPU_3558_io_fcsr_flags_valid;
  wire [4:0] FPU_3558_io_fcsr_flags_bits;
  wire [63:0] FPU_3558_io_store_data;
  wire [63:0] FPU_3558_io_toint_data;
  wire  FPU_3558_io_dmem_resp_val;
  wire [2:0] FPU_3558_io_dmem_resp_type;
  wire [4:0] FPU_3558_io_dmem_resp_tag;
  wire [63:0] FPU_3558_io_dmem_resp_data;
  wire  FPU_3558_io_valid;
  wire  FPU_3558_io_fcsr_rdy;
  wire  FPU_3558_io_nack_mem;
  wire  FPU_3558_io_illegal_rm;
  wire  FPU_3558_io_killx;
  wire  FPU_3558_io_killm;
  wire [4:0] FPU_3558_io_dec_cmd;
  wire  FPU_3558_io_dec_ldst;
  wire  FPU_3558_io_dec_wen;
  wire  FPU_3558_io_dec_ren1;
  wire  FPU_3558_io_dec_ren2;
  wire  FPU_3558_io_dec_ren3;
  wire  FPU_3558_io_dec_swap12;
  wire  FPU_3558_io_dec_swap23;
  wire  FPU_3558_io_dec_single;
  wire  FPU_3558_io_dec_fromint;
  wire  FPU_3558_io_dec_toint;
  wire  FPU_3558_io_dec_fastpipe;
  wire  FPU_3558_io_dec_fma;
  wire  FPU_3558_io_dec_div;
  wire  FPU_3558_io_dec_sqrt;
  wire  FPU_3558_io_dec_round;
  wire  FPU_3558_io_dec_wflags;
  wire  FPU_3558_io_sboard_set;
  wire  FPU_3558_io_sboard_clr;
  wire [4:0] FPU_3558_io_sboard_clra;
  wire  FPU_3558_io_cp_req_ready;
  wire  FPU_3558_io_cp_req_valid;
  wire [4:0] FPU_3558_io_cp_req_bits_cmd;
  wire  FPU_3558_io_cp_req_bits_ldst;
  wire  FPU_3558_io_cp_req_bits_wen;
  wire  FPU_3558_io_cp_req_bits_ren1;
  wire  FPU_3558_io_cp_req_bits_ren2;
  wire  FPU_3558_io_cp_req_bits_ren3;
  wire  FPU_3558_io_cp_req_bits_swap12;
  wire  FPU_3558_io_cp_req_bits_swap23;
  wire  FPU_3558_io_cp_req_bits_single;
  wire  FPU_3558_io_cp_req_bits_fromint;
  wire  FPU_3558_io_cp_req_bits_toint;
  wire  FPU_3558_io_cp_req_bits_fastpipe;
  wire  FPU_3558_io_cp_req_bits_fma;
  wire  FPU_3558_io_cp_req_bits_div;
  wire  FPU_3558_io_cp_req_bits_sqrt;
  wire  FPU_3558_io_cp_req_bits_round;
  wire  FPU_3558_io_cp_req_bits_wflags;
  wire [2:0] FPU_3558_io_cp_req_bits_rm;
  wire [1:0] FPU_3558_io_cp_req_bits_typ;
  wire [64:0] FPU_3558_io_cp_req_bits_in1;
  wire [64:0] FPU_3558_io_cp_req_bits_in2;
  wire [64:0] FPU_3558_io_cp_req_bits_in3;
  wire  FPU_3558_io_cp_resp_ready;
  wire  FPU_3558_io_cp_resp_valid;
  wire [64:0] FPU_3558_io_cp_resp_bits_data;
  wire [4:0] FPU_3558_io_cp_resp_bits_exc;
  wire  uncachedArb_clk;
  wire  uncachedArb_reset;
  wire  uncachedArb_io_in_0_acquire_ready;
  wire  uncachedArb_io_in_0_acquire_valid;
  wire [25:0] uncachedArb_io_in_0_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_in_0_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_addr_beat;
  wire  uncachedArb_io_in_0_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_in_0_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_in_0_acquire_bits_union;
  wire [63:0] uncachedArb_io_in_0_acquire_bits_data;
  wire  uncachedArb_io_in_0_grant_ready;
  wire  uncachedArb_io_in_0_grant_valid;
  wire [2:0] uncachedArb_io_in_0_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_in_0_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_in_0_grant_bits_manager_xact_id;
  wire  uncachedArb_io_in_0_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_in_0_grant_bits_g_type;
  wire [63:0] uncachedArb_io_in_0_grant_bits_data;
  wire  uncachedArb_io_out_acquire_ready;
  wire  uncachedArb_io_out_acquire_valid;
  wire [25:0] uncachedArb_io_out_acquire_bits_addr_block;
  wire [1:0] uncachedArb_io_out_acquire_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_acquire_bits_addr_beat;
  wire  uncachedArb_io_out_acquire_bits_is_builtin_type;
  wire [2:0] uncachedArb_io_out_acquire_bits_a_type;
  wire [11:0] uncachedArb_io_out_acquire_bits_union;
  wire [63:0] uncachedArb_io_out_acquire_bits_data;
  wire  uncachedArb_io_out_grant_ready;
  wire  uncachedArb_io_out_grant_valid;
  wire [2:0] uncachedArb_io_out_grant_bits_addr_beat;
  wire [1:0] uncachedArb_io_out_grant_bits_client_xact_id;
  wire [2:0] uncachedArb_io_out_grant_bits_manager_xact_id;
  wire  uncachedArb_io_out_grant_bits_is_builtin_type;
  wire [3:0] uncachedArb_io_out_grant_bits_g_type;
  wire [63:0] uncachedArb_io_out_grant_bits_data;
  wire  PTW_3559_clk;
  wire  PTW_3559_reset;
  wire  PTW_3559_io_requestor_0_req_ready;
  wire  PTW_3559_io_requestor_0_req_valid;
  wire [26:0] PTW_3559_io_requestor_0_req_bits_addr;
  wire [1:0] PTW_3559_io_requestor_0_req_bits_prv;
  wire  PTW_3559_io_requestor_0_req_bits_store;
  wire  PTW_3559_io_requestor_0_req_bits_fetch;
  wire  PTW_3559_io_requestor_0_resp_valid;
  wire [19:0] PTW_3559_io_requestor_0_resp_bits_pte_ppn;
  wire [2:0] PTW_3559_io_requestor_0_resp_bits_pte_reserved_for_software;
  wire  PTW_3559_io_requestor_0_resp_bits_pte_d;
  wire  PTW_3559_io_requestor_0_resp_bits_pte_r;
  wire [3:0] PTW_3559_io_requestor_0_resp_bits_pte_typ;
  wire  PTW_3559_io_requestor_0_resp_bits_pte_v;
  wire  PTW_3559_io_requestor_0_status_debug;
  wire [1:0] PTW_3559_io_requestor_0_status_prv;
  wire  PTW_3559_io_requestor_0_status_sd;
  wire [30:0] PTW_3559_io_requestor_0_status_zero3;
  wire  PTW_3559_io_requestor_0_status_sd_rv32;
  wire [1:0] PTW_3559_io_requestor_0_status_zero2;
  wire [4:0] PTW_3559_io_requestor_0_status_vm;
  wire [4:0] PTW_3559_io_requestor_0_status_zero1;
  wire  PTW_3559_io_requestor_0_status_pum;
  wire  PTW_3559_io_requestor_0_status_mprv;
  wire [1:0] PTW_3559_io_requestor_0_status_xs;
  wire [1:0] PTW_3559_io_requestor_0_status_fs;
  wire [1:0] PTW_3559_io_requestor_0_status_mpp;
  wire [1:0] PTW_3559_io_requestor_0_status_hpp;
  wire  PTW_3559_io_requestor_0_status_spp;
  wire  PTW_3559_io_requestor_0_status_mpie;
  wire  PTW_3559_io_requestor_0_status_hpie;
  wire  PTW_3559_io_requestor_0_status_spie;
  wire  PTW_3559_io_requestor_0_status_upie;
  wire  PTW_3559_io_requestor_0_status_mie;
  wire  PTW_3559_io_requestor_0_status_hie;
  wire  PTW_3559_io_requestor_0_status_sie;
  wire  PTW_3559_io_requestor_0_status_uie;
  wire  PTW_3559_io_requestor_0_invalidate;
  wire  PTW_3559_io_requestor_1_req_ready;
  wire  PTW_3559_io_requestor_1_req_valid;
  wire [26:0] PTW_3559_io_requestor_1_req_bits_addr;
  wire [1:0] PTW_3559_io_requestor_1_req_bits_prv;
  wire  PTW_3559_io_requestor_1_req_bits_store;
  wire  PTW_3559_io_requestor_1_req_bits_fetch;
  wire  PTW_3559_io_requestor_1_resp_valid;
  wire [19:0] PTW_3559_io_requestor_1_resp_bits_pte_ppn;
  wire [2:0] PTW_3559_io_requestor_1_resp_bits_pte_reserved_for_software;
  wire  PTW_3559_io_requestor_1_resp_bits_pte_d;
  wire  PTW_3559_io_requestor_1_resp_bits_pte_r;
  wire [3:0] PTW_3559_io_requestor_1_resp_bits_pte_typ;
  wire  PTW_3559_io_requestor_1_resp_bits_pte_v;
  wire  PTW_3559_io_requestor_1_status_debug;
  wire [1:0] PTW_3559_io_requestor_1_status_prv;
  wire  PTW_3559_io_requestor_1_status_sd;
  wire [30:0] PTW_3559_io_requestor_1_status_zero3;
  wire  PTW_3559_io_requestor_1_status_sd_rv32;
  wire [1:0] PTW_3559_io_requestor_1_status_zero2;
  wire [4:0] PTW_3559_io_requestor_1_status_vm;
  wire [4:0] PTW_3559_io_requestor_1_status_zero1;
  wire  PTW_3559_io_requestor_1_status_pum;
  wire  PTW_3559_io_requestor_1_status_mprv;
  wire [1:0] PTW_3559_io_requestor_1_status_xs;
  wire [1:0] PTW_3559_io_requestor_1_status_fs;
  wire [1:0] PTW_3559_io_requestor_1_status_mpp;
  wire [1:0] PTW_3559_io_requestor_1_status_hpp;
  wire  PTW_3559_io_requestor_1_status_spp;
  wire  PTW_3559_io_requestor_1_status_mpie;
  wire  PTW_3559_io_requestor_1_status_hpie;
  wire  PTW_3559_io_requestor_1_status_spie;
  wire  PTW_3559_io_requestor_1_status_upie;
  wire  PTW_3559_io_requestor_1_status_mie;
  wire  PTW_3559_io_requestor_1_status_hie;
  wire  PTW_3559_io_requestor_1_status_sie;
  wire  PTW_3559_io_requestor_1_status_uie;
  wire  PTW_3559_io_requestor_1_invalidate;
  wire  PTW_3559_io_mem_req_ready;
  wire  PTW_3559_io_mem_req_valid;
  wire [39:0] PTW_3559_io_mem_req_bits_addr;
  wire [8:0] PTW_3559_io_mem_req_bits_tag;
  wire [4:0] PTW_3559_io_mem_req_bits_cmd;
  wire [2:0] PTW_3559_io_mem_req_bits_typ;
  wire  PTW_3559_io_mem_req_bits_phys;
  wire [63:0] PTW_3559_io_mem_req_bits_data;
  wire  PTW_3559_io_mem_s1_kill;
  wire [63:0] PTW_3559_io_mem_s1_data;
  wire  PTW_3559_io_mem_s2_nack;
  wire  PTW_3559_io_mem_resp_valid;
  wire [39:0] PTW_3559_io_mem_resp_bits_addr;
  wire [8:0] PTW_3559_io_mem_resp_bits_tag;
  wire [4:0] PTW_3559_io_mem_resp_bits_cmd;
  wire [2:0] PTW_3559_io_mem_resp_bits_typ;
  wire [63:0] PTW_3559_io_mem_resp_bits_data;
  wire  PTW_3559_io_mem_resp_bits_replay;
  wire  PTW_3559_io_mem_resp_bits_has_data;
  wire [63:0] PTW_3559_io_mem_resp_bits_data_word_bypass;
  wire [63:0] PTW_3559_io_mem_resp_bits_store_data;
  wire  PTW_3559_io_mem_replay_next;
  wire  PTW_3559_io_mem_xcpt_ma_ld;
  wire  PTW_3559_io_mem_xcpt_ma_st;
  wire  PTW_3559_io_mem_xcpt_pf_ld;
  wire  PTW_3559_io_mem_xcpt_pf_st;
  wire  PTW_3559_io_mem_invalidate_lr;
  wire  PTW_3559_io_mem_ordered;
  wire [19:0] PTW_3559_io_dpath_ptbr;
  wire  PTW_3559_io_dpath_invalidate;
  wire  PTW_3559_io_dpath_status_debug;
  wire [1:0] PTW_3559_io_dpath_status_prv;
  wire  PTW_3559_io_dpath_status_sd;
  wire [30:0] PTW_3559_io_dpath_status_zero3;
  wire  PTW_3559_io_dpath_status_sd_rv32;
  wire [1:0] PTW_3559_io_dpath_status_zero2;
  wire [4:0] PTW_3559_io_dpath_status_vm;
  wire [4:0] PTW_3559_io_dpath_status_zero1;
  wire  PTW_3559_io_dpath_status_pum;
  wire  PTW_3559_io_dpath_status_mprv;
  wire [1:0] PTW_3559_io_dpath_status_xs;
  wire [1:0] PTW_3559_io_dpath_status_fs;
  wire [1:0] PTW_3559_io_dpath_status_mpp;
  wire [1:0] PTW_3559_io_dpath_status_hpp;
  wire  PTW_3559_io_dpath_status_spp;
  wire  PTW_3559_io_dpath_status_mpie;
  wire  PTW_3559_io_dpath_status_hpie;
  wire  PTW_3559_io_dpath_status_spie;
  wire  PTW_3559_io_dpath_status_upie;
  wire  PTW_3559_io_dpath_status_mie;
  wire  PTW_3559_io_dpath_status_hie;
  wire  PTW_3559_io_dpath_status_sie;
  wire  PTW_3559_io_dpath_status_uie;
  wire  dcArb_clk;
  wire  dcArb_reset;
  wire  dcArb_io_requestor_0_req_ready;
  wire  dcArb_io_requestor_0_req_valid;
  wire [39:0] dcArb_io_requestor_0_req_bits_addr;
  wire [8:0] dcArb_io_requestor_0_req_bits_tag;
  wire [4:0] dcArb_io_requestor_0_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_req_bits_typ;
  wire  dcArb_io_requestor_0_req_bits_phys;
  wire [63:0] dcArb_io_requestor_0_req_bits_data;
  wire  dcArb_io_requestor_0_s1_kill;
  wire [63:0] dcArb_io_requestor_0_s1_data;
  wire  dcArb_io_requestor_0_s2_nack;
  wire  dcArb_io_requestor_0_resp_valid;
  wire [39:0] dcArb_io_requestor_0_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_0_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_0_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_0_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data;
  wire  dcArb_io_requestor_0_resp_bits_replay;
  wire  dcArb_io_requestor_0_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_0_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_0_resp_bits_store_data;
  wire  dcArb_io_requestor_0_replay_next;
  wire  dcArb_io_requestor_0_xcpt_ma_ld;
  wire  dcArb_io_requestor_0_xcpt_ma_st;
  wire  dcArb_io_requestor_0_xcpt_pf_ld;
  wire  dcArb_io_requestor_0_xcpt_pf_st;
  wire  dcArb_io_requestor_0_invalidate_lr;
  wire  dcArb_io_requestor_0_ordered;
  wire  dcArb_io_requestor_1_req_ready;
  wire  dcArb_io_requestor_1_req_valid;
  wire [39:0] dcArb_io_requestor_1_req_bits_addr;
  wire [8:0] dcArb_io_requestor_1_req_bits_tag;
  wire [4:0] dcArb_io_requestor_1_req_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_req_bits_typ;
  wire  dcArb_io_requestor_1_req_bits_phys;
  wire [63:0] dcArb_io_requestor_1_req_bits_data;
  wire  dcArb_io_requestor_1_s1_kill;
  wire [63:0] dcArb_io_requestor_1_s1_data;
  wire  dcArb_io_requestor_1_s2_nack;
  wire  dcArb_io_requestor_1_resp_valid;
  wire [39:0] dcArb_io_requestor_1_resp_bits_addr;
  wire [8:0] dcArb_io_requestor_1_resp_bits_tag;
  wire [4:0] dcArb_io_requestor_1_resp_bits_cmd;
  wire [2:0] dcArb_io_requestor_1_resp_bits_typ;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data;
  wire  dcArb_io_requestor_1_resp_bits_replay;
  wire  dcArb_io_requestor_1_resp_bits_has_data;
  wire [63:0] dcArb_io_requestor_1_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_requestor_1_resp_bits_store_data;
  wire  dcArb_io_requestor_1_replay_next;
  wire  dcArb_io_requestor_1_xcpt_ma_ld;
  wire  dcArb_io_requestor_1_xcpt_ma_st;
  wire  dcArb_io_requestor_1_xcpt_pf_ld;
  wire  dcArb_io_requestor_1_xcpt_pf_st;
  wire  dcArb_io_requestor_1_invalidate_lr;
  wire  dcArb_io_requestor_1_ordered;
  wire  dcArb_io_mem_req_ready;
  wire  dcArb_io_mem_req_valid;
  wire [39:0] dcArb_io_mem_req_bits_addr;
  wire [8:0] dcArb_io_mem_req_bits_tag;
  wire [4:0] dcArb_io_mem_req_bits_cmd;
  wire [2:0] dcArb_io_mem_req_bits_typ;
  wire  dcArb_io_mem_req_bits_phys;
  wire [63:0] dcArb_io_mem_req_bits_data;
  wire  dcArb_io_mem_s1_kill;
  wire [63:0] dcArb_io_mem_s1_data;
  wire  dcArb_io_mem_s2_nack;
  wire  dcArb_io_mem_resp_valid;
  wire [39:0] dcArb_io_mem_resp_bits_addr;
  wire [8:0] dcArb_io_mem_resp_bits_tag;
  wire [4:0] dcArb_io_mem_resp_bits_cmd;
  wire [2:0] dcArb_io_mem_resp_bits_typ;
  wire [63:0] dcArb_io_mem_resp_bits_data;
  wire  dcArb_io_mem_resp_bits_replay;
  wire  dcArb_io_mem_resp_bits_has_data;
  wire [63:0] dcArb_io_mem_resp_bits_data_word_bypass;
  wire [63:0] dcArb_io_mem_resp_bits_store_data;
  wire  dcArb_io_mem_replay_next;
  wire  dcArb_io_mem_xcpt_ma_ld;
  wire  dcArb_io_mem_xcpt_ma_st;
  wire  dcArb_io_mem_xcpt_pf_ld;
  wire  dcArb_io_mem_xcpt_pf_st;
  wire  dcArb_io_mem_invalidate_lr;
  wire  dcArb_io_mem_ordered;
  reg  GEN_0;
  reg [31:0] GEN_58;
  reg [1:0] GEN_1;
  reg [31:0] GEN_59;
  reg  GEN_2;
  reg [31:0] GEN_60;
  reg [2:0] GEN_3;
  reg [31:0] GEN_61;
  reg [31:0] GEN_4;
  reg [31:0] GEN_62;
  reg [31:0] GEN_5;
  reg [31:0] GEN_63;
  reg [31:0] GEN_6;
  reg [31:0] GEN_64;
  reg [1:0] GEN_7;
  reg [31:0] GEN_65;
  reg  GEN_8;
  reg [31:0] GEN_66;
  reg  GEN_9;
  reg [31:0] GEN_67;
  reg  GEN_10;
  reg [31:0] GEN_68;
  reg [4:0] GEN_11;
  reg [31:0] GEN_69;
  reg [63:0] GEN_12;
  reg [63:0] GEN_70;
  reg  GEN_13;
  reg [31:0] GEN_71;
  reg [39:0] GEN_14;
  reg [63:0] GEN_72;
  reg [8:0] GEN_15;
  reg [31:0] GEN_73;
  reg [4:0] GEN_16;
  reg [31:0] GEN_74;
  reg [2:0] GEN_17;
  reg [31:0] GEN_75;
  reg  GEN_18;
  reg [31:0] GEN_76;
  reg [63:0] GEN_19;
  reg [63:0] GEN_77;
  reg  GEN_20;
  reg [31:0] GEN_78;
  reg [63:0] GEN_21;
  reg [63:0] GEN_79;
  reg  GEN_22;
  reg [31:0] GEN_80;
  reg  GEN_23;
  reg [31:0] GEN_81;
  reg  GEN_24;
  reg [31:0] GEN_82;
  reg  GEN_25;
  reg [31:0] GEN_83;
  reg [25:0] GEN_26;
  reg [31:0] GEN_84;
  reg [1:0] GEN_27;
  reg [31:0] GEN_85;
  reg [2:0] GEN_28;
  reg [31:0] GEN_86;
  reg  GEN_29;
  reg [31:0] GEN_87;
  reg [2:0] GEN_30;
  reg [31:0] GEN_88;
  reg [11:0] GEN_31;
  reg [31:0] GEN_89;
  reg [63:0] GEN_32;
  reg [63:0] GEN_90;
  reg  GEN_33;
  reg [31:0] GEN_91;
  reg  GEN_34;
  reg [31:0] GEN_92;
  reg [4:0] GEN_35;
  reg [31:0] GEN_93;
  reg  GEN_36;
  reg [31:0] GEN_94;
  reg  GEN_37;
  reg [31:0] GEN_95;
  reg  GEN_38;
  reg [31:0] GEN_96;
  reg  GEN_39;
  reg [31:0] GEN_97;
  reg  GEN_40;
  reg [31:0] GEN_98;
  reg  GEN_41;
  reg [31:0] GEN_99;
  reg  GEN_42;
  reg [31:0] GEN_100;
  reg  GEN_43;
  reg [31:0] GEN_101;
  reg  GEN_44;
  reg [31:0] GEN_102;
  reg  GEN_45;
  reg [31:0] GEN_103;
  reg  GEN_46;
  reg [31:0] GEN_104;
  reg  GEN_47;
  reg [31:0] GEN_105;
  reg  GEN_48;
  reg [31:0] GEN_106;
  reg  GEN_49;
  reg [31:0] GEN_107;
  reg  GEN_50;
  reg [31:0] GEN_108;
  reg  GEN_51;
  reg [31:0] GEN_109;
  reg [2:0] GEN_52;
  reg [31:0] GEN_110;
  reg [1:0] GEN_53;
  reg [31:0] GEN_111;
  reg [64:0] GEN_54;
  reg [95:0] GEN_112;
  reg [64:0] GEN_55;
  reg [95:0] GEN_113;
  reg [64:0] GEN_56;
  reg [95:0] GEN_114;
  reg  GEN_57;
  reg [31:0] GEN_115;
  Rocket core (
    .clk(core_clk),
    .reset(core_reset),
    .io_prci_reset(core_io_prci_reset),
    .io_prci_id(core_io_prci_id),
    .io_prci_interrupts_mtip(core_io_prci_interrupts_mtip),
    .io_prci_interrupts_meip(core_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(core_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(core_io_prci_interrupts_debug),
    .io_prci_interrupts_msip(core_io_prci_interrupts_msip),
    .io_imem_req_valid(core_io_imem_req_valid),
    .io_imem_req_bits_pc(core_io_imem_req_bits_pc),
    .io_imem_resp_ready(core_io_imem_resp_ready),
    .io_imem_resp_valid(core_io_imem_resp_valid),
    .io_imem_resp_bits_pc(core_io_imem_resp_bits_pc),
    .io_imem_resp_bits_data_0(core_io_imem_resp_bits_data_0),
    .io_imem_resp_bits_mask(core_io_imem_resp_bits_mask),
    .io_imem_resp_bits_xcpt_if(core_io_imem_resp_bits_xcpt_if),
    .io_imem_btb_resp_valid(core_io_imem_btb_resp_valid),
    .io_imem_btb_resp_bits_taken(core_io_imem_btb_resp_bits_taken),
    .io_imem_btb_resp_bits_mask(core_io_imem_btb_resp_bits_mask),
    .io_imem_btb_resp_bits_bridx(core_io_imem_btb_resp_bits_bridx),
    .io_imem_btb_resp_bits_target(core_io_imem_btb_resp_bits_target),
    .io_imem_btb_resp_bits_entry(core_io_imem_btb_resp_bits_entry),
    .io_imem_btb_resp_bits_bht_history(core_io_imem_btb_resp_bits_bht_history),
    .io_imem_btb_resp_bits_bht_value(core_io_imem_btb_resp_bits_bht_value),
    .io_imem_btb_update_valid(core_io_imem_btb_update_valid),
    .io_imem_btb_update_bits_prediction_valid(core_io_imem_btb_update_bits_prediction_valid),
    .io_imem_btb_update_bits_prediction_bits_taken(core_io_imem_btb_update_bits_prediction_bits_taken),
    .io_imem_btb_update_bits_prediction_bits_mask(core_io_imem_btb_update_bits_prediction_bits_mask),
    .io_imem_btb_update_bits_prediction_bits_bridx(core_io_imem_btb_update_bits_prediction_bits_bridx),
    .io_imem_btb_update_bits_prediction_bits_target(core_io_imem_btb_update_bits_prediction_bits_target),
    .io_imem_btb_update_bits_prediction_bits_entry(core_io_imem_btb_update_bits_prediction_bits_entry),
    .io_imem_btb_update_bits_prediction_bits_bht_history(core_io_imem_btb_update_bits_prediction_bits_bht_history),
    .io_imem_btb_update_bits_prediction_bits_bht_value(core_io_imem_btb_update_bits_prediction_bits_bht_value),
    .io_imem_btb_update_bits_pc(core_io_imem_btb_update_bits_pc),
    .io_imem_btb_update_bits_target(core_io_imem_btb_update_bits_target),
    .io_imem_btb_update_bits_taken(core_io_imem_btb_update_bits_taken),
    .io_imem_btb_update_bits_isJump(core_io_imem_btb_update_bits_isJump),
    .io_imem_btb_update_bits_isReturn(core_io_imem_btb_update_bits_isReturn),
    .io_imem_btb_update_bits_br_pc(core_io_imem_btb_update_bits_br_pc),
    .io_imem_bht_update_valid(core_io_imem_bht_update_valid),
    .io_imem_bht_update_bits_prediction_valid(core_io_imem_bht_update_bits_prediction_valid),
    .io_imem_bht_update_bits_prediction_bits_taken(core_io_imem_bht_update_bits_prediction_bits_taken),
    .io_imem_bht_update_bits_prediction_bits_mask(core_io_imem_bht_update_bits_prediction_bits_mask),
    .io_imem_bht_update_bits_prediction_bits_bridx(core_io_imem_bht_update_bits_prediction_bits_bridx),
    .io_imem_bht_update_bits_prediction_bits_target(core_io_imem_bht_update_bits_prediction_bits_target),
    .io_imem_bht_update_bits_prediction_bits_entry(core_io_imem_bht_update_bits_prediction_bits_entry),
    .io_imem_bht_update_bits_prediction_bits_bht_history(core_io_imem_bht_update_bits_prediction_bits_bht_history),
    .io_imem_bht_update_bits_prediction_bits_bht_value(core_io_imem_bht_update_bits_prediction_bits_bht_value),
    .io_imem_bht_update_bits_pc(core_io_imem_bht_update_bits_pc),
    .io_imem_bht_update_bits_taken(core_io_imem_bht_update_bits_taken),
    .io_imem_bht_update_bits_mispredict(core_io_imem_bht_update_bits_mispredict),
    .io_imem_ras_update_valid(core_io_imem_ras_update_valid),
    .io_imem_ras_update_bits_isCall(core_io_imem_ras_update_bits_isCall),
    .io_imem_ras_update_bits_isReturn(core_io_imem_ras_update_bits_isReturn),
    .io_imem_ras_update_bits_returnAddr(core_io_imem_ras_update_bits_returnAddr),
    .io_imem_ras_update_bits_prediction_valid(core_io_imem_ras_update_bits_prediction_valid),
    .io_imem_ras_update_bits_prediction_bits_taken(core_io_imem_ras_update_bits_prediction_bits_taken),
    .io_imem_ras_update_bits_prediction_bits_mask(core_io_imem_ras_update_bits_prediction_bits_mask),
    .io_imem_ras_update_bits_prediction_bits_bridx(core_io_imem_ras_update_bits_prediction_bits_bridx),
    .io_imem_ras_update_bits_prediction_bits_target(core_io_imem_ras_update_bits_prediction_bits_target),
    .io_imem_ras_update_bits_prediction_bits_entry(core_io_imem_ras_update_bits_prediction_bits_entry),
    .io_imem_ras_update_bits_prediction_bits_bht_history(core_io_imem_ras_update_bits_prediction_bits_bht_history),
    .io_imem_ras_update_bits_prediction_bits_bht_value(core_io_imem_ras_update_bits_prediction_bits_bht_value),
    .io_imem_flush_icache(core_io_imem_flush_icache),
    .io_imem_flush_tlb(core_io_imem_flush_tlb),
    .io_imem_npc(core_io_imem_npc),
    .io_dmem_req_ready(core_io_dmem_req_ready),
    .io_dmem_req_valid(core_io_dmem_req_valid),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_tag(core_io_dmem_req_bits_tag),
    .io_dmem_req_bits_cmd(core_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_req_bits_phys(core_io_dmem_req_bits_phys),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_s1_kill(core_io_dmem_s1_kill),
    .io_dmem_s1_data(core_io_dmem_s1_data),
    .io_dmem_s2_nack(core_io_dmem_s2_nack),
    .io_dmem_resp_valid(core_io_dmem_resp_valid),
    .io_dmem_resp_bits_addr(core_io_dmem_resp_bits_addr),
    .io_dmem_resp_bits_tag(core_io_dmem_resp_bits_tag),
    .io_dmem_resp_bits_cmd(core_io_dmem_resp_bits_cmd),
    .io_dmem_resp_bits_typ(core_io_dmem_resp_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    .io_dmem_resp_bits_replay(core_io_dmem_resp_bits_replay),
    .io_dmem_resp_bits_has_data(core_io_dmem_resp_bits_has_data),
    .io_dmem_resp_bits_data_word_bypass(core_io_dmem_resp_bits_data_word_bypass),
    .io_dmem_resp_bits_store_data(core_io_dmem_resp_bits_store_data),
    .io_dmem_replay_next(core_io_dmem_replay_next),
    .io_dmem_xcpt_ma_ld(core_io_dmem_xcpt_ma_ld),
    .io_dmem_xcpt_ma_st(core_io_dmem_xcpt_ma_st),
    .io_dmem_xcpt_pf_ld(core_io_dmem_xcpt_pf_ld),
    .io_dmem_xcpt_pf_st(core_io_dmem_xcpt_pf_st),
    .io_dmem_invalidate_lr(core_io_dmem_invalidate_lr),
    .io_dmem_ordered(core_io_dmem_ordered),
    .io_ptw_ptbr(core_io_ptw_ptbr),
    .io_ptw_invalidate(core_io_ptw_invalidate),
    .io_ptw_status_debug(core_io_ptw_status_debug),
    .io_ptw_status_prv(core_io_ptw_status_prv),
    .io_ptw_status_sd(core_io_ptw_status_sd),
    .io_ptw_status_zero3(core_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(core_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(core_io_ptw_status_zero2),
    .io_ptw_status_vm(core_io_ptw_status_vm),
    .io_ptw_status_zero1(core_io_ptw_status_zero1),
    .io_ptw_status_pum(core_io_ptw_status_pum),
    .io_ptw_status_mprv(core_io_ptw_status_mprv),
    .io_ptw_status_xs(core_io_ptw_status_xs),
    .io_ptw_status_fs(core_io_ptw_status_fs),
    .io_ptw_status_mpp(core_io_ptw_status_mpp),
    .io_ptw_status_hpp(core_io_ptw_status_hpp),
    .io_ptw_status_spp(core_io_ptw_status_spp),
    .io_ptw_status_mpie(core_io_ptw_status_mpie),
    .io_ptw_status_hpie(core_io_ptw_status_hpie),
    .io_ptw_status_spie(core_io_ptw_status_spie),
    .io_ptw_status_upie(core_io_ptw_status_upie),
    .io_ptw_status_mie(core_io_ptw_status_mie),
    .io_ptw_status_hie(core_io_ptw_status_hie),
    .io_ptw_status_sie(core_io_ptw_status_sie),
    .io_ptw_status_uie(core_io_ptw_status_uie),
    .io_fpu_inst(core_io_fpu_inst),
    .io_fpu_fromint_data(core_io_fpu_fromint_data),
    .io_fpu_fcsr_rm(core_io_fpu_fcsr_rm),
    .io_fpu_fcsr_flags_valid(core_io_fpu_fcsr_flags_valid),
    .io_fpu_fcsr_flags_bits(core_io_fpu_fcsr_flags_bits),
    .io_fpu_store_data(core_io_fpu_store_data),
    .io_fpu_toint_data(core_io_fpu_toint_data),
    .io_fpu_dmem_resp_val(core_io_fpu_dmem_resp_val),
    .io_fpu_dmem_resp_type(core_io_fpu_dmem_resp_type),
    .io_fpu_dmem_resp_tag(core_io_fpu_dmem_resp_tag),
    .io_fpu_dmem_resp_data(core_io_fpu_dmem_resp_data),
    .io_fpu_valid(core_io_fpu_valid),
    .io_fpu_fcsr_rdy(core_io_fpu_fcsr_rdy),
    .io_fpu_nack_mem(core_io_fpu_nack_mem),
    .io_fpu_illegal_rm(core_io_fpu_illegal_rm),
    .io_fpu_killx(core_io_fpu_killx),
    .io_fpu_killm(core_io_fpu_killm),
    .io_fpu_dec_cmd(core_io_fpu_dec_cmd),
    .io_fpu_dec_ldst(core_io_fpu_dec_ldst),
    .io_fpu_dec_wen(core_io_fpu_dec_wen),
    .io_fpu_dec_ren1(core_io_fpu_dec_ren1),
    .io_fpu_dec_ren2(core_io_fpu_dec_ren2),
    .io_fpu_dec_ren3(core_io_fpu_dec_ren3),
    .io_fpu_dec_swap12(core_io_fpu_dec_swap12),
    .io_fpu_dec_swap23(core_io_fpu_dec_swap23),
    .io_fpu_dec_single(core_io_fpu_dec_single),
    .io_fpu_dec_fromint(core_io_fpu_dec_fromint),
    .io_fpu_dec_toint(core_io_fpu_dec_toint),
    .io_fpu_dec_fastpipe(core_io_fpu_dec_fastpipe),
    .io_fpu_dec_fma(core_io_fpu_dec_fma),
    .io_fpu_dec_div(core_io_fpu_dec_div),
    .io_fpu_dec_sqrt(core_io_fpu_dec_sqrt),
    .io_fpu_dec_round(core_io_fpu_dec_round),
    .io_fpu_dec_wflags(core_io_fpu_dec_wflags),
    .io_fpu_sboard_set(core_io_fpu_sboard_set),
    .io_fpu_sboard_clr(core_io_fpu_sboard_clr),
    .io_fpu_sboard_clra(core_io_fpu_sboard_clra),
    .io_fpu_cp_req_ready(core_io_fpu_cp_req_ready),
    .io_fpu_cp_req_valid(core_io_fpu_cp_req_valid),
    .io_fpu_cp_req_bits_cmd(core_io_fpu_cp_req_bits_cmd),
    .io_fpu_cp_req_bits_ldst(core_io_fpu_cp_req_bits_ldst),
    .io_fpu_cp_req_bits_wen(core_io_fpu_cp_req_bits_wen),
    .io_fpu_cp_req_bits_ren1(core_io_fpu_cp_req_bits_ren1),
    .io_fpu_cp_req_bits_ren2(core_io_fpu_cp_req_bits_ren2),
    .io_fpu_cp_req_bits_ren3(core_io_fpu_cp_req_bits_ren3),
    .io_fpu_cp_req_bits_swap12(core_io_fpu_cp_req_bits_swap12),
    .io_fpu_cp_req_bits_swap23(core_io_fpu_cp_req_bits_swap23),
    .io_fpu_cp_req_bits_single(core_io_fpu_cp_req_bits_single),
    .io_fpu_cp_req_bits_fromint(core_io_fpu_cp_req_bits_fromint),
    .io_fpu_cp_req_bits_toint(core_io_fpu_cp_req_bits_toint),
    .io_fpu_cp_req_bits_fastpipe(core_io_fpu_cp_req_bits_fastpipe),
    .io_fpu_cp_req_bits_fma(core_io_fpu_cp_req_bits_fma),
    .io_fpu_cp_req_bits_div(core_io_fpu_cp_req_bits_div),
    .io_fpu_cp_req_bits_sqrt(core_io_fpu_cp_req_bits_sqrt),
    .io_fpu_cp_req_bits_round(core_io_fpu_cp_req_bits_round),
    .io_fpu_cp_req_bits_wflags(core_io_fpu_cp_req_bits_wflags),
    .io_fpu_cp_req_bits_rm(core_io_fpu_cp_req_bits_rm),
    .io_fpu_cp_req_bits_typ(core_io_fpu_cp_req_bits_typ),
    .io_fpu_cp_req_bits_in1(core_io_fpu_cp_req_bits_in1),
    .io_fpu_cp_req_bits_in2(core_io_fpu_cp_req_bits_in2),
    .io_fpu_cp_req_bits_in3(core_io_fpu_cp_req_bits_in3),
    .io_fpu_cp_resp_ready(core_io_fpu_cp_resp_ready),
    .io_fpu_cp_resp_valid(core_io_fpu_cp_resp_valid),
    .io_fpu_cp_resp_bits_data(core_io_fpu_cp_resp_bits_data),
    .io_fpu_cp_resp_bits_exc(core_io_fpu_cp_resp_bits_exc),
    .io_rocc_cmd_ready(core_io_rocc_cmd_ready),
    .io_rocc_cmd_valid(core_io_rocc_cmd_valid),
    .io_rocc_cmd_bits_inst_funct(core_io_rocc_cmd_bits_inst_funct),
    .io_rocc_cmd_bits_inst_rs2(core_io_rocc_cmd_bits_inst_rs2),
    .io_rocc_cmd_bits_inst_rs1(core_io_rocc_cmd_bits_inst_rs1),
    .io_rocc_cmd_bits_inst_xd(core_io_rocc_cmd_bits_inst_xd),
    .io_rocc_cmd_bits_inst_xs1(core_io_rocc_cmd_bits_inst_xs1),
    .io_rocc_cmd_bits_inst_xs2(core_io_rocc_cmd_bits_inst_xs2),
    .io_rocc_cmd_bits_inst_rd(core_io_rocc_cmd_bits_inst_rd),
    .io_rocc_cmd_bits_inst_opcode(core_io_rocc_cmd_bits_inst_opcode),
    .io_rocc_cmd_bits_rs1(core_io_rocc_cmd_bits_rs1),
    .io_rocc_cmd_bits_rs2(core_io_rocc_cmd_bits_rs2),
    .io_rocc_resp_ready(core_io_rocc_resp_ready),
    .io_rocc_resp_valid(core_io_rocc_resp_valid),
    .io_rocc_resp_bits_rd(core_io_rocc_resp_bits_rd),
    .io_rocc_resp_bits_data(core_io_rocc_resp_bits_data),
    .io_rocc_mem_req_ready(core_io_rocc_mem_req_ready),
    .io_rocc_mem_req_valid(core_io_rocc_mem_req_valid),
    .io_rocc_mem_req_bits_addr(core_io_rocc_mem_req_bits_addr),
    .io_rocc_mem_req_bits_tag(core_io_rocc_mem_req_bits_tag),
    .io_rocc_mem_req_bits_cmd(core_io_rocc_mem_req_bits_cmd),
    .io_rocc_mem_req_bits_typ(core_io_rocc_mem_req_bits_typ),
    .io_rocc_mem_req_bits_phys(core_io_rocc_mem_req_bits_phys),
    .io_rocc_mem_req_bits_data(core_io_rocc_mem_req_bits_data),
    .io_rocc_mem_s1_kill(core_io_rocc_mem_s1_kill),
    .io_rocc_mem_s1_data(core_io_rocc_mem_s1_data),
    .io_rocc_mem_s2_nack(core_io_rocc_mem_s2_nack),
    .io_rocc_mem_resp_valid(core_io_rocc_mem_resp_valid),
    .io_rocc_mem_resp_bits_addr(core_io_rocc_mem_resp_bits_addr),
    .io_rocc_mem_resp_bits_tag(core_io_rocc_mem_resp_bits_tag),
    .io_rocc_mem_resp_bits_cmd(core_io_rocc_mem_resp_bits_cmd),
    .io_rocc_mem_resp_bits_typ(core_io_rocc_mem_resp_bits_typ),
    .io_rocc_mem_resp_bits_data(core_io_rocc_mem_resp_bits_data),
    .io_rocc_mem_resp_bits_replay(core_io_rocc_mem_resp_bits_replay),
    .io_rocc_mem_resp_bits_has_data(core_io_rocc_mem_resp_bits_has_data),
    .io_rocc_mem_resp_bits_data_word_bypass(core_io_rocc_mem_resp_bits_data_word_bypass),
    .io_rocc_mem_resp_bits_store_data(core_io_rocc_mem_resp_bits_store_data),
    .io_rocc_mem_replay_next(core_io_rocc_mem_replay_next),
    .io_rocc_mem_xcpt_ma_ld(core_io_rocc_mem_xcpt_ma_ld),
    .io_rocc_mem_xcpt_ma_st(core_io_rocc_mem_xcpt_ma_st),
    .io_rocc_mem_xcpt_pf_ld(core_io_rocc_mem_xcpt_pf_ld),
    .io_rocc_mem_xcpt_pf_st(core_io_rocc_mem_xcpt_pf_st),
    .io_rocc_mem_invalidate_lr(core_io_rocc_mem_invalidate_lr),
    .io_rocc_mem_ordered(core_io_rocc_mem_ordered),
    .io_rocc_busy(core_io_rocc_busy),
    .io_rocc_status_debug(core_io_rocc_status_debug),
    .io_rocc_status_prv(core_io_rocc_status_prv),
    .io_rocc_status_sd(core_io_rocc_status_sd),
    .io_rocc_status_zero3(core_io_rocc_status_zero3),
    .io_rocc_status_sd_rv32(core_io_rocc_status_sd_rv32),
    .io_rocc_status_zero2(core_io_rocc_status_zero2),
    .io_rocc_status_vm(core_io_rocc_status_vm),
    .io_rocc_status_zero1(core_io_rocc_status_zero1),
    .io_rocc_status_pum(core_io_rocc_status_pum),
    .io_rocc_status_mprv(core_io_rocc_status_mprv),
    .io_rocc_status_xs(core_io_rocc_status_xs),
    .io_rocc_status_fs(core_io_rocc_status_fs),
    .io_rocc_status_mpp(core_io_rocc_status_mpp),
    .io_rocc_status_hpp(core_io_rocc_status_hpp),
    .io_rocc_status_spp(core_io_rocc_status_spp),
    .io_rocc_status_mpie(core_io_rocc_status_mpie),
    .io_rocc_status_hpie(core_io_rocc_status_hpie),
    .io_rocc_status_spie(core_io_rocc_status_spie),
    .io_rocc_status_upie(core_io_rocc_status_upie),
    .io_rocc_status_mie(core_io_rocc_status_mie),
    .io_rocc_status_hie(core_io_rocc_status_hie),
    .io_rocc_status_sie(core_io_rocc_status_sie),
    .io_rocc_status_uie(core_io_rocc_status_uie),
    .io_rocc_interrupt(core_io_rocc_interrupt),
    .io_rocc_autl_acquire_ready(core_io_rocc_autl_acquire_ready),
    .io_rocc_autl_acquire_valid(core_io_rocc_autl_acquire_valid),
    .io_rocc_autl_acquire_bits_addr_block(core_io_rocc_autl_acquire_bits_addr_block),
    .io_rocc_autl_acquire_bits_client_xact_id(core_io_rocc_autl_acquire_bits_client_xact_id),
    .io_rocc_autl_acquire_bits_addr_beat(core_io_rocc_autl_acquire_bits_addr_beat),
    .io_rocc_autl_acquire_bits_is_builtin_type(core_io_rocc_autl_acquire_bits_is_builtin_type),
    .io_rocc_autl_acquire_bits_a_type(core_io_rocc_autl_acquire_bits_a_type),
    .io_rocc_autl_acquire_bits_union(core_io_rocc_autl_acquire_bits_union),
    .io_rocc_autl_acquire_bits_data(core_io_rocc_autl_acquire_bits_data),
    .io_rocc_autl_grant_ready(core_io_rocc_autl_grant_ready),
    .io_rocc_autl_grant_valid(core_io_rocc_autl_grant_valid),
    .io_rocc_autl_grant_bits_addr_beat(core_io_rocc_autl_grant_bits_addr_beat),
    .io_rocc_autl_grant_bits_client_xact_id(core_io_rocc_autl_grant_bits_client_xact_id),
    .io_rocc_autl_grant_bits_manager_xact_id(core_io_rocc_autl_grant_bits_manager_xact_id),
    .io_rocc_autl_grant_bits_is_builtin_type(core_io_rocc_autl_grant_bits_is_builtin_type),
    .io_rocc_autl_grant_bits_g_type(core_io_rocc_autl_grant_bits_g_type),
    .io_rocc_autl_grant_bits_data(core_io_rocc_autl_grant_bits_data),
    .io_rocc_fpu_req_ready(core_io_rocc_fpu_req_ready),
    .io_rocc_fpu_req_valid(core_io_rocc_fpu_req_valid),
    .io_rocc_fpu_req_bits_cmd(core_io_rocc_fpu_req_bits_cmd),
    .io_rocc_fpu_req_bits_ldst(core_io_rocc_fpu_req_bits_ldst),
    .io_rocc_fpu_req_bits_wen(core_io_rocc_fpu_req_bits_wen),
    .io_rocc_fpu_req_bits_ren1(core_io_rocc_fpu_req_bits_ren1),
    .io_rocc_fpu_req_bits_ren2(core_io_rocc_fpu_req_bits_ren2),
    .io_rocc_fpu_req_bits_ren3(core_io_rocc_fpu_req_bits_ren3),
    .io_rocc_fpu_req_bits_swap12(core_io_rocc_fpu_req_bits_swap12),
    .io_rocc_fpu_req_bits_swap23(core_io_rocc_fpu_req_bits_swap23),
    .io_rocc_fpu_req_bits_single(core_io_rocc_fpu_req_bits_single),
    .io_rocc_fpu_req_bits_fromint(core_io_rocc_fpu_req_bits_fromint),
    .io_rocc_fpu_req_bits_toint(core_io_rocc_fpu_req_bits_toint),
    .io_rocc_fpu_req_bits_fastpipe(core_io_rocc_fpu_req_bits_fastpipe),
    .io_rocc_fpu_req_bits_fma(core_io_rocc_fpu_req_bits_fma),
    .io_rocc_fpu_req_bits_div(core_io_rocc_fpu_req_bits_div),
    .io_rocc_fpu_req_bits_sqrt(core_io_rocc_fpu_req_bits_sqrt),
    .io_rocc_fpu_req_bits_round(core_io_rocc_fpu_req_bits_round),
    .io_rocc_fpu_req_bits_wflags(core_io_rocc_fpu_req_bits_wflags),
    .io_rocc_fpu_req_bits_rm(core_io_rocc_fpu_req_bits_rm),
    .io_rocc_fpu_req_bits_typ(core_io_rocc_fpu_req_bits_typ),
    .io_rocc_fpu_req_bits_in1(core_io_rocc_fpu_req_bits_in1),
    .io_rocc_fpu_req_bits_in2(core_io_rocc_fpu_req_bits_in2),
    .io_rocc_fpu_req_bits_in3(core_io_rocc_fpu_req_bits_in3),
    .io_rocc_fpu_resp_ready(core_io_rocc_fpu_resp_ready),
    .io_rocc_fpu_resp_valid(core_io_rocc_fpu_resp_valid),
    .io_rocc_fpu_resp_bits_data(core_io_rocc_fpu_resp_bits_data),
    .io_rocc_fpu_resp_bits_exc(core_io_rocc_fpu_resp_bits_exc),
    .io_rocc_exception(core_io_rocc_exception),
    .io_rocc_csr_waddr(core_io_rocc_csr_waddr),
    .io_rocc_csr_wdata(core_io_rocc_csr_wdata),
    .io_rocc_csr_wen(core_io_rocc_csr_wen),
    .io_rocc_host_id(core_io_rocc_host_id)
  );
  Frontend icache (
    .clk(icache_clk),
    .reset(icache_reset),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_pc(icache_io_cpu_req_bits_pc),
    .io_cpu_resp_ready(icache_io_cpu_resp_ready),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(icache_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_data_0(icache_io_cpu_resp_bits_data_0),
    .io_cpu_resp_bits_mask(icache_io_cpu_resp_bits_mask),
    .io_cpu_resp_bits_xcpt_if(icache_io_cpu_resp_bits_xcpt_if),
    .io_cpu_btb_resp_valid(icache_io_cpu_btb_resp_valid),
    .io_cpu_btb_resp_bits_taken(icache_io_cpu_btb_resp_bits_taken),
    .io_cpu_btb_resp_bits_mask(icache_io_cpu_btb_resp_bits_mask),
    .io_cpu_btb_resp_bits_bridx(icache_io_cpu_btb_resp_bits_bridx),
    .io_cpu_btb_resp_bits_target(icache_io_cpu_btb_resp_bits_target),
    .io_cpu_btb_resp_bits_entry(icache_io_cpu_btb_resp_bits_entry),
    .io_cpu_btb_resp_bits_bht_history(icache_io_cpu_btb_resp_bits_bht_history),
    .io_cpu_btb_resp_bits_bht_value(icache_io_cpu_btb_resp_bits_bht_value),
    .io_cpu_btb_update_valid(icache_io_cpu_btb_update_valid),
    .io_cpu_btb_update_bits_prediction_valid(icache_io_cpu_btb_update_bits_prediction_valid),
    .io_cpu_btb_update_bits_prediction_bits_taken(icache_io_cpu_btb_update_bits_prediction_bits_taken),
    .io_cpu_btb_update_bits_prediction_bits_mask(icache_io_cpu_btb_update_bits_prediction_bits_mask),
    .io_cpu_btb_update_bits_prediction_bits_bridx(icache_io_cpu_btb_update_bits_prediction_bits_bridx),
    .io_cpu_btb_update_bits_prediction_bits_target(icache_io_cpu_btb_update_bits_prediction_bits_target),
    .io_cpu_btb_update_bits_prediction_bits_entry(icache_io_cpu_btb_update_bits_prediction_bits_entry),
    .io_cpu_btb_update_bits_prediction_bits_bht_history(icache_io_cpu_btb_update_bits_prediction_bits_bht_history),
    .io_cpu_btb_update_bits_prediction_bits_bht_value(icache_io_cpu_btb_update_bits_prediction_bits_bht_value),
    .io_cpu_btb_update_bits_pc(icache_io_cpu_btb_update_bits_pc),
    .io_cpu_btb_update_bits_target(icache_io_cpu_btb_update_bits_target),
    .io_cpu_btb_update_bits_taken(icache_io_cpu_btb_update_bits_taken),
    .io_cpu_btb_update_bits_isJump(icache_io_cpu_btb_update_bits_isJump),
    .io_cpu_btb_update_bits_isReturn(icache_io_cpu_btb_update_bits_isReturn),
    .io_cpu_btb_update_bits_br_pc(icache_io_cpu_btb_update_bits_br_pc),
    .io_cpu_bht_update_valid(icache_io_cpu_bht_update_valid),
    .io_cpu_bht_update_bits_prediction_valid(icache_io_cpu_bht_update_bits_prediction_valid),
    .io_cpu_bht_update_bits_prediction_bits_taken(icache_io_cpu_bht_update_bits_prediction_bits_taken),
    .io_cpu_bht_update_bits_prediction_bits_mask(icache_io_cpu_bht_update_bits_prediction_bits_mask),
    .io_cpu_bht_update_bits_prediction_bits_bridx(icache_io_cpu_bht_update_bits_prediction_bits_bridx),
    .io_cpu_bht_update_bits_prediction_bits_target(icache_io_cpu_bht_update_bits_prediction_bits_target),
    .io_cpu_bht_update_bits_prediction_bits_entry(icache_io_cpu_bht_update_bits_prediction_bits_entry),
    .io_cpu_bht_update_bits_prediction_bits_bht_history(icache_io_cpu_bht_update_bits_prediction_bits_bht_history),
    .io_cpu_bht_update_bits_prediction_bits_bht_value(icache_io_cpu_bht_update_bits_prediction_bits_bht_value),
    .io_cpu_bht_update_bits_pc(icache_io_cpu_bht_update_bits_pc),
    .io_cpu_bht_update_bits_taken(icache_io_cpu_bht_update_bits_taken),
    .io_cpu_bht_update_bits_mispredict(icache_io_cpu_bht_update_bits_mispredict),
    .io_cpu_ras_update_valid(icache_io_cpu_ras_update_valid),
    .io_cpu_ras_update_bits_isCall(icache_io_cpu_ras_update_bits_isCall),
    .io_cpu_ras_update_bits_isReturn(icache_io_cpu_ras_update_bits_isReturn),
    .io_cpu_ras_update_bits_returnAddr(icache_io_cpu_ras_update_bits_returnAddr),
    .io_cpu_ras_update_bits_prediction_valid(icache_io_cpu_ras_update_bits_prediction_valid),
    .io_cpu_ras_update_bits_prediction_bits_taken(icache_io_cpu_ras_update_bits_prediction_bits_taken),
    .io_cpu_ras_update_bits_prediction_bits_mask(icache_io_cpu_ras_update_bits_prediction_bits_mask),
    .io_cpu_ras_update_bits_prediction_bits_bridx(icache_io_cpu_ras_update_bits_prediction_bits_bridx),
    .io_cpu_ras_update_bits_prediction_bits_target(icache_io_cpu_ras_update_bits_prediction_bits_target),
    .io_cpu_ras_update_bits_prediction_bits_entry(icache_io_cpu_ras_update_bits_prediction_bits_entry),
    .io_cpu_ras_update_bits_prediction_bits_bht_history(icache_io_cpu_ras_update_bits_prediction_bits_bht_history),
    .io_cpu_ras_update_bits_prediction_bits_bht_value(icache_io_cpu_ras_update_bits_prediction_bits_bht_value),
    .io_cpu_flush_icache(icache_io_cpu_flush_icache),
    .io_cpu_flush_tlb(icache_io_cpu_flush_tlb),
    .io_cpu_npc(icache_io_cpu_npc),
    .io_ptw_req_ready(icache_io_ptw_req_ready),
    .io_ptw_req_valid(icache_io_ptw_req_valid),
    .io_ptw_req_bits_addr(icache_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(icache_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(icache_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(icache_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(icache_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(icache_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(icache_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(icache_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(icache_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(icache_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(icache_io_ptw_resp_bits_pte_v),
    .io_ptw_status_debug(icache_io_ptw_status_debug),
    .io_ptw_status_prv(icache_io_ptw_status_prv),
    .io_ptw_status_sd(icache_io_ptw_status_sd),
    .io_ptw_status_zero3(icache_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(icache_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(icache_io_ptw_status_zero2),
    .io_ptw_status_vm(icache_io_ptw_status_vm),
    .io_ptw_status_zero1(icache_io_ptw_status_zero1),
    .io_ptw_status_pum(icache_io_ptw_status_pum),
    .io_ptw_status_mprv(icache_io_ptw_status_mprv),
    .io_ptw_status_xs(icache_io_ptw_status_xs),
    .io_ptw_status_fs(icache_io_ptw_status_fs),
    .io_ptw_status_mpp(icache_io_ptw_status_mpp),
    .io_ptw_status_hpp(icache_io_ptw_status_hpp),
    .io_ptw_status_spp(icache_io_ptw_status_spp),
    .io_ptw_status_mpie(icache_io_ptw_status_mpie),
    .io_ptw_status_hpie(icache_io_ptw_status_hpie),
    .io_ptw_status_spie(icache_io_ptw_status_spie),
    .io_ptw_status_upie(icache_io_ptw_status_upie),
    .io_ptw_status_mie(icache_io_ptw_status_mie),
    .io_ptw_status_hie(icache_io_ptw_status_hie),
    .io_ptw_status_sie(icache_io_ptw_status_sie),
    .io_ptw_status_uie(icache_io_ptw_status_uie),
    .io_ptw_invalidate(icache_io_ptw_invalidate),
    .io_mem_acquire_ready(icache_io_mem_acquire_ready),
    .io_mem_acquire_valid(icache_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(icache_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(icache_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(icache_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(icache_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(icache_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(icache_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(icache_io_mem_acquire_bits_data),
    .io_mem_grant_ready(icache_io_mem_grant_ready),
    .io_mem_grant_valid(icache_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(icache_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(icache_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(icache_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(icache_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(icache_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(icache_io_mem_grant_bits_data)
  );
  HellaCache HellaCache_3557 (
    .clk(HellaCache_3557_clk),
    .reset(HellaCache_3557_reset),
    .io_cpu_req_ready(HellaCache_3557_io_cpu_req_ready),
    .io_cpu_req_valid(HellaCache_3557_io_cpu_req_valid),
    .io_cpu_req_bits_addr(HellaCache_3557_io_cpu_req_bits_addr),
    .io_cpu_req_bits_tag(HellaCache_3557_io_cpu_req_bits_tag),
    .io_cpu_req_bits_cmd(HellaCache_3557_io_cpu_req_bits_cmd),
    .io_cpu_req_bits_typ(HellaCache_3557_io_cpu_req_bits_typ),
    .io_cpu_req_bits_phys(HellaCache_3557_io_cpu_req_bits_phys),
    .io_cpu_req_bits_data(HellaCache_3557_io_cpu_req_bits_data),
    .io_cpu_s1_kill(HellaCache_3557_io_cpu_s1_kill),
    .io_cpu_s1_data(HellaCache_3557_io_cpu_s1_data),
    .io_cpu_s2_nack(HellaCache_3557_io_cpu_s2_nack),
    .io_cpu_resp_valid(HellaCache_3557_io_cpu_resp_valid),
    .io_cpu_resp_bits_addr(HellaCache_3557_io_cpu_resp_bits_addr),
    .io_cpu_resp_bits_tag(HellaCache_3557_io_cpu_resp_bits_tag),
    .io_cpu_resp_bits_cmd(HellaCache_3557_io_cpu_resp_bits_cmd),
    .io_cpu_resp_bits_typ(HellaCache_3557_io_cpu_resp_bits_typ),
    .io_cpu_resp_bits_data(HellaCache_3557_io_cpu_resp_bits_data),
    .io_cpu_resp_bits_replay(HellaCache_3557_io_cpu_resp_bits_replay),
    .io_cpu_resp_bits_has_data(HellaCache_3557_io_cpu_resp_bits_has_data),
    .io_cpu_resp_bits_data_word_bypass(HellaCache_3557_io_cpu_resp_bits_data_word_bypass),
    .io_cpu_resp_bits_store_data(HellaCache_3557_io_cpu_resp_bits_store_data),
    .io_cpu_replay_next(HellaCache_3557_io_cpu_replay_next),
    .io_cpu_xcpt_ma_ld(HellaCache_3557_io_cpu_xcpt_ma_ld),
    .io_cpu_xcpt_ma_st(HellaCache_3557_io_cpu_xcpt_ma_st),
    .io_cpu_xcpt_pf_ld(HellaCache_3557_io_cpu_xcpt_pf_ld),
    .io_cpu_xcpt_pf_st(HellaCache_3557_io_cpu_xcpt_pf_st),
    .io_cpu_invalidate_lr(HellaCache_3557_io_cpu_invalidate_lr),
    .io_cpu_ordered(HellaCache_3557_io_cpu_ordered),
    .io_ptw_req_ready(HellaCache_3557_io_ptw_req_ready),
    .io_ptw_req_valid(HellaCache_3557_io_ptw_req_valid),
    .io_ptw_req_bits_addr(HellaCache_3557_io_ptw_req_bits_addr),
    .io_ptw_req_bits_prv(HellaCache_3557_io_ptw_req_bits_prv),
    .io_ptw_req_bits_store(HellaCache_3557_io_ptw_req_bits_store),
    .io_ptw_req_bits_fetch(HellaCache_3557_io_ptw_req_bits_fetch),
    .io_ptw_resp_valid(HellaCache_3557_io_ptw_resp_valid),
    .io_ptw_resp_bits_pte_ppn(HellaCache_3557_io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_reserved_for_software(HellaCache_3557_io_ptw_resp_bits_pte_reserved_for_software),
    .io_ptw_resp_bits_pte_d(HellaCache_3557_io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_r(HellaCache_3557_io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_typ(HellaCache_3557_io_ptw_resp_bits_pte_typ),
    .io_ptw_resp_bits_pte_v(HellaCache_3557_io_ptw_resp_bits_pte_v),
    .io_ptw_status_debug(HellaCache_3557_io_ptw_status_debug),
    .io_ptw_status_prv(HellaCache_3557_io_ptw_status_prv),
    .io_ptw_status_sd(HellaCache_3557_io_ptw_status_sd),
    .io_ptw_status_zero3(HellaCache_3557_io_ptw_status_zero3),
    .io_ptw_status_sd_rv32(HellaCache_3557_io_ptw_status_sd_rv32),
    .io_ptw_status_zero2(HellaCache_3557_io_ptw_status_zero2),
    .io_ptw_status_vm(HellaCache_3557_io_ptw_status_vm),
    .io_ptw_status_zero1(HellaCache_3557_io_ptw_status_zero1),
    .io_ptw_status_pum(HellaCache_3557_io_ptw_status_pum),
    .io_ptw_status_mprv(HellaCache_3557_io_ptw_status_mprv),
    .io_ptw_status_xs(HellaCache_3557_io_ptw_status_xs),
    .io_ptw_status_fs(HellaCache_3557_io_ptw_status_fs),
    .io_ptw_status_mpp(HellaCache_3557_io_ptw_status_mpp),
    .io_ptw_status_hpp(HellaCache_3557_io_ptw_status_hpp),
    .io_ptw_status_spp(HellaCache_3557_io_ptw_status_spp),
    .io_ptw_status_mpie(HellaCache_3557_io_ptw_status_mpie),
    .io_ptw_status_hpie(HellaCache_3557_io_ptw_status_hpie),
    .io_ptw_status_spie(HellaCache_3557_io_ptw_status_spie),
    .io_ptw_status_upie(HellaCache_3557_io_ptw_status_upie),
    .io_ptw_status_mie(HellaCache_3557_io_ptw_status_mie),
    .io_ptw_status_hie(HellaCache_3557_io_ptw_status_hie),
    .io_ptw_status_sie(HellaCache_3557_io_ptw_status_sie),
    .io_ptw_status_uie(HellaCache_3557_io_ptw_status_uie),
    .io_ptw_invalidate(HellaCache_3557_io_ptw_invalidate),
    .io_mem_acquire_ready(HellaCache_3557_io_mem_acquire_ready),
    .io_mem_acquire_valid(HellaCache_3557_io_mem_acquire_valid),
    .io_mem_acquire_bits_addr_block(HellaCache_3557_io_mem_acquire_bits_addr_block),
    .io_mem_acquire_bits_client_xact_id(HellaCache_3557_io_mem_acquire_bits_client_xact_id),
    .io_mem_acquire_bits_addr_beat(HellaCache_3557_io_mem_acquire_bits_addr_beat),
    .io_mem_acquire_bits_is_builtin_type(HellaCache_3557_io_mem_acquire_bits_is_builtin_type),
    .io_mem_acquire_bits_a_type(HellaCache_3557_io_mem_acquire_bits_a_type),
    .io_mem_acquire_bits_union(HellaCache_3557_io_mem_acquire_bits_union),
    .io_mem_acquire_bits_data(HellaCache_3557_io_mem_acquire_bits_data),
    .io_mem_probe_ready(HellaCache_3557_io_mem_probe_ready),
    .io_mem_probe_valid(HellaCache_3557_io_mem_probe_valid),
    .io_mem_probe_bits_addr_block(HellaCache_3557_io_mem_probe_bits_addr_block),
    .io_mem_probe_bits_p_type(HellaCache_3557_io_mem_probe_bits_p_type),
    .io_mem_release_ready(HellaCache_3557_io_mem_release_ready),
    .io_mem_release_valid(HellaCache_3557_io_mem_release_valid),
    .io_mem_release_bits_addr_beat(HellaCache_3557_io_mem_release_bits_addr_beat),
    .io_mem_release_bits_addr_block(HellaCache_3557_io_mem_release_bits_addr_block),
    .io_mem_release_bits_client_xact_id(HellaCache_3557_io_mem_release_bits_client_xact_id),
    .io_mem_release_bits_voluntary(HellaCache_3557_io_mem_release_bits_voluntary),
    .io_mem_release_bits_r_type(HellaCache_3557_io_mem_release_bits_r_type),
    .io_mem_release_bits_data(HellaCache_3557_io_mem_release_bits_data),
    .io_mem_grant_ready(HellaCache_3557_io_mem_grant_ready),
    .io_mem_grant_valid(HellaCache_3557_io_mem_grant_valid),
    .io_mem_grant_bits_addr_beat(HellaCache_3557_io_mem_grant_bits_addr_beat),
    .io_mem_grant_bits_client_xact_id(HellaCache_3557_io_mem_grant_bits_client_xact_id),
    .io_mem_grant_bits_manager_xact_id(HellaCache_3557_io_mem_grant_bits_manager_xact_id),
    .io_mem_grant_bits_is_builtin_type(HellaCache_3557_io_mem_grant_bits_is_builtin_type),
    .io_mem_grant_bits_g_type(HellaCache_3557_io_mem_grant_bits_g_type),
    .io_mem_grant_bits_data(HellaCache_3557_io_mem_grant_bits_data),
    .io_mem_grant_bits_manager_id(HellaCache_3557_io_mem_grant_bits_manager_id),
    .io_mem_finish_ready(HellaCache_3557_io_mem_finish_ready),
    .io_mem_finish_valid(HellaCache_3557_io_mem_finish_valid),
    .io_mem_finish_bits_manager_xact_id(HellaCache_3557_io_mem_finish_bits_manager_xact_id),
    .io_mem_finish_bits_manager_id(HellaCache_3557_io_mem_finish_bits_manager_id)
  );
  FPU FPU_3558 (
    .clk(FPU_3558_clk),
    .reset(FPU_3558_reset),
    .io_inst(FPU_3558_io_inst),
    .io_fromint_data(FPU_3558_io_fromint_data),
    .io_fcsr_rm(FPU_3558_io_fcsr_rm),
    .io_fcsr_flags_valid(FPU_3558_io_fcsr_flags_valid),
    .io_fcsr_flags_bits(FPU_3558_io_fcsr_flags_bits),
    .io_store_data(FPU_3558_io_store_data),
    .io_toint_data(FPU_3558_io_toint_data),
    .io_dmem_resp_val(FPU_3558_io_dmem_resp_val),
    .io_dmem_resp_type(FPU_3558_io_dmem_resp_type),
    .io_dmem_resp_tag(FPU_3558_io_dmem_resp_tag),
    .io_dmem_resp_data(FPU_3558_io_dmem_resp_data),
    .io_valid(FPU_3558_io_valid),
    .io_fcsr_rdy(FPU_3558_io_fcsr_rdy),
    .io_nack_mem(FPU_3558_io_nack_mem),
    .io_illegal_rm(FPU_3558_io_illegal_rm),
    .io_killx(FPU_3558_io_killx),
    .io_killm(FPU_3558_io_killm),
    .io_dec_cmd(FPU_3558_io_dec_cmd),
    .io_dec_ldst(FPU_3558_io_dec_ldst),
    .io_dec_wen(FPU_3558_io_dec_wen),
    .io_dec_ren1(FPU_3558_io_dec_ren1),
    .io_dec_ren2(FPU_3558_io_dec_ren2),
    .io_dec_ren3(FPU_3558_io_dec_ren3),
    .io_dec_swap12(FPU_3558_io_dec_swap12),
    .io_dec_swap23(FPU_3558_io_dec_swap23),
    .io_dec_single(FPU_3558_io_dec_single),
    .io_dec_fromint(FPU_3558_io_dec_fromint),
    .io_dec_toint(FPU_3558_io_dec_toint),
    .io_dec_fastpipe(FPU_3558_io_dec_fastpipe),
    .io_dec_fma(FPU_3558_io_dec_fma),
    .io_dec_div(FPU_3558_io_dec_div),
    .io_dec_sqrt(FPU_3558_io_dec_sqrt),
    .io_dec_round(FPU_3558_io_dec_round),
    .io_dec_wflags(FPU_3558_io_dec_wflags),
    .io_sboard_set(FPU_3558_io_sboard_set),
    .io_sboard_clr(FPU_3558_io_sboard_clr),
    .io_sboard_clra(FPU_3558_io_sboard_clra),
    .io_cp_req_ready(FPU_3558_io_cp_req_ready),
    .io_cp_req_valid(FPU_3558_io_cp_req_valid),
    .io_cp_req_bits_cmd(FPU_3558_io_cp_req_bits_cmd),
    .io_cp_req_bits_ldst(FPU_3558_io_cp_req_bits_ldst),
    .io_cp_req_bits_wen(FPU_3558_io_cp_req_bits_wen),
    .io_cp_req_bits_ren1(FPU_3558_io_cp_req_bits_ren1),
    .io_cp_req_bits_ren2(FPU_3558_io_cp_req_bits_ren2),
    .io_cp_req_bits_ren3(FPU_3558_io_cp_req_bits_ren3),
    .io_cp_req_bits_swap12(FPU_3558_io_cp_req_bits_swap12),
    .io_cp_req_bits_swap23(FPU_3558_io_cp_req_bits_swap23),
    .io_cp_req_bits_single(FPU_3558_io_cp_req_bits_single),
    .io_cp_req_bits_fromint(FPU_3558_io_cp_req_bits_fromint),
    .io_cp_req_bits_toint(FPU_3558_io_cp_req_bits_toint),
    .io_cp_req_bits_fastpipe(FPU_3558_io_cp_req_bits_fastpipe),
    .io_cp_req_bits_fma(FPU_3558_io_cp_req_bits_fma),
    .io_cp_req_bits_div(FPU_3558_io_cp_req_bits_div),
    .io_cp_req_bits_sqrt(FPU_3558_io_cp_req_bits_sqrt),
    .io_cp_req_bits_round(FPU_3558_io_cp_req_bits_round),
    .io_cp_req_bits_wflags(FPU_3558_io_cp_req_bits_wflags),
    .io_cp_req_bits_rm(FPU_3558_io_cp_req_bits_rm),
    .io_cp_req_bits_typ(FPU_3558_io_cp_req_bits_typ),
    .io_cp_req_bits_in1(FPU_3558_io_cp_req_bits_in1),
    .io_cp_req_bits_in2(FPU_3558_io_cp_req_bits_in2),
    .io_cp_req_bits_in3(FPU_3558_io_cp_req_bits_in3),
    .io_cp_resp_ready(FPU_3558_io_cp_resp_ready),
    .io_cp_resp_valid(FPU_3558_io_cp_resp_valid),
    .io_cp_resp_bits_data(FPU_3558_io_cp_resp_bits_data),
    .io_cp_resp_bits_exc(FPU_3558_io_cp_resp_bits_exc)
  );
  ClientUncachedTileLinkIOArbiter_101 uncachedArb (
    .clk(uncachedArb_clk),
    .reset(uncachedArb_reset),
    .io_in_0_acquire_ready(uncachedArb_io_in_0_acquire_ready),
    .io_in_0_acquire_valid(uncachedArb_io_in_0_acquire_valid),
    .io_in_0_acquire_bits_addr_block(uncachedArb_io_in_0_acquire_bits_addr_block),
    .io_in_0_acquire_bits_client_xact_id(uncachedArb_io_in_0_acquire_bits_client_xact_id),
    .io_in_0_acquire_bits_addr_beat(uncachedArb_io_in_0_acquire_bits_addr_beat),
    .io_in_0_acquire_bits_is_builtin_type(uncachedArb_io_in_0_acquire_bits_is_builtin_type),
    .io_in_0_acquire_bits_a_type(uncachedArb_io_in_0_acquire_bits_a_type),
    .io_in_0_acquire_bits_union(uncachedArb_io_in_0_acquire_bits_union),
    .io_in_0_acquire_bits_data(uncachedArb_io_in_0_acquire_bits_data),
    .io_in_0_grant_ready(uncachedArb_io_in_0_grant_ready),
    .io_in_0_grant_valid(uncachedArb_io_in_0_grant_valid),
    .io_in_0_grant_bits_addr_beat(uncachedArb_io_in_0_grant_bits_addr_beat),
    .io_in_0_grant_bits_client_xact_id(uncachedArb_io_in_0_grant_bits_client_xact_id),
    .io_in_0_grant_bits_manager_xact_id(uncachedArb_io_in_0_grant_bits_manager_xact_id),
    .io_in_0_grant_bits_is_builtin_type(uncachedArb_io_in_0_grant_bits_is_builtin_type),
    .io_in_0_grant_bits_g_type(uncachedArb_io_in_0_grant_bits_g_type),
    .io_in_0_grant_bits_data(uncachedArb_io_in_0_grant_bits_data),
    .io_out_acquire_ready(uncachedArb_io_out_acquire_ready),
    .io_out_acquire_valid(uncachedArb_io_out_acquire_valid),
    .io_out_acquire_bits_addr_block(uncachedArb_io_out_acquire_bits_addr_block),
    .io_out_acquire_bits_client_xact_id(uncachedArb_io_out_acquire_bits_client_xact_id),
    .io_out_acquire_bits_addr_beat(uncachedArb_io_out_acquire_bits_addr_beat),
    .io_out_acquire_bits_is_builtin_type(uncachedArb_io_out_acquire_bits_is_builtin_type),
    .io_out_acquire_bits_a_type(uncachedArb_io_out_acquire_bits_a_type),
    .io_out_acquire_bits_union(uncachedArb_io_out_acquire_bits_union),
    .io_out_acquire_bits_data(uncachedArb_io_out_acquire_bits_data),
    .io_out_grant_ready(uncachedArb_io_out_grant_ready),
    .io_out_grant_valid(uncachedArb_io_out_grant_valid),
    .io_out_grant_bits_addr_beat(uncachedArb_io_out_grant_bits_addr_beat),
    .io_out_grant_bits_client_xact_id(uncachedArb_io_out_grant_bits_client_xact_id),
    .io_out_grant_bits_manager_xact_id(uncachedArb_io_out_grant_bits_manager_xact_id),
    .io_out_grant_bits_is_builtin_type(uncachedArb_io_out_grant_bits_is_builtin_type),
    .io_out_grant_bits_g_type(uncachedArb_io_out_grant_bits_g_type),
    .io_out_grant_bits_data(uncachedArb_io_out_grant_bits_data)
  );
  PTW PTW_3559 (
    .clk(PTW_3559_clk),
    .reset(PTW_3559_reset),
    .io_requestor_0_req_ready(PTW_3559_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(PTW_3559_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(PTW_3559_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_prv(PTW_3559_io_requestor_0_req_bits_prv),
    .io_requestor_0_req_bits_store(PTW_3559_io_requestor_0_req_bits_store),
    .io_requestor_0_req_bits_fetch(PTW_3559_io_requestor_0_req_bits_fetch),
    .io_requestor_0_resp_valid(PTW_3559_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_pte_ppn(PTW_3559_io_requestor_0_resp_bits_pte_ppn),
    .io_requestor_0_resp_bits_pte_reserved_for_software(PTW_3559_io_requestor_0_resp_bits_pte_reserved_for_software),
    .io_requestor_0_resp_bits_pte_d(PTW_3559_io_requestor_0_resp_bits_pte_d),
    .io_requestor_0_resp_bits_pte_r(PTW_3559_io_requestor_0_resp_bits_pte_r),
    .io_requestor_0_resp_bits_pte_typ(PTW_3559_io_requestor_0_resp_bits_pte_typ),
    .io_requestor_0_resp_bits_pte_v(PTW_3559_io_requestor_0_resp_bits_pte_v),
    .io_requestor_0_status_debug(PTW_3559_io_requestor_0_status_debug),
    .io_requestor_0_status_prv(PTW_3559_io_requestor_0_status_prv),
    .io_requestor_0_status_sd(PTW_3559_io_requestor_0_status_sd),
    .io_requestor_0_status_zero3(PTW_3559_io_requestor_0_status_zero3),
    .io_requestor_0_status_sd_rv32(PTW_3559_io_requestor_0_status_sd_rv32),
    .io_requestor_0_status_zero2(PTW_3559_io_requestor_0_status_zero2),
    .io_requestor_0_status_vm(PTW_3559_io_requestor_0_status_vm),
    .io_requestor_0_status_zero1(PTW_3559_io_requestor_0_status_zero1),
    .io_requestor_0_status_pum(PTW_3559_io_requestor_0_status_pum),
    .io_requestor_0_status_mprv(PTW_3559_io_requestor_0_status_mprv),
    .io_requestor_0_status_xs(PTW_3559_io_requestor_0_status_xs),
    .io_requestor_0_status_fs(PTW_3559_io_requestor_0_status_fs),
    .io_requestor_0_status_mpp(PTW_3559_io_requestor_0_status_mpp),
    .io_requestor_0_status_hpp(PTW_3559_io_requestor_0_status_hpp),
    .io_requestor_0_status_spp(PTW_3559_io_requestor_0_status_spp),
    .io_requestor_0_status_mpie(PTW_3559_io_requestor_0_status_mpie),
    .io_requestor_0_status_hpie(PTW_3559_io_requestor_0_status_hpie),
    .io_requestor_0_status_spie(PTW_3559_io_requestor_0_status_spie),
    .io_requestor_0_status_upie(PTW_3559_io_requestor_0_status_upie),
    .io_requestor_0_status_mie(PTW_3559_io_requestor_0_status_mie),
    .io_requestor_0_status_hie(PTW_3559_io_requestor_0_status_hie),
    .io_requestor_0_status_sie(PTW_3559_io_requestor_0_status_sie),
    .io_requestor_0_status_uie(PTW_3559_io_requestor_0_status_uie),
    .io_requestor_0_invalidate(PTW_3559_io_requestor_0_invalidate),
    .io_requestor_1_req_ready(PTW_3559_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(PTW_3559_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(PTW_3559_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_prv(PTW_3559_io_requestor_1_req_bits_prv),
    .io_requestor_1_req_bits_store(PTW_3559_io_requestor_1_req_bits_store),
    .io_requestor_1_req_bits_fetch(PTW_3559_io_requestor_1_req_bits_fetch),
    .io_requestor_1_resp_valid(PTW_3559_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_pte_ppn(PTW_3559_io_requestor_1_resp_bits_pte_ppn),
    .io_requestor_1_resp_bits_pte_reserved_for_software(PTW_3559_io_requestor_1_resp_bits_pte_reserved_for_software),
    .io_requestor_1_resp_bits_pte_d(PTW_3559_io_requestor_1_resp_bits_pte_d),
    .io_requestor_1_resp_bits_pte_r(PTW_3559_io_requestor_1_resp_bits_pte_r),
    .io_requestor_1_resp_bits_pte_typ(PTW_3559_io_requestor_1_resp_bits_pte_typ),
    .io_requestor_1_resp_bits_pte_v(PTW_3559_io_requestor_1_resp_bits_pte_v),
    .io_requestor_1_status_debug(PTW_3559_io_requestor_1_status_debug),
    .io_requestor_1_status_prv(PTW_3559_io_requestor_1_status_prv),
    .io_requestor_1_status_sd(PTW_3559_io_requestor_1_status_sd),
    .io_requestor_1_status_zero3(PTW_3559_io_requestor_1_status_zero3),
    .io_requestor_1_status_sd_rv32(PTW_3559_io_requestor_1_status_sd_rv32),
    .io_requestor_1_status_zero2(PTW_3559_io_requestor_1_status_zero2),
    .io_requestor_1_status_vm(PTW_3559_io_requestor_1_status_vm),
    .io_requestor_1_status_zero1(PTW_3559_io_requestor_1_status_zero1),
    .io_requestor_1_status_pum(PTW_3559_io_requestor_1_status_pum),
    .io_requestor_1_status_mprv(PTW_3559_io_requestor_1_status_mprv),
    .io_requestor_1_status_xs(PTW_3559_io_requestor_1_status_xs),
    .io_requestor_1_status_fs(PTW_3559_io_requestor_1_status_fs),
    .io_requestor_1_status_mpp(PTW_3559_io_requestor_1_status_mpp),
    .io_requestor_1_status_hpp(PTW_3559_io_requestor_1_status_hpp),
    .io_requestor_1_status_spp(PTW_3559_io_requestor_1_status_spp),
    .io_requestor_1_status_mpie(PTW_3559_io_requestor_1_status_mpie),
    .io_requestor_1_status_hpie(PTW_3559_io_requestor_1_status_hpie),
    .io_requestor_1_status_spie(PTW_3559_io_requestor_1_status_spie),
    .io_requestor_1_status_upie(PTW_3559_io_requestor_1_status_upie),
    .io_requestor_1_status_mie(PTW_3559_io_requestor_1_status_mie),
    .io_requestor_1_status_hie(PTW_3559_io_requestor_1_status_hie),
    .io_requestor_1_status_sie(PTW_3559_io_requestor_1_status_sie),
    .io_requestor_1_status_uie(PTW_3559_io_requestor_1_status_uie),
    .io_requestor_1_invalidate(PTW_3559_io_requestor_1_invalidate),
    .io_mem_req_ready(PTW_3559_io_mem_req_ready),
    .io_mem_req_valid(PTW_3559_io_mem_req_valid),
    .io_mem_req_bits_addr(PTW_3559_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(PTW_3559_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(PTW_3559_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(PTW_3559_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(PTW_3559_io_mem_req_bits_phys),
    .io_mem_req_bits_data(PTW_3559_io_mem_req_bits_data),
    .io_mem_s1_kill(PTW_3559_io_mem_s1_kill),
    .io_mem_s1_data(PTW_3559_io_mem_s1_data),
    .io_mem_s2_nack(PTW_3559_io_mem_s2_nack),
    .io_mem_resp_valid(PTW_3559_io_mem_resp_valid),
    .io_mem_resp_bits_addr(PTW_3559_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(PTW_3559_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(PTW_3559_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(PTW_3559_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(PTW_3559_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(PTW_3559_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(PTW_3559_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(PTW_3559_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(PTW_3559_io_mem_resp_bits_store_data),
    .io_mem_replay_next(PTW_3559_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(PTW_3559_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(PTW_3559_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(PTW_3559_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(PTW_3559_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(PTW_3559_io_mem_invalidate_lr),
    .io_mem_ordered(PTW_3559_io_mem_ordered),
    .io_dpath_ptbr(PTW_3559_io_dpath_ptbr),
    .io_dpath_invalidate(PTW_3559_io_dpath_invalidate),
    .io_dpath_status_debug(PTW_3559_io_dpath_status_debug),
    .io_dpath_status_prv(PTW_3559_io_dpath_status_prv),
    .io_dpath_status_sd(PTW_3559_io_dpath_status_sd),
    .io_dpath_status_zero3(PTW_3559_io_dpath_status_zero3),
    .io_dpath_status_sd_rv32(PTW_3559_io_dpath_status_sd_rv32),
    .io_dpath_status_zero2(PTW_3559_io_dpath_status_zero2),
    .io_dpath_status_vm(PTW_3559_io_dpath_status_vm),
    .io_dpath_status_zero1(PTW_3559_io_dpath_status_zero1),
    .io_dpath_status_pum(PTW_3559_io_dpath_status_pum),
    .io_dpath_status_mprv(PTW_3559_io_dpath_status_mprv),
    .io_dpath_status_xs(PTW_3559_io_dpath_status_xs),
    .io_dpath_status_fs(PTW_3559_io_dpath_status_fs),
    .io_dpath_status_mpp(PTW_3559_io_dpath_status_mpp),
    .io_dpath_status_hpp(PTW_3559_io_dpath_status_hpp),
    .io_dpath_status_spp(PTW_3559_io_dpath_status_spp),
    .io_dpath_status_mpie(PTW_3559_io_dpath_status_mpie),
    .io_dpath_status_hpie(PTW_3559_io_dpath_status_hpie),
    .io_dpath_status_spie(PTW_3559_io_dpath_status_spie),
    .io_dpath_status_upie(PTW_3559_io_dpath_status_upie),
    .io_dpath_status_mie(PTW_3559_io_dpath_status_mie),
    .io_dpath_status_hie(PTW_3559_io_dpath_status_hie),
    .io_dpath_status_sie(PTW_3559_io_dpath_status_sie),
    .io_dpath_status_uie(PTW_3559_io_dpath_status_uie)
  );
  HellaCacheArbiter dcArb (
    .clk(dcArb_clk),
    .reset(dcArb_reset),
    .io_requestor_0_req_ready(dcArb_io_requestor_0_req_ready),
    .io_requestor_0_req_valid(dcArb_io_requestor_0_req_valid),
    .io_requestor_0_req_bits_addr(dcArb_io_requestor_0_req_bits_addr),
    .io_requestor_0_req_bits_tag(dcArb_io_requestor_0_req_bits_tag),
    .io_requestor_0_req_bits_cmd(dcArb_io_requestor_0_req_bits_cmd),
    .io_requestor_0_req_bits_typ(dcArb_io_requestor_0_req_bits_typ),
    .io_requestor_0_req_bits_phys(dcArb_io_requestor_0_req_bits_phys),
    .io_requestor_0_req_bits_data(dcArb_io_requestor_0_req_bits_data),
    .io_requestor_0_s1_kill(dcArb_io_requestor_0_s1_kill),
    .io_requestor_0_s1_data(dcArb_io_requestor_0_s1_data),
    .io_requestor_0_s2_nack(dcArb_io_requestor_0_s2_nack),
    .io_requestor_0_resp_valid(dcArb_io_requestor_0_resp_valid),
    .io_requestor_0_resp_bits_addr(dcArb_io_requestor_0_resp_bits_addr),
    .io_requestor_0_resp_bits_tag(dcArb_io_requestor_0_resp_bits_tag),
    .io_requestor_0_resp_bits_cmd(dcArb_io_requestor_0_resp_bits_cmd),
    .io_requestor_0_resp_bits_typ(dcArb_io_requestor_0_resp_bits_typ),
    .io_requestor_0_resp_bits_data(dcArb_io_requestor_0_resp_bits_data),
    .io_requestor_0_resp_bits_replay(dcArb_io_requestor_0_resp_bits_replay),
    .io_requestor_0_resp_bits_has_data(dcArb_io_requestor_0_resp_bits_has_data),
    .io_requestor_0_resp_bits_data_word_bypass(dcArb_io_requestor_0_resp_bits_data_word_bypass),
    .io_requestor_0_resp_bits_store_data(dcArb_io_requestor_0_resp_bits_store_data),
    .io_requestor_0_replay_next(dcArb_io_requestor_0_replay_next),
    .io_requestor_0_xcpt_ma_ld(dcArb_io_requestor_0_xcpt_ma_ld),
    .io_requestor_0_xcpt_ma_st(dcArb_io_requestor_0_xcpt_ma_st),
    .io_requestor_0_xcpt_pf_ld(dcArb_io_requestor_0_xcpt_pf_ld),
    .io_requestor_0_xcpt_pf_st(dcArb_io_requestor_0_xcpt_pf_st),
    .io_requestor_0_invalidate_lr(dcArb_io_requestor_0_invalidate_lr),
    .io_requestor_0_ordered(dcArb_io_requestor_0_ordered),
    .io_requestor_1_req_ready(dcArb_io_requestor_1_req_ready),
    .io_requestor_1_req_valid(dcArb_io_requestor_1_req_valid),
    .io_requestor_1_req_bits_addr(dcArb_io_requestor_1_req_bits_addr),
    .io_requestor_1_req_bits_tag(dcArb_io_requestor_1_req_bits_tag),
    .io_requestor_1_req_bits_cmd(dcArb_io_requestor_1_req_bits_cmd),
    .io_requestor_1_req_bits_typ(dcArb_io_requestor_1_req_bits_typ),
    .io_requestor_1_req_bits_phys(dcArb_io_requestor_1_req_bits_phys),
    .io_requestor_1_req_bits_data(dcArb_io_requestor_1_req_bits_data),
    .io_requestor_1_s1_kill(dcArb_io_requestor_1_s1_kill),
    .io_requestor_1_s1_data(dcArb_io_requestor_1_s1_data),
    .io_requestor_1_s2_nack(dcArb_io_requestor_1_s2_nack),
    .io_requestor_1_resp_valid(dcArb_io_requestor_1_resp_valid),
    .io_requestor_1_resp_bits_addr(dcArb_io_requestor_1_resp_bits_addr),
    .io_requestor_1_resp_bits_tag(dcArb_io_requestor_1_resp_bits_tag),
    .io_requestor_1_resp_bits_cmd(dcArb_io_requestor_1_resp_bits_cmd),
    .io_requestor_1_resp_bits_typ(dcArb_io_requestor_1_resp_bits_typ),
    .io_requestor_1_resp_bits_data(dcArb_io_requestor_1_resp_bits_data),
    .io_requestor_1_resp_bits_replay(dcArb_io_requestor_1_resp_bits_replay),
    .io_requestor_1_resp_bits_has_data(dcArb_io_requestor_1_resp_bits_has_data),
    .io_requestor_1_resp_bits_data_word_bypass(dcArb_io_requestor_1_resp_bits_data_word_bypass),
    .io_requestor_1_resp_bits_store_data(dcArb_io_requestor_1_resp_bits_store_data),
    .io_requestor_1_replay_next(dcArb_io_requestor_1_replay_next),
    .io_requestor_1_xcpt_ma_ld(dcArb_io_requestor_1_xcpt_ma_ld),
    .io_requestor_1_xcpt_ma_st(dcArb_io_requestor_1_xcpt_ma_st),
    .io_requestor_1_xcpt_pf_ld(dcArb_io_requestor_1_xcpt_pf_ld),
    .io_requestor_1_xcpt_pf_st(dcArb_io_requestor_1_xcpt_pf_st),
    .io_requestor_1_invalidate_lr(dcArb_io_requestor_1_invalidate_lr),
    .io_requestor_1_ordered(dcArb_io_requestor_1_ordered),
    .io_mem_req_ready(dcArb_io_mem_req_ready),
    .io_mem_req_valid(dcArb_io_mem_req_valid),
    .io_mem_req_bits_addr(dcArb_io_mem_req_bits_addr),
    .io_mem_req_bits_tag(dcArb_io_mem_req_bits_tag),
    .io_mem_req_bits_cmd(dcArb_io_mem_req_bits_cmd),
    .io_mem_req_bits_typ(dcArb_io_mem_req_bits_typ),
    .io_mem_req_bits_phys(dcArb_io_mem_req_bits_phys),
    .io_mem_req_bits_data(dcArb_io_mem_req_bits_data),
    .io_mem_s1_kill(dcArb_io_mem_s1_kill),
    .io_mem_s1_data(dcArb_io_mem_s1_data),
    .io_mem_s2_nack(dcArb_io_mem_s2_nack),
    .io_mem_resp_valid(dcArb_io_mem_resp_valid),
    .io_mem_resp_bits_addr(dcArb_io_mem_resp_bits_addr),
    .io_mem_resp_bits_tag(dcArb_io_mem_resp_bits_tag),
    .io_mem_resp_bits_cmd(dcArb_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_typ(dcArb_io_mem_resp_bits_typ),
    .io_mem_resp_bits_data(dcArb_io_mem_resp_bits_data),
    .io_mem_resp_bits_replay(dcArb_io_mem_resp_bits_replay),
    .io_mem_resp_bits_has_data(dcArb_io_mem_resp_bits_has_data),
    .io_mem_resp_bits_data_word_bypass(dcArb_io_mem_resp_bits_data_word_bypass),
    .io_mem_resp_bits_store_data(dcArb_io_mem_resp_bits_store_data),
    .io_mem_replay_next(dcArb_io_mem_replay_next),
    .io_mem_xcpt_ma_ld(dcArb_io_mem_xcpt_ma_ld),
    .io_mem_xcpt_ma_st(dcArb_io_mem_xcpt_ma_st),
    .io_mem_xcpt_pf_ld(dcArb_io_mem_xcpt_pf_ld),
    .io_mem_xcpt_pf_st(dcArb_io_mem_xcpt_pf_st),
    .io_mem_invalidate_lr(dcArb_io_mem_invalidate_lr),
    .io_mem_ordered(dcArb_io_mem_ordered)
  );
  assign io_cached_0_acquire_valid = HellaCache_3557_io_mem_acquire_valid;
  assign io_cached_0_acquire_bits_addr_block = HellaCache_3557_io_mem_acquire_bits_addr_block;
  assign io_cached_0_acquire_bits_client_xact_id = HellaCache_3557_io_mem_acquire_bits_client_xact_id;
  assign io_cached_0_acquire_bits_addr_beat = HellaCache_3557_io_mem_acquire_bits_addr_beat;
  assign io_cached_0_acquire_bits_is_builtin_type = HellaCache_3557_io_mem_acquire_bits_is_builtin_type;
  assign io_cached_0_acquire_bits_a_type = HellaCache_3557_io_mem_acquire_bits_a_type;
  assign io_cached_0_acquire_bits_union = HellaCache_3557_io_mem_acquire_bits_union;
  assign io_cached_0_acquire_bits_data = HellaCache_3557_io_mem_acquire_bits_data;
  assign io_cached_0_probe_ready = HellaCache_3557_io_mem_probe_ready;
  assign io_cached_0_release_valid = HellaCache_3557_io_mem_release_valid;
  assign io_cached_0_release_bits_addr_beat = HellaCache_3557_io_mem_release_bits_addr_beat;
  assign io_cached_0_release_bits_addr_block = HellaCache_3557_io_mem_release_bits_addr_block;
  assign io_cached_0_release_bits_client_xact_id = HellaCache_3557_io_mem_release_bits_client_xact_id;
  assign io_cached_0_release_bits_voluntary = HellaCache_3557_io_mem_release_bits_voluntary;
  assign io_cached_0_release_bits_r_type = HellaCache_3557_io_mem_release_bits_r_type;
  assign io_cached_0_release_bits_data = HellaCache_3557_io_mem_release_bits_data;
  assign io_cached_0_grant_ready = HellaCache_3557_io_mem_grant_ready;
  assign io_cached_0_finish_valid = HellaCache_3557_io_mem_finish_valid;
  assign io_cached_0_finish_bits_manager_xact_id = HellaCache_3557_io_mem_finish_bits_manager_xact_id;
  assign io_cached_0_finish_bits_manager_id = HellaCache_3557_io_mem_finish_bits_manager_id;
  assign io_uncached_0_acquire_valid = uncachedArb_io_out_acquire_valid;
  assign io_uncached_0_acquire_bits_addr_block = uncachedArb_io_out_acquire_bits_addr_block;
  assign io_uncached_0_acquire_bits_client_xact_id = uncachedArb_io_out_acquire_bits_client_xact_id;
  assign io_uncached_0_acquire_bits_addr_beat = uncachedArb_io_out_acquire_bits_addr_beat;
  assign io_uncached_0_acquire_bits_is_builtin_type = uncachedArb_io_out_acquire_bits_is_builtin_type;
  assign io_uncached_0_acquire_bits_a_type = uncachedArb_io_out_acquire_bits_a_type;
  assign io_uncached_0_acquire_bits_union = uncachedArb_io_out_acquire_bits_union;
  assign io_uncached_0_acquire_bits_data = uncachedArb_io_out_acquire_bits_data;
  assign io_uncached_0_grant_ready = uncachedArb_io_out_grant_ready;
  assign io_dma_req_valid = GEN_0;
  assign io_dma_req_bits_xact_id = GEN_1;
  assign io_dma_req_bits_client_id = GEN_2;
  assign io_dma_req_bits_cmd = GEN_3;
  assign io_dma_req_bits_source = GEN_4;
  assign io_dma_req_bits_dest = GEN_5;
  assign io_dma_req_bits_length = GEN_6;
  assign io_dma_req_bits_size = GEN_7;
  assign io_dma_resp_ready = GEN_8;
  assign core_clk = clk;
  assign core_reset = reset;
  assign core_io_prci_reset = io_prci_reset;
  assign core_io_prci_id = io_prci_id;
  assign core_io_prci_interrupts_mtip = io_prci_interrupts_mtip;
  assign core_io_prci_interrupts_meip = io_prci_interrupts_meip;
  assign core_io_prci_interrupts_seip = io_prci_interrupts_seip;
  assign core_io_prci_interrupts_debug = io_prci_interrupts_debug;
  assign core_io_prci_interrupts_msip = io_prci_interrupts_msip;
  assign core_io_imem_resp_valid = icache_io_cpu_resp_valid;
  assign core_io_imem_resp_bits_pc = icache_io_cpu_resp_bits_pc;
  assign core_io_imem_resp_bits_data_0 = icache_io_cpu_resp_bits_data_0;
  assign core_io_imem_resp_bits_mask = icache_io_cpu_resp_bits_mask;
  assign core_io_imem_resp_bits_xcpt_if = icache_io_cpu_resp_bits_xcpt_if;
  assign core_io_imem_btb_resp_valid = icache_io_cpu_btb_resp_valid;
  assign core_io_imem_btb_resp_bits_taken = icache_io_cpu_btb_resp_bits_taken;
  assign core_io_imem_btb_resp_bits_mask = icache_io_cpu_btb_resp_bits_mask;
  assign core_io_imem_btb_resp_bits_bridx = icache_io_cpu_btb_resp_bits_bridx;
  assign core_io_imem_btb_resp_bits_target = icache_io_cpu_btb_resp_bits_target;
  assign core_io_imem_btb_resp_bits_entry = icache_io_cpu_btb_resp_bits_entry;
  assign core_io_imem_btb_resp_bits_bht_history = icache_io_cpu_btb_resp_bits_bht_history;
  assign core_io_imem_btb_resp_bits_bht_value = icache_io_cpu_btb_resp_bits_bht_value;
  assign core_io_imem_npc = icache_io_cpu_npc;
  assign core_io_dmem_req_ready = dcArb_io_requestor_1_req_ready;
  assign core_io_dmem_s2_nack = dcArb_io_requestor_1_s2_nack;
  assign core_io_dmem_resp_valid = dcArb_io_requestor_1_resp_valid;
  assign core_io_dmem_resp_bits_addr = dcArb_io_requestor_1_resp_bits_addr;
  assign core_io_dmem_resp_bits_tag = dcArb_io_requestor_1_resp_bits_tag;
  assign core_io_dmem_resp_bits_cmd = dcArb_io_requestor_1_resp_bits_cmd;
  assign core_io_dmem_resp_bits_typ = dcArb_io_requestor_1_resp_bits_typ;
  assign core_io_dmem_resp_bits_data = dcArb_io_requestor_1_resp_bits_data;
  assign core_io_dmem_resp_bits_replay = dcArb_io_requestor_1_resp_bits_replay;
  assign core_io_dmem_resp_bits_has_data = dcArb_io_requestor_1_resp_bits_has_data;
  assign core_io_dmem_resp_bits_data_word_bypass = dcArb_io_requestor_1_resp_bits_data_word_bypass;
  assign core_io_dmem_resp_bits_store_data = dcArb_io_requestor_1_resp_bits_store_data;
  assign core_io_dmem_replay_next = dcArb_io_requestor_1_replay_next;
  assign core_io_dmem_xcpt_ma_ld = dcArb_io_requestor_1_xcpt_ma_ld;
  assign core_io_dmem_xcpt_ma_st = dcArb_io_requestor_1_xcpt_ma_st;
  assign core_io_dmem_xcpt_pf_ld = dcArb_io_requestor_1_xcpt_pf_ld;
  assign core_io_dmem_xcpt_pf_st = dcArb_io_requestor_1_xcpt_pf_st;
  assign core_io_dmem_ordered = dcArb_io_requestor_1_ordered;
  assign core_io_fpu_fcsr_flags_valid = FPU_3558_io_fcsr_flags_valid;
  assign core_io_fpu_fcsr_flags_bits = FPU_3558_io_fcsr_flags_bits;
  assign core_io_fpu_store_data = FPU_3558_io_store_data;
  assign core_io_fpu_toint_data = FPU_3558_io_toint_data;
  assign core_io_fpu_fcsr_rdy = FPU_3558_io_fcsr_rdy;
  assign core_io_fpu_nack_mem = FPU_3558_io_nack_mem;
  assign core_io_fpu_illegal_rm = FPU_3558_io_illegal_rm;
  assign core_io_fpu_dec_cmd = FPU_3558_io_dec_cmd;
  assign core_io_fpu_dec_ldst = FPU_3558_io_dec_ldst;
  assign core_io_fpu_dec_wen = FPU_3558_io_dec_wen;
  assign core_io_fpu_dec_ren1 = FPU_3558_io_dec_ren1;
  assign core_io_fpu_dec_ren2 = FPU_3558_io_dec_ren2;
  assign core_io_fpu_dec_ren3 = FPU_3558_io_dec_ren3;
  assign core_io_fpu_dec_swap12 = FPU_3558_io_dec_swap12;
  assign core_io_fpu_dec_swap23 = FPU_3558_io_dec_swap23;
  assign core_io_fpu_dec_single = FPU_3558_io_dec_single;
  assign core_io_fpu_dec_fromint = FPU_3558_io_dec_fromint;
  assign core_io_fpu_dec_toint = FPU_3558_io_dec_toint;
  assign core_io_fpu_dec_fastpipe = FPU_3558_io_dec_fastpipe;
  assign core_io_fpu_dec_fma = FPU_3558_io_dec_fma;
  assign core_io_fpu_dec_div = FPU_3558_io_dec_div;
  assign core_io_fpu_dec_sqrt = FPU_3558_io_dec_sqrt;
  assign core_io_fpu_dec_round = FPU_3558_io_dec_round;
  assign core_io_fpu_dec_wflags = FPU_3558_io_dec_wflags;
  assign core_io_fpu_sboard_set = FPU_3558_io_sboard_set;
  assign core_io_fpu_sboard_clr = FPU_3558_io_sboard_clr;
  assign core_io_fpu_sboard_clra = FPU_3558_io_sboard_clra;
  assign core_io_fpu_cp_req_ready = FPU_3558_io_cp_req_ready;
  assign core_io_fpu_cp_resp_valid = FPU_3558_io_cp_resp_valid;
  assign core_io_fpu_cp_resp_bits_data = FPU_3558_io_cp_resp_bits_data;
  assign core_io_fpu_cp_resp_bits_exc = FPU_3558_io_cp_resp_bits_exc;
  assign core_io_rocc_cmd_ready = GEN_9;
  assign core_io_rocc_resp_valid = GEN_10;
  assign core_io_rocc_resp_bits_rd = GEN_11;
  assign core_io_rocc_resp_bits_data = GEN_12;
  assign core_io_rocc_mem_req_valid = GEN_13;
  assign core_io_rocc_mem_req_bits_addr = GEN_14;
  assign core_io_rocc_mem_req_bits_tag = GEN_15;
  assign core_io_rocc_mem_req_bits_cmd = GEN_16;
  assign core_io_rocc_mem_req_bits_typ = GEN_17;
  assign core_io_rocc_mem_req_bits_phys = GEN_18;
  assign core_io_rocc_mem_req_bits_data = GEN_19;
  assign core_io_rocc_mem_s1_kill = GEN_20;
  assign core_io_rocc_mem_s1_data = GEN_21;
  assign core_io_rocc_mem_invalidate_lr = GEN_22;
  assign core_io_rocc_busy = GEN_23;
  assign core_io_rocc_interrupt = GEN_24;
  assign core_io_rocc_autl_acquire_valid = GEN_25;
  assign core_io_rocc_autl_acquire_bits_addr_block = GEN_26;
  assign core_io_rocc_autl_acquire_bits_client_xact_id = GEN_27;
  assign core_io_rocc_autl_acquire_bits_addr_beat = GEN_28;
  assign core_io_rocc_autl_acquire_bits_is_builtin_type = GEN_29;
  assign core_io_rocc_autl_acquire_bits_a_type = GEN_30;
  assign core_io_rocc_autl_acquire_bits_union = GEN_31;
  assign core_io_rocc_autl_acquire_bits_data = GEN_32;
  assign core_io_rocc_autl_grant_ready = GEN_33;
  assign core_io_rocc_fpu_req_valid = GEN_34;
  assign core_io_rocc_fpu_req_bits_cmd = GEN_35;
  assign core_io_rocc_fpu_req_bits_ldst = GEN_36;
  assign core_io_rocc_fpu_req_bits_wen = GEN_37;
  assign core_io_rocc_fpu_req_bits_ren1 = GEN_38;
  assign core_io_rocc_fpu_req_bits_ren2 = GEN_39;
  assign core_io_rocc_fpu_req_bits_ren3 = GEN_40;
  assign core_io_rocc_fpu_req_bits_swap12 = GEN_41;
  assign core_io_rocc_fpu_req_bits_swap23 = GEN_42;
  assign core_io_rocc_fpu_req_bits_single = GEN_43;
  assign core_io_rocc_fpu_req_bits_fromint = GEN_44;
  assign core_io_rocc_fpu_req_bits_toint = GEN_45;
  assign core_io_rocc_fpu_req_bits_fastpipe = GEN_46;
  assign core_io_rocc_fpu_req_bits_fma = GEN_47;
  assign core_io_rocc_fpu_req_bits_div = GEN_48;
  assign core_io_rocc_fpu_req_bits_sqrt = GEN_49;
  assign core_io_rocc_fpu_req_bits_round = GEN_50;
  assign core_io_rocc_fpu_req_bits_wflags = GEN_51;
  assign core_io_rocc_fpu_req_bits_rm = GEN_52;
  assign core_io_rocc_fpu_req_bits_typ = GEN_53;
  assign core_io_rocc_fpu_req_bits_in1 = GEN_54;
  assign core_io_rocc_fpu_req_bits_in2 = GEN_55;
  assign core_io_rocc_fpu_req_bits_in3 = GEN_56;
  assign core_io_rocc_fpu_resp_ready = GEN_57;
  assign icache_clk = clk;
  assign icache_reset = reset;
  assign icache_io_cpu_req_valid = core_io_imem_req_valid;
  assign icache_io_cpu_req_bits_pc = core_io_imem_req_bits_pc;
  assign icache_io_cpu_resp_ready = core_io_imem_resp_ready;
  assign icache_io_cpu_btb_update_valid = core_io_imem_btb_update_valid;
  assign icache_io_cpu_btb_update_bits_prediction_valid = core_io_imem_btb_update_bits_prediction_valid;
  assign icache_io_cpu_btb_update_bits_prediction_bits_taken = core_io_imem_btb_update_bits_prediction_bits_taken;
  assign icache_io_cpu_btb_update_bits_prediction_bits_mask = core_io_imem_btb_update_bits_prediction_bits_mask;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bridx = core_io_imem_btb_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_btb_update_bits_prediction_bits_target = core_io_imem_btb_update_bits_prediction_bits_target;
  assign icache_io_cpu_btb_update_bits_prediction_bits_entry = core_io_imem_btb_update_bits_prediction_bits_entry;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_history = core_io_imem_btb_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_btb_update_bits_prediction_bits_bht_value = core_io_imem_btb_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
  assign icache_io_cpu_btb_update_bits_target = core_io_imem_btb_update_bits_target;
  assign icache_io_cpu_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
  assign icache_io_cpu_btb_update_bits_isJump = core_io_imem_btb_update_bits_isJump;
  assign icache_io_cpu_btb_update_bits_isReturn = core_io_imem_btb_update_bits_isReturn;
  assign icache_io_cpu_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
  assign icache_io_cpu_bht_update_valid = core_io_imem_bht_update_valid;
  assign icache_io_cpu_bht_update_bits_prediction_valid = core_io_imem_bht_update_bits_prediction_valid;
  assign icache_io_cpu_bht_update_bits_prediction_bits_taken = core_io_imem_bht_update_bits_prediction_bits_taken;
  assign icache_io_cpu_bht_update_bits_prediction_bits_mask = core_io_imem_bht_update_bits_prediction_bits_mask;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bridx = core_io_imem_bht_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_bht_update_bits_prediction_bits_target = core_io_imem_bht_update_bits_prediction_bits_target;
  assign icache_io_cpu_bht_update_bits_prediction_bits_entry = core_io_imem_bht_update_bits_prediction_bits_entry;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_history = core_io_imem_bht_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_bht_update_bits_prediction_bits_bht_value = core_io_imem_bht_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
  assign icache_io_cpu_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
  assign icache_io_cpu_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
  assign icache_io_cpu_ras_update_valid = core_io_imem_ras_update_valid;
  assign icache_io_cpu_ras_update_bits_isCall = core_io_imem_ras_update_bits_isCall;
  assign icache_io_cpu_ras_update_bits_isReturn = core_io_imem_ras_update_bits_isReturn;
  assign icache_io_cpu_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
  assign icache_io_cpu_ras_update_bits_prediction_valid = core_io_imem_ras_update_bits_prediction_valid;
  assign icache_io_cpu_ras_update_bits_prediction_bits_taken = core_io_imem_ras_update_bits_prediction_bits_taken;
  assign icache_io_cpu_ras_update_bits_prediction_bits_mask = core_io_imem_ras_update_bits_prediction_bits_mask;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bridx = core_io_imem_ras_update_bits_prediction_bits_bridx;
  assign icache_io_cpu_ras_update_bits_prediction_bits_target = core_io_imem_ras_update_bits_prediction_bits_target;
  assign icache_io_cpu_ras_update_bits_prediction_bits_entry = core_io_imem_ras_update_bits_prediction_bits_entry;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_history = core_io_imem_ras_update_bits_prediction_bits_bht_history;
  assign icache_io_cpu_ras_update_bits_prediction_bits_bht_value = core_io_imem_ras_update_bits_prediction_bits_bht_value;
  assign icache_io_cpu_flush_icache = core_io_imem_flush_icache;
  assign icache_io_cpu_flush_tlb = core_io_imem_flush_tlb;
  assign icache_io_ptw_req_ready = PTW_3559_io_requestor_0_req_ready;
  assign icache_io_ptw_resp_valid = PTW_3559_io_requestor_0_resp_valid;
  assign icache_io_ptw_resp_bits_pte_ppn = PTW_3559_io_requestor_0_resp_bits_pte_ppn;
  assign icache_io_ptw_resp_bits_pte_reserved_for_software = PTW_3559_io_requestor_0_resp_bits_pte_reserved_for_software;
  assign icache_io_ptw_resp_bits_pte_d = PTW_3559_io_requestor_0_resp_bits_pte_d;
  assign icache_io_ptw_resp_bits_pte_r = PTW_3559_io_requestor_0_resp_bits_pte_r;
  assign icache_io_ptw_resp_bits_pte_typ = PTW_3559_io_requestor_0_resp_bits_pte_typ;
  assign icache_io_ptw_resp_bits_pte_v = PTW_3559_io_requestor_0_resp_bits_pte_v;
  assign icache_io_ptw_status_debug = PTW_3559_io_requestor_0_status_debug;
  assign icache_io_ptw_status_prv = PTW_3559_io_requestor_0_status_prv;
  assign icache_io_ptw_status_sd = PTW_3559_io_requestor_0_status_sd;
  assign icache_io_ptw_status_zero3 = PTW_3559_io_requestor_0_status_zero3;
  assign icache_io_ptw_status_sd_rv32 = PTW_3559_io_requestor_0_status_sd_rv32;
  assign icache_io_ptw_status_zero2 = PTW_3559_io_requestor_0_status_zero2;
  assign icache_io_ptw_status_vm = PTW_3559_io_requestor_0_status_vm;
  assign icache_io_ptw_status_zero1 = PTW_3559_io_requestor_0_status_zero1;
  assign icache_io_ptw_status_pum = PTW_3559_io_requestor_0_status_pum;
  assign icache_io_ptw_status_mprv = PTW_3559_io_requestor_0_status_mprv;
  assign icache_io_ptw_status_xs = PTW_3559_io_requestor_0_status_xs;
  assign icache_io_ptw_status_fs = PTW_3559_io_requestor_0_status_fs;
  assign icache_io_ptw_status_mpp = PTW_3559_io_requestor_0_status_mpp;
  assign icache_io_ptw_status_hpp = PTW_3559_io_requestor_0_status_hpp;
  assign icache_io_ptw_status_spp = PTW_3559_io_requestor_0_status_spp;
  assign icache_io_ptw_status_mpie = PTW_3559_io_requestor_0_status_mpie;
  assign icache_io_ptw_status_hpie = PTW_3559_io_requestor_0_status_hpie;
  assign icache_io_ptw_status_spie = PTW_3559_io_requestor_0_status_spie;
  assign icache_io_ptw_status_upie = PTW_3559_io_requestor_0_status_upie;
  assign icache_io_ptw_status_mie = PTW_3559_io_requestor_0_status_mie;
  assign icache_io_ptw_status_hie = PTW_3559_io_requestor_0_status_hie;
  assign icache_io_ptw_status_sie = PTW_3559_io_requestor_0_status_sie;
  assign icache_io_ptw_status_uie = PTW_3559_io_requestor_0_status_uie;
  assign icache_io_ptw_invalidate = PTW_3559_io_requestor_0_invalidate;
  assign icache_io_mem_acquire_ready = uncachedArb_io_in_0_acquire_ready;
  assign icache_io_mem_grant_valid = uncachedArb_io_in_0_grant_valid;
  assign icache_io_mem_grant_bits_addr_beat = uncachedArb_io_in_0_grant_bits_addr_beat;
  assign icache_io_mem_grant_bits_client_xact_id = uncachedArb_io_in_0_grant_bits_client_xact_id;
  assign icache_io_mem_grant_bits_manager_xact_id = uncachedArb_io_in_0_grant_bits_manager_xact_id;
  assign icache_io_mem_grant_bits_is_builtin_type = uncachedArb_io_in_0_grant_bits_is_builtin_type;
  assign icache_io_mem_grant_bits_g_type = uncachedArb_io_in_0_grant_bits_g_type;
  assign icache_io_mem_grant_bits_data = uncachedArb_io_in_0_grant_bits_data;
  assign HellaCache_3557_clk = clk;
  assign HellaCache_3557_reset = reset;
  assign HellaCache_3557_io_cpu_req_valid = dcArb_io_mem_req_valid;
  assign HellaCache_3557_io_cpu_req_bits_addr = dcArb_io_mem_req_bits_addr;
  assign HellaCache_3557_io_cpu_req_bits_tag = dcArb_io_mem_req_bits_tag;
  assign HellaCache_3557_io_cpu_req_bits_cmd = dcArb_io_mem_req_bits_cmd;
  assign HellaCache_3557_io_cpu_req_bits_typ = dcArb_io_mem_req_bits_typ;
  assign HellaCache_3557_io_cpu_req_bits_phys = dcArb_io_mem_req_bits_phys;
  assign HellaCache_3557_io_cpu_req_bits_data = dcArb_io_mem_req_bits_data;
  assign HellaCache_3557_io_cpu_s1_kill = dcArb_io_mem_s1_kill;
  assign HellaCache_3557_io_cpu_s1_data = dcArb_io_mem_s1_data;
  assign HellaCache_3557_io_cpu_invalidate_lr = dcArb_io_mem_invalidate_lr;
  assign HellaCache_3557_io_ptw_req_ready = PTW_3559_io_requestor_1_req_ready;
  assign HellaCache_3557_io_ptw_resp_valid = PTW_3559_io_requestor_1_resp_valid;
  assign HellaCache_3557_io_ptw_resp_bits_pte_ppn = PTW_3559_io_requestor_1_resp_bits_pte_ppn;
  assign HellaCache_3557_io_ptw_resp_bits_pte_reserved_for_software = PTW_3559_io_requestor_1_resp_bits_pte_reserved_for_software;
  assign HellaCache_3557_io_ptw_resp_bits_pte_d = PTW_3559_io_requestor_1_resp_bits_pte_d;
  assign HellaCache_3557_io_ptw_resp_bits_pte_r = PTW_3559_io_requestor_1_resp_bits_pte_r;
  assign HellaCache_3557_io_ptw_resp_bits_pte_typ = PTW_3559_io_requestor_1_resp_bits_pte_typ;
  assign HellaCache_3557_io_ptw_resp_bits_pte_v = PTW_3559_io_requestor_1_resp_bits_pte_v;
  assign HellaCache_3557_io_ptw_status_debug = PTW_3559_io_requestor_1_status_debug;
  assign HellaCache_3557_io_ptw_status_prv = PTW_3559_io_requestor_1_status_prv;
  assign HellaCache_3557_io_ptw_status_sd = PTW_3559_io_requestor_1_status_sd;
  assign HellaCache_3557_io_ptw_status_zero3 = PTW_3559_io_requestor_1_status_zero3;
  assign HellaCache_3557_io_ptw_status_sd_rv32 = PTW_3559_io_requestor_1_status_sd_rv32;
  assign HellaCache_3557_io_ptw_status_zero2 = PTW_3559_io_requestor_1_status_zero2;
  assign HellaCache_3557_io_ptw_status_vm = PTW_3559_io_requestor_1_status_vm;
  assign HellaCache_3557_io_ptw_status_zero1 = PTW_3559_io_requestor_1_status_zero1;
  assign HellaCache_3557_io_ptw_status_pum = PTW_3559_io_requestor_1_status_pum;
  assign HellaCache_3557_io_ptw_status_mprv = PTW_3559_io_requestor_1_status_mprv;
  assign HellaCache_3557_io_ptw_status_xs = PTW_3559_io_requestor_1_status_xs;
  assign HellaCache_3557_io_ptw_status_fs = PTW_3559_io_requestor_1_status_fs;
  assign HellaCache_3557_io_ptw_status_mpp = PTW_3559_io_requestor_1_status_mpp;
  assign HellaCache_3557_io_ptw_status_hpp = PTW_3559_io_requestor_1_status_hpp;
  assign HellaCache_3557_io_ptw_status_spp = PTW_3559_io_requestor_1_status_spp;
  assign HellaCache_3557_io_ptw_status_mpie = PTW_3559_io_requestor_1_status_mpie;
  assign HellaCache_3557_io_ptw_status_hpie = PTW_3559_io_requestor_1_status_hpie;
  assign HellaCache_3557_io_ptw_status_spie = PTW_3559_io_requestor_1_status_spie;
  assign HellaCache_3557_io_ptw_status_upie = PTW_3559_io_requestor_1_status_upie;
  assign HellaCache_3557_io_ptw_status_mie = PTW_3559_io_requestor_1_status_mie;
  assign HellaCache_3557_io_ptw_status_hie = PTW_3559_io_requestor_1_status_hie;
  assign HellaCache_3557_io_ptw_status_sie = PTW_3559_io_requestor_1_status_sie;
  assign HellaCache_3557_io_ptw_status_uie = PTW_3559_io_requestor_1_status_uie;
  assign HellaCache_3557_io_ptw_invalidate = PTW_3559_io_requestor_1_invalidate;
  assign HellaCache_3557_io_mem_acquire_ready = io_cached_0_acquire_ready;
  assign HellaCache_3557_io_mem_probe_valid = io_cached_0_probe_valid;
  assign HellaCache_3557_io_mem_probe_bits_addr_block = io_cached_0_probe_bits_addr_block;
  assign HellaCache_3557_io_mem_probe_bits_p_type = io_cached_0_probe_bits_p_type;
  assign HellaCache_3557_io_mem_release_ready = io_cached_0_release_ready;
  assign HellaCache_3557_io_mem_grant_valid = io_cached_0_grant_valid;
  assign HellaCache_3557_io_mem_grant_bits_addr_beat = io_cached_0_grant_bits_addr_beat;
  assign HellaCache_3557_io_mem_grant_bits_client_xact_id = io_cached_0_grant_bits_client_xact_id;
  assign HellaCache_3557_io_mem_grant_bits_manager_xact_id = io_cached_0_grant_bits_manager_xact_id;
  assign HellaCache_3557_io_mem_grant_bits_is_builtin_type = io_cached_0_grant_bits_is_builtin_type;
  assign HellaCache_3557_io_mem_grant_bits_g_type = io_cached_0_grant_bits_g_type;
  assign HellaCache_3557_io_mem_grant_bits_data = io_cached_0_grant_bits_data;
  assign HellaCache_3557_io_mem_grant_bits_manager_id = io_cached_0_grant_bits_manager_id;
  assign HellaCache_3557_io_mem_finish_ready = io_cached_0_finish_ready;
  assign FPU_3558_clk = clk;
  assign FPU_3558_reset = reset;
  assign FPU_3558_io_inst = core_io_fpu_inst;
  assign FPU_3558_io_fromint_data = core_io_fpu_fromint_data;
  assign FPU_3558_io_fcsr_rm = core_io_fpu_fcsr_rm;
  assign FPU_3558_io_dmem_resp_val = core_io_fpu_dmem_resp_val;
  assign FPU_3558_io_dmem_resp_type = core_io_fpu_dmem_resp_type;
  assign FPU_3558_io_dmem_resp_tag = core_io_fpu_dmem_resp_tag;
  assign FPU_3558_io_dmem_resp_data = core_io_fpu_dmem_resp_data;
  assign FPU_3558_io_valid = core_io_fpu_valid;
  assign FPU_3558_io_killx = core_io_fpu_killx;
  assign FPU_3558_io_killm = core_io_fpu_killm;
  assign FPU_3558_io_cp_req_valid = 1'h0;
  assign FPU_3558_io_cp_req_bits_cmd = core_io_fpu_cp_req_bits_cmd;
  assign FPU_3558_io_cp_req_bits_ldst = core_io_fpu_cp_req_bits_ldst;
  assign FPU_3558_io_cp_req_bits_wen = core_io_fpu_cp_req_bits_wen;
  assign FPU_3558_io_cp_req_bits_ren1 = core_io_fpu_cp_req_bits_ren1;
  assign FPU_3558_io_cp_req_bits_ren2 = core_io_fpu_cp_req_bits_ren2;
  assign FPU_3558_io_cp_req_bits_ren3 = core_io_fpu_cp_req_bits_ren3;
  assign FPU_3558_io_cp_req_bits_swap12 = core_io_fpu_cp_req_bits_swap12;
  assign FPU_3558_io_cp_req_bits_swap23 = core_io_fpu_cp_req_bits_swap23;
  assign FPU_3558_io_cp_req_bits_single = core_io_fpu_cp_req_bits_single;
  assign FPU_3558_io_cp_req_bits_fromint = core_io_fpu_cp_req_bits_fromint;
  assign FPU_3558_io_cp_req_bits_toint = core_io_fpu_cp_req_bits_toint;
  assign FPU_3558_io_cp_req_bits_fastpipe = core_io_fpu_cp_req_bits_fastpipe;
  assign FPU_3558_io_cp_req_bits_fma = core_io_fpu_cp_req_bits_fma;
  assign FPU_3558_io_cp_req_bits_div = core_io_fpu_cp_req_bits_div;
  assign FPU_3558_io_cp_req_bits_sqrt = core_io_fpu_cp_req_bits_sqrt;
  assign FPU_3558_io_cp_req_bits_round = core_io_fpu_cp_req_bits_round;
  assign FPU_3558_io_cp_req_bits_wflags = core_io_fpu_cp_req_bits_wflags;
  assign FPU_3558_io_cp_req_bits_rm = core_io_fpu_cp_req_bits_rm;
  assign FPU_3558_io_cp_req_bits_typ = core_io_fpu_cp_req_bits_typ;
  assign FPU_3558_io_cp_req_bits_in1 = core_io_fpu_cp_req_bits_in1;
  assign FPU_3558_io_cp_req_bits_in2 = core_io_fpu_cp_req_bits_in2;
  assign FPU_3558_io_cp_req_bits_in3 = core_io_fpu_cp_req_bits_in3;
  assign FPU_3558_io_cp_resp_ready = 1'h0;
  assign uncachedArb_clk = clk;
  assign uncachedArb_reset = reset;
  assign uncachedArb_io_in_0_acquire_valid = icache_io_mem_acquire_valid;
  assign uncachedArb_io_in_0_acquire_bits_addr_block = icache_io_mem_acquire_bits_addr_block;
  assign uncachedArb_io_in_0_acquire_bits_client_xact_id = icache_io_mem_acquire_bits_client_xact_id;
  assign uncachedArb_io_in_0_acquire_bits_addr_beat = icache_io_mem_acquire_bits_addr_beat;
  assign uncachedArb_io_in_0_acquire_bits_is_builtin_type = icache_io_mem_acquire_bits_is_builtin_type;
  assign uncachedArb_io_in_0_acquire_bits_a_type = icache_io_mem_acquire_bits_a_type;
  assign uncachedArb_io_in_0_acquire_bits_union = icache_io_mem_acquire_bits_union;
  assign uncachedArb_io_in_0_acquire_bits_data = icache_io_mem_acquire_bits_data;
  assign uncachedArb_io_in_0_grant_ready = icache_io_mem_grant_ready;
  assign uncachedArb_io_out_acquire_ready = io_uncached_0_acquire_ready;
  assign uncachedArb_io_out_grant_valid = io_uncached_0_grant_valid;
  assign uncachedArb_io_out_grant_bits_addr_beat = io_uncached_0_grant_bits_addr_beat;
  assign uncachedArb_io_out_grant_bits_client_xact_id = io_uncached_0_grant_bits_client_xact_id;
  assign uncachedArb_io_out_grant_bits_manager_xact_id = io_uncached_0_grant_bits_manager_xact_id;
  assign uncachedArb_io_out_grant_bits_is_builtin_type = io_uncached_0_grant_bits_is_builtin_type;
  assign uncachedArb_io_out_grant_bits_g_type = io_uncached_0_grant_bits_g_type;
  assign uncachedArb_io_out_grant_bits_data = io_uncached_0_grant_bits_data;
  assign PTW_3559_clk = clk;
  assign PTW_3559_reset = reset;
  assign PTW_3559_io_requestor_0_req_valid = icache_io_ptw_req_valid;
  assign PTW_3559_io_requestor_0_req_bits_addr = icache_io_ptw_req_bits_addr;
  assign PTW_3559_io_requestor_0_req_bits_prv = icache_io_ptw_req_bits_prv;
  assign PTW_3559_io_requestor_0_req_bits_store = icache_io_ptw_req_bits_store;
  assign PTW_3559_io_requestor_0_req_bits_fetch = icache_io_ptw_req_bits_fetch;
  assign PTW_3559_io_requestor_1_req_valid = HellaCache_3557_io_ptw_req_valid;
  assign PTW_3559_io_requestor_1_req_bits_addr = HellaCache_3557_io_ptw_req_bits_addr;
  assign PTW_3559_io_requestor_1_req_bits_prv = HellaCache_3557_io_ptw_req_bits_prv;
  assign PTW_3559_io_requestor_1_req_bits_store = HellaCache_3557_io_ptw_req_bits_store;
  assign PTW_3559_io_requestor_1_req_bits_fetch = HellaCache_3557_io_ptw_req_bits_fetch;
  assign PTW_3559_io_mem_req_ready = dcArb_io_requestor_0_req_ready;
  assign PTW_3559_io_mem_s2_nack = dcArb_io_requestor_0_s2_nack;
  assign PTW_3559_io_mem_resp_valid = dcArb_io_requestor_0_resp_valid;
  assign PTW_3559_io_mem_resp_bits_addr = dcArb_io_requestor_0_resp_bits_addr;
  assign PTW_3559_io_mem_resp_bits_tag = dcArb_io_requestor_0_resp_bits_tag;
  assign PTW_3559_io_mem_resp_bits_cmd = dcArb_io_requestor_0_resp_bits_cmd;
  assign PTW_3559_io_mem_resp_bits_typ = dcArb_io_requestor_0_resp_bits_typ;
  assign PTW_3559_io_mem_resp_bits_data = dcArb_io_requestor_0_resp_bits_data;
  assign PTW_3559_io_mem_resp_bits_replay = dcArb_io_requestor_0_resp_bits_replay;
  assign PTW_3559_io_mem_resp_bits_has_data = dcArb_io_requestor_0_resp_bits_has_data;
  assign PTW_3559_io_mem_resp_bits_data_word_bypass = dcArb_io_requestor_0_resp_bits_data_word_bypass;
  assign PTW_3559_io_mem_resp_bits_store_data = dcArb_io_requestor_0_resp_bits_store_data;
  assign PTW_3559_io_mem_replay_next = dcArb_io_requestor_0_replay_next;
  assign PTW_3559_io_mem_xcpt_ma_ld = dcArb_io_requestor_0_xcpt_ma_ld;
  assign PTW_3559_io_mem_xcpt_ma_st = dcArb_io_requestor_0_xcpt_ma_st;
  assign PTW_3559_io_mem_xcpt_pf_ld = dcArb_io_requestor_0_xcpt_pf_ld;
  assign PTW_3559_io_mem_xcpt_pf_st = dcArb_io_requestor_0_xcpt_pf_st;
  assign PTW_3559_io_mem_ordered = dcArb_io_requestor_0_ordered;
  assign PTW_3559_io_dpath_ptbr = core_io_ptw_ptbr;
  assign PTW_3559_io_dpath_invalidate = core_io_ptw_invalidate;
  assign PTW_3559_io_dpath_status_debug = core_io_ptw_status_debug;
  assign PTW_3559_io_dpath_status_prv = core_io_ptw_status_prv;
  assign PTW_3559_io_dpath_status_sd = core_io_ptw_status_sd;
  assign PTW_3559_io_dpath_status_zero3 = core_io_ptw_status_zero3;
  assign PTW_3559_io_dpath_status_sd_rv32 = core_io_ptw_status_sd_rv32;
  assign PTW_3559_io_dpath_status_zero2 = core_io_ptw_status_zero2;
  assign PTW_3559_io_dpath_status_vm = core_io_ptw_status_vm;
  assign PTW_3559_io_dpath_status_zero1 = core_io_ptw_status_zero1;
  assign PTW_3559_io_dpath_status_pum = core_io_ptw_status_pum;
  assign PTW_3559_io_dpath_status_mprv = core_io_ptw_status_mprv;
  assign PTW_3559_io_dpath_status_xs = core_io_ptw_status_xs;
  assign PTW_3559_io_dpath_status_fs = core_io_ptw_status_fs;
  assign PTW_3559_io_dpath_status_mpp = core_io_ptw_status_mpp;
  assign PTW_3559_io_dpath_status_hpp = core_io_ptw_status_hpp;
  assign PTW_3559_io_dpath_status_spp = core_io_ptw_status_spp;
  assign PTW_3559_io_dpath_status_mpie = core_io_ptw_status_mpie;
  assign PTW_3559_io_dpath_status_hpie = core_io_ptw_status_hpie;
  assign PTW_3559_io_dpath_status_spie = core_io_ptw_status_spie;
  assign PTW_3559_io_dpath_status_upie = core_io_ptw_status_upie;
  assign PTW_3559_io_dpath_status_mie = core_io_ptw_status_mie;
  assign PTW_3559_io_dpath_status_hie = core_io_ptw_status_hie;
  assign PTW_3559_io_dpath_status_sie = core_io_ptw_status_sie;
  assign PTW_3559_io_dpath_status_uie = core_io_ptw_status_uie;
  assign dcArb_clk = clk;
  assign dcArb_reset = reset;
  assign dcArb_io_requestor_0_req_valid = PTW_3559_io_mem_req_valid;
  assign dcArb_io_requestor_0_req_bits_addr = PTW_3559_io_mem_req_bits_addr;
  assign dcArb_io_requestor_0_req_bits_tag = PTW_3559_io_mem_req_bits_tag;
  assign dcArb_io_requestor_0_req_bits_cmd = PTW_3559_io_mem_req_bits_cmd;
  assign dcArb_io_requestor_0_req_bits_typ = PTW_3559_io_mem_req_bits_typ;
  assign dcArb_io_requestor_0_req_bits_phys = PTW_3559_io_mem_req_bits_phys;
  assign dcArb_io_requestor_0_req_bits_data = PTW_3559_io_mem_req_bits_data;
  assign dcArb_io_requestor_0_s1_kill = PTW_3559_io_mem_s1_kill;
  assign dcArb_io_requestor_0_s1_data = PTW_3559_io_mem_s1_data;
  assign dcArb_io_requestor_0_invalidate_lr = PTW_3559_io_mem_invalidate_lr;
  assign dcArb_io_requestor_1_req_valid = core_io_dmem_req_valid;
  assign dcArb_io_requestor_1_req_bits_addr = core_io_dmem_req_bits_addr;
  assign dcArb_io_requestor_1_req_bits_tag = core_io_dmem_req_bits_tag;
  assign dcArb_io_requestor_1_req_bits_cmd = core_io_dmem_req_bits_cmd;
  assign dcArb_io_requestor_1_req_bits_typ = core_io_dmem_req_bits_typ;
  assign dcArb_io_requestor_1_req_bits_phys = core_io_dmem_req_bits_phys;
  assign dcArb_io_requestor_1_req_bits_data = core_io_dmem_req_bits_data;
  assign dcArb_io_requestor_1_s1_kill = core_io_dmem_s1_kill;
  assign dcArb_io_requestor_1_s1_data = core_io_dmem_s1_data;
  assign dcArb_io_requestor_1_invalidate_lr = core_io_dmem_invalidate_lr;
  assign dcArb_io_mem_req_ready = HellaCache_3557_io_cpu_req_ready;
  assign dcArb_io_mem_s2_nack = HellaCache_3557_io_cpu_s2_nack;
  assign dcArb_io_mem_resp_valid = HellaCache_3557_io_cpu_resp_valid;
  assign dcArb_io_mem_resp_bits_addr = HellaCache_3557_io_cpu_resp_bits_addr;
  assign dcArb_io_mem_resp_bits_tag = HellaCache_3557_io_cpu_resp_bits_tag;
  assign dcArb_io_mem_resp_bits_cmd = HellaCache_3557_io_cpu_resp_bits_cmd;
  assign dcArb_io_mem_resp_bits_typ = HellaCache_3557_io_cpu_resp_bits_typ;
  assign dcArb_io_mem_resp_bits_data = HellaCache_3557_io_cpu_resp_bits_data;
  assign dcArb_io_mem_resp_bits_replay = HellaCache_3557_io_cpu_resp_bits_replay;
  assign dcArb_io_mem_resp_bits_has_data = HellaCache_3557_io_cpu_resp_bits_has_data;
  assign dcArb_io_mem_resp_bits_data_word_bypass = HellaCache_3557_io_cpu_resp_bits_data_word_bypass;
  assign dcArb_io_mem_resp_bits_store_data = HellaCache_3557_io_cpu_resp_bits_store_data;
  assign dcArb_io_mem_replay_next = HellaCache_3557_io_cpu_replay_next;
  assign dcArb_io_mem_xcpt_ma_ld = HellaCache_3557_io_cpu_xcpt_ma_ld;
  assign dcArb_io_mem_xcpt_ma_st = HellaCache_3557_io_cpu_xcpt_ma_st;
  assign dcArb_io_mem_xcpt_pf_ld = HellaCache_3557_io_cpu_xcpt_pf_ld;
  assign dcArb_io_mem_xcpt_pf_st = HellaCache_3557_io_cpu_xcpt_pf_st;
  assign dcArb_io_mem_ordered = HellaCache_3557_io_cpu_ordered;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_58 = {1{$random}};
  GEN_0 = GEN_58[0:0];
  GEN_59 = {1{$random}};
  GEN_1 = GEN_59[1:0];
  GEN_60 = {1{$random}};
  GEN_2 = GEN_60[0:0];
  GEN_61 = {1{$random}};
  GEN_3 = GEN_61[2:0];
  GEN_62 = {1{$random}};
  GEN_4 = GEN_62[31:0];
  GEN_63 = {1{$random}};
  GEN_5 = GEN_63[31:0];
  GEN_64 = {1{$random}};
  GEN_6 = GEN_64[31:0];
  GEN_65 = {1{$random}};
  GEN_7 = GEN_65[1:0];
  GEN_66 = {1{$random}};
  GEN_8 = GEN_66[0:0];
  GEN_67 = {1{$random}};
  GEN_9 = GEN_67[0:0];
  GEN_68 = {1{$random}};
  GEN_10 = GEN_68[0:0];
  GEN_69 = {1{$random}};
  GEN_11 = GEN_69[4:0];
  GEN_70 = {2{$random}};
  GEN_12 = GEN_70[63:0];
  GEN_71 = {1{$random}};
  GEN_13 = GEN_71[0:0];
  GEN_72 = {2{$random}};
  GEN_14 = GEN_72[39:0];
  GEN_73 = {1{$random}};
  GEN_15 = GEN_73[8:0];
  GEN_74 = {1{$random}};
  GEN_16 = GEN_74[4:0];
  GEN_75 = {1{$random}};
  GEN_17 = GEN_75[2:0];
  GEN_76 = {1{$random}};
  GEN_18 = GEN_76[0:0];
  GEN_77 = {2{$random}};
  GEN_19 = GEN_77[63:0];
  GEN_78 = {1{$random}};
  GEN_20 = GEN_78[0:0];
  GEN_79 = {2{$random}};
  GEN_21 = GEN_79[63:0];
  GEN_80 = {1{$random}};
  GEN_22 = GEN_80[0:0];
  GEN_81 = {1{$random}};
  GEN_23 = GEN_81[0:0];
  GEN_82 = {1{$random}};
  GEN_24 = GEN_82[0:0];
  GEN_83 = {1{$random}};
  GEN_25 = GEN_83[0:0];
  GEN_84 = {1{$random}};
  GEN_26 = GEN_84[25:0];
  GEN_85 = {1{$random}};
  GEN_27 = GEN_85[1:0];
  GEN_86 = {1{$random}};
  GEN_28 = GEN_86[2:0];
  GEN_87 = {1{$random}};
  GEN_29 = GEN_87[0:0];
  GEN_88 = {1{$random}};
  GEN_30 = GEN_88[2:0];
  GEN_89 = {1{$random}};
  GEN_31 = GEN_89[11:0];
  GEN_90 = {2{$random}};
  GEN_32 = GEN_90[63:0];
  GEN_91 = {1{$random}};
  GEN_33 = GEN_91[0:0];
  GEN_92 = {1{$random}};
  GEN_34 = GEN_92[0:0];
  GEN_93 = {1{$random}};
  GEN_35 = GEN_93[4:0];
  GEN_94 = {1{$random}};
  GEN_36 = GEN_94[0:0];
  GEN_95 = {1{$random}};
  GEN_37 = GEN_95[0:0];
  GEN_96 = {1{$random}};
  GEN_38 = GEN_96[0:0];
  GEN_97 = {1{$random}};
  GEN_39 = GEN_97[0:0];
  GEN_98 = {1{$random}};
  GEN_40 = GEN_98[0:0];
  GEN_99 = {1{$random}};
  GEN_41 = GEN_99[0:0];
  GEN_100 = {1{$random}};
  GEN_42 = GEN_100[0:0];
  GEN_101 = {1{$random}};
  GEN_43 = GEN_101[0:0];
  GEN_102 = {1{$random}};
  GEN_44 = GEN_102[0:0];
  GEN_103 = {1{$random}};
  GEN_45 = GEN_103[0:0];
  GEN_104 = {1{$random}};
  GEN_46 = GEN_104[0:0];
  GEN_105 = {1{$random}};
  GEN_47 = GEN_105[0:0];
  GEN_106 = {1{$random}};
  GEN_48 = GEN_106[0:0];
  GEN_107 = {1{$random}};
  GEN_49 = GEN_107[0:0];
  GEN_108 = {1{$random}};
  GEN_50 = GEN_108[0:0];
  GEN_109 = {1{$random}};
  GEN_51 = GEN_109[0:0];
  GEN_110 = {1{$random}};
  GEN_52 = GEN_110[2:0];
  GEN_111 = {1{$random}};
  GEN_53 = GEN_111[1:0];
  GEN_112 = {3{$random}};
  GEN_54 = GEN_112[64:0];
  GEN_113 = {3{$random}};
  GEN_55 = GEN_113[64:0];
  GEN_114 = {3{$random}};
  GEN_56 = GEN_114[64:0];
  GEN_115 = {1{$random}};
  GEN_57 = GEN_115[0:0];
  end
`endif
endmodule
module Top(
  input   clk,
  input   reset,
  output  io_host_clk,
  output  io_host_clk_edge,
  output  io_host_in_ready,
  input   io_host_in_valid,
  input  [15:0] io_host_in_bits,
  input   io_host_out_ready,
  output  io_host_out_valid,
  output [15:0] io_host_out_bits,
  input   io_mem_axi_0_aw_ready,
  output  io_mem_axi_0_aw_valid,
  output [31:0] io_mem_axi_0_aw_bits_addr,
  output [7:0] io_mem_axi_0_aw_bits_len,
  output [2:0] io_mem_axi_0_aw_bits_size,
  output [1:0] io_mem_axi_0_aw_bits_burst,
  output  io_mem_axi_0_aw_bits_lock,
  output [3:0] io_mem_axi_0_aw_bits_cache,
  output [2:0] io_mem_axi_0_aw_bits_prot,
  output [3:0] io_mem_axi_0_aw_bits_qos,
  output [3:0] io_mem_axi_0_aw_bits_region,
  output [4:0] io_mem_axi_0_aw_bits_id,
  output  io_mem_axi_0_aw_bits_user,
  input   io_mem_axi_0_w_ready,
  output  io_mem_axi_0_w_valid,
  output [63:0] io_mem_axi_0_w_bits_data,
  output  io_mem_axi_0_w_bits_last,
  output [4:0] io_mem_axi_0_w_bits_id,
  output [7:0] io_mem_axi_0_w_bits_strb,
  output  io_mem_axi_0_w_bits_user,
  output  io_mem_axi_0_b_ready,
  input   io_mem_axi_0_b_valid,
  input  [1:0] io_mem_axi_0_b_bits_resp,
  input  [4:0] io_mem_axi_0_b_bits_id,
  input   io_mem_axi_0_b_bits_user,
  input   io_mem_axi_0_ar_ready,
  output  io_mem_axi_0_ar_valid,
  output [31:0] io_mem_axi_0_ar_bits_addr,
  output [7:0] io_mem_axi_0_ar_bits_len,
  output [2:0] io_mem_axi_0_ar_bits_size,
  output [1:0] io_mem_axi_0_ar_bits_burst,
  output  io_mem_axi_0_ar_bits_lock,
  output [3:0] io_mem_axi_0_ar_bits_cache,
  output [2:0] io_mem_axi_0_ar_bits_prot,
  output [3:0] io_mem_axi_0_ar_bits_qos,
  output [3:0] io_mem_axi_0_ar_bits_region,
  output [4:0] io_mem_axi_0_ar_bits_id,
  output  io_mem_axi_0_ar_bits_user,
  output  io_mem_axi_0_r_ready,
  input   io_mem_axi_0_r_valid,
  input  [1:0] io_mem_axi_0_r_bits_resp,
  input  [63:0] io_mem_axi_0_r_bits_data,
  input   io_mem_axi_0_r_bits_last,
  input  [4:0] io_mem_axi_0_r_bits_id,
  input   io_mem_axi_0_r_bits_user,
  input   io_interrupts_0,
  input   io_interrupts_1,
  output  io_debug_req_ready,
  input   io_debug_req_valid,
  input  [4:0] io_debug_req_bits_addr,
  input  [1:0] io_debug_req_bits_op,
  input  [33:0] io_debug_req_bits_data,
  input   io_debug_resp_ready,
  output  io_debug_resp_valid,
  output [1:0] io_debug_resp_bits_resp,
  output [33:0] io_debug_resp_bits_data
);
  wire  uncore_clk;
  wire  uncore_reset;
  wire  uncore_io_host_clk;
  wire  uncore_io_host_clk_edge;
  wire  uncore_io_host_in_ready;
  wire  uncore_io_host_in_valid;
  wire [15:0] uncore_io_host_in_bits;
  wire  uncore_io_host_out_ready;
  wire  uncore_io_host_out_valid;
  wire [15:0] uncore_io_host_out_bits;
  wire  uncore_io_mem_axi_0_aw_ready;
  wire  uncore_io_mem_axi_0_aw_valid;
  wire [31:0] uncore_io_mem_axi_0_aw_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_aw_bits_len;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_size;
  wire [1:0] uncore_io_mem_axi_0_aw_bits_burst;
  wire  uncore_io_mem_axi_0_aw_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_aw_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_aw_bits_region;
  wire [4:0] uncore_io_mem_axi_0_aw_bits_id;
  wire  uncore_io_mem_axi_0_aw_bits_user;
  wire  uncore_io_mem_axi_0_w_ready;
  wire  uncore_io_mem_axi_0_w_valid;
  wire [63:0] uncore_io_mem_axi_0_w_bits_data;
  wire  uncore_io_mem_axi_0_w_bits_last;
  wire [4:0] uncore_io_mem_axi_0_w_bits_id;
  wire [7:0] uncore_io_mem_axi_0_w_bits_strb;
  wire  uncore_io_mem_axi_0_w_bits_user;
  wire  uncore_io_mem_axi_0_b_ready;
  wire  uncore_io_mem_axi_0_b_valid;
  wire [1:0] uncore_io_mem_axi_0_b_bits_resp;
  wire [4:0] uncore_io_mem_axi_0_b_bits_id;
  wire  uncore_io_mem_axi_0_b_bits_user;
  wire  uncore_io_mem_axi_0_ar_ready;
  wire  uncore_io_mem_axi_0_ar_valid;
  wire [31:0] uncore_io_mem_axi_0_ar_bits_addr;
  wire [7:0] uncore_io_mem_axi_0_ar_bits_len;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_size;
  wire [1:0] uncore_io_mem_axi_0_ar_bits_burst;
  wire  uncore_io_mem_axi_0_ar_bits_lock;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_cache;
  wire [2:0] uncore_io_mem_axi_0_ar_bits_prot;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_qos;
  wire [3:0] uncore_io_mem_axi_0_ar_bits_region;
  wire [4:0] uncore_io_mem_axi_0_ar_bits_id;
  wire  uncore_io_mem_axi_0_ar_bits_user;
  wire  uncore_io_mem_axi_0_r_ready;
  wire  uncore_io_mem_axi_0_r_valid;
  wire [1:0] uncore_io_mem_axi_0_r_bits_resp;
  wire [63:0] uncore_io_mem_axi_0_r_bits_data;
  wire  uncore_io_mem_axi_0_r_bits_last;
  wire [4:0] uncore_io_mem_axi_0_r_bits_id;
  wire  uncore_io_mem_axi_0_r_bits_user;
  wire  uncore_io_tiles_cached_0_acquire_ready;
  wire  uncore_io_tiles_cached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_cached_0_acquire_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_cached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_cached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_cached_0_acquire_bits_data;
  wire  uncore_io_tiles_cached_0_probe_ready;
  wire  uncore_io_tiles_cached_0_probe_valid;
  wire [25:0] uncore_io_tiles_cached_0_probe_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_probe_bits_p_type;
  wire  uncore_io_tiles_cached_0_release_ready;
  wire  uncore_io_tiles_cached_0_release_valid;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_addr_beat;
  wire [25:0] uncore_io_tiles_cached_0_release_bits_addr_block;
  wire [1:0] uncore_io_tiles_cached_0_release_bits_client_xact_id;
  wire  uncore_io_tiles_cached_0_release_bits_voluntary;
  wire [2:0] uncore_io_tiles_cached_0_release_bits_r_type;
  wire [63:0] uncore_io_tiles_cached_0_release_bits_data;
  wire  uncore_io_tiles_cached_0_grant_ready;
  wire  uncore_io_tiles_cached_0_grant_valid;
  wire [2:0] uncore_io_tiles_cached_0_grant_bits_addr_beat;
  wire [1:0] uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_cached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_cached_0_grant_bits_data;
  wire  uncore_io_tiles_cached_0_grant_bits_manager_id;
  wire  uncore_io_tiles_cached_0_finish_ready;
  wire  uncore_io_tiles_cached_0_finish_valid;
  wire [2:0] uncore_io_tiles_cached_0_finish_bits_manager_xact_id;
  wire  uncore_io_tiles_cached_0_finish_bits_manager_id;
  wire  uncore_io_tiles_uncached_0_acquire_ready;
  wire  uncore_io_tiles_uncached_0_acquire_valid;
  wire [25:0] uncore_io_tiles_uncached_0_acquire_bits_addr_block;
  wire [1:0] uncore_io_tiles_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_addr_beat;
  wire  uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] uncore_io_tiles_uncached_0_acquire_bits_a_type;
  wire [11:0] uncore_io_tiles_uncached_0_acquire_bits_union;
  wire [63:0] uncore_io_tiles_uncached_0_acquire_bits_data;
  wire  uncore_io_tiles_uncached_0_grant_ready;
  wire  uncore_io_tiles_uncached_0_grant_valid;
  wire [2:0] uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  wire [1:0] uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  wire [2:0] uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  wire  uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] uncore_io_tiles_uncached_0_grant_bits_g_type;
  wire [63:0] uncore_io_tiles_uncached_0_grant_bits_data;
  wire  uncore_io_prci_0_reset;
  wire  uncore_io_prci_0_id;
  wire  uncore_io_prci_0_interrupts_mtip;
  wire  uncore_io_prci_0_interrupts_meip;
  wire  uncore_io_prci_0_interrupts_seip;
  wire  uncore_io_prci_0_interrupts_debug;
  wire  uncore_io_prci_0_interrupts_msip;
  wire  uncore_io_interrupts_0;
  wire  uncore_io_interrupts_1;
  wire  uncore_io_debugBus_req_ready;
  wire  uncore_io_debugBus_req_valid;
  wire [4:0] uncore_io_debugBus_req_bits_addr;
  wire [1:0] uncore_io_debugBus_req_bits_op;
  wire [33:0] uncore_io_debugBus_req_bits_data;
  wire  uncore_io_debugBus_resp_ready;
  wire  uncore_io_debugBus_resp_valid;
  wire [1:0] uncore_io_debugBus_resp_bits_resp;
  wire [33:0] uncore_io_debugBus_resp_bits_data;
  wire  RocketTile_1325_clk;
  wire  RocketTile_1325_reset;
  wire  RocketTile_1325_io_cached_0_acquire_ready;
  wire  RocketTile_1325_io_cached_0_acquire_valid;
  wire [25:0] RocketTile_1325_io_cached_0_acquire_bits_addr_block;
  wire [1:0] RocketTile_1325_io_cached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1325_io_cached_0_acquire_bits_addr_beat;
  wire  RocketTile_1325_io_cached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1325_io_cached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1325_io_cached_0_acquire_bits_union;
  wire [63:0] RocketTile_1325_io_cached_0_acquire_bits_data;
  wire  RocketTile_1325_io_cached_0_probe_ready;
  wire  RocketTile_1325_io_cached_0_probe_valid;
  wire [25:0] RocketTile_1325_io_cached_0_probe_bits_addr_block;
  wire [1:0] RocketTile_1325_io_cached_0_probe_bits_p_type;
  wire  RocketTile_1325_io_cached_0_release_ready;
  wire  RocketTile_1325_io_cached_0_release_valid;
  wire [2:0] RocketTile_1325_io_cached_0_release_bits_addr_beat;
  wire [25:0] RocketTile_1325_io_cached_0_release_bits_addr_block;
  wire [1:0] RocketTile_1325_io_cached_0_release_bits_client_xact_id;
  wire  RocketTile_1325_io_cached_0_release_bits_voluntary;
  wire [2:0] RocketTile_1325_io_cached_0_release_bits_r_type;
  wire [63:0] RocketTile_1325_io_cached_0_release_bits_data;
  wire  RocketTile_1325_io_cached_0_grant_ready;
  wire  RocketTile_1325_io_cached_0_grant_valid;
  wire [2:0] RocketTile_1325_io_cached_0_grant_bits_addr_beat;
  wire [1:0] RocketTile_1325_io_cached_0_grant_bits_client_xact_id;
  wire [2:0] RocketTile_1325_io_cached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1325_io_cached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1325_io_cached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1325_io_cached_0_grant_bits_data;
  wire  RocketTile_1325_io_cached_0_grant_bits_manager_id;
  wire  RocketTile_1325_io_cached_0_finish_ready;
  wire  RocketTile_1325_io_cached_0_finish_valid;
  wire [2:0] RocketTile_1325_io_cached_0_finish_bits_manager_xact_id;
  wire  RocketTile_1325_io_cached_0_finish_bits_manager_id;
  wire  RocketTile_1325_io_uncached_0_acquire_ready;
  wire  RocketTile_1325_io_uncached_0_acquire_valid;
  wire [25:0] RocketTile_1325_io_uncached_0_acquire_bits_addr_block;
  wire [1:0] RocketTile_1325_io_uncached_0_acquire_bits_client_xact_id;
  wire [2:0] RocketTile_1325_io_uncached_0_acquire_bits_addr_beat;
  wire  RocketTile_1325_io_uncached_0_acquire_bits_is_builtin_type;
  wire [2:0] RocketTile_1325_io_uncached_0_acquire_bits_a_type;
  wire [11:0] RocketTile_1325_io_uncached_0_acquire_bits_union;
  wire [63:0] RocketTile_1325_io_uncached_0_acquire_bits_data;
  wire  RocketTile_1325_io_uncached_0_grant_ready;
  wire  RocketTile_1325_io_uncached_0_grant_valid;
  wire [2:0] RocketTile_1325_io_uncached_0_grant_bits_addr_beat;
  wire [1:0] RocketTile_1325_io_uncached_0_grant_bits_client_xact_id;
  wire [2:0] RocketTile_1325_io_uncached_0_grant_bits_manager_xact_id;
  wire  RocketTile_1325_io_uncached_0_grant_bits_is_builtin_type;
  wire [3:0] RocketTile_1325_io_uncached_0_grant_bits_g_type;
  wire [63:0] RocketTile_1325_io_uncached_0_grant_bits_data;
  wire  RocketTile_1325_io_prci_reset;
  wire  RocketTile_1325_io_prci_id;
  wire  RocketTile_1325_io_prci_interrupts_mtip;
  wire  RocketTile_1325_io_prci_interrupts_meip;
  wire  RocketTile_1325_io_prci_interrupts_seip;
  wire  RocketTile_1325_io_prci_interrupts_debug;
  wire  RocketTile_1325_io_prci_interrupts_msip;
  wire  RocketTile_1325_io_dma_req_ready;
  wire  RocketTile_1325_io_dma_req_valid;
  wire [1:0] RocketTile_1325_io_dma_req_bits_xact_id;
  wire  RocketTile_1325_io_dma_req_bits_client_id;
  wire [2:0] RocketTile_1325_io_dma_req_bits_cmd;
  wire [31:0] RocketTile_1325_io_dma_req_bits_source;
  wire [31:0] RocketTile_1325_io_dma_req_bits_dest;
  wire [31:0] RocketTile_1325_io_dma_req_bits_length;
  wire [1:0] RocketTile_1325_io_dma_req_bits_size;
  wire  RocketTile_1325_io_dma_resp_ready;
  wire  RocketTile_1325_io_dma_resp_valid;
  wire [1:0] RocketTile_1325_io_dma_resp_bits_xact_id;
  wire  RocketTile_1325_io_dma_resp_bits_client_id;
  wire [1:0] RocketTile_1325_io_dma_resp_bits_status;
  reg  GEN_0;
  reg [31:0] GEN_5;
  reg  GEN_1;
  reg [31:0] GEN_6;
  reg [1:0] GEN_2;
  reg [31:0] GEN_7;
  reg  GEN_3;
  reg [31:0] GEN_8;
  reg [1:0] GEN_4;
  reg [31:0] GEN_9;
  Uncore uncore (
    .clk(uncore_clk),
    .reset(uncore_reset),
    .io_host_clk(uncore_io_host_clk),
    .io_host_clk_edge(uncore_io_host_clk_edge),
    .io_host_in_ready(uncore_io_host_in_ready),
    .io_host_in_valid(uncore_io_host_in_valid),
    .io_host_in_bits(uncore_io_host_in_bits),
    .io_host_out_ready(uncore_io_host_out_ready),
    .io_host_out_valid(uncore_io_host_out_valid),
    .io_host_out_bits(uncore_io_host_out_bits),
    .io_mem_axi_0_aw_ready(uncore_io_mem_axi_0_aw_ready),
    .io_mem_axi_0_aw_valid(uncore_io_mem_axi_0_aw_valid),
    .io_mem_axi_0_aw_bits_addr(uncore_io_mem_axi_0_aw_bits_addr),
    .io_mem_axi_0_aw_bits_len(uncore_io_mem_axi_0_aw_bits_len),
    .io_mem_axi_0_aw_bits_size(uncore_io_mem_axi_0_aw_bits_size),
    .io_mem_axi_0_aw_bits_burst(uncore_io_mem_axi_0_aw_bits_burst),
    .io_mem_axi_0_aw_bits_lock(uncore_io_mem_axi_0_aw_bits_lock),
    .io_mem_axi_0_aw_bits_cache(uncore_io_mem_axi_0_aw_bits_cache),
    .io_mem_axi_0_aw_bits_prot(uncore_io_mem_axi_0_aw_bits_prot),
    .io_mem_axi_0_aw_bits_qos(uncore_io_mem_axi_0_aw_bits_qos),
    .io_mem_axi_0_aw_bits_region(uncore_io_mem_axi_0_aw_bits_region),
    .io_mem_axi_0_aw_bits_id(uncore_io_mem_axi_0_aw_bits_id),
    .io_mem_axi_0_aw_bits_user(uncore_io_mem_axi_0_aw_bits_user),
    .io_mem_axi_0_w_ready(uncore_io_mem_axi_0_w_ready),
    .io_mem_axi_0_w_valid(uncore_io_mem_axi_0_w_valid),
    .io_mem_axi_0_w_bits_data(uncore_io_mem_axi_0_w_bits_data),
    .io_mem_axi_0_w_bits_last(uncore_io_mem_axi_0_w_bits_last),
    .io_mem_axi_0_w_bits_id(uncore_io_mem_axi_0_w_bits_id),
    .io_mem_axi_0_w_bits_strb(uncore_io_mem_axi_0_w_bits_strb),
    .io_mem_axi_0_w_bits_user(uncore_io_mem_axi_0_w_bits_user),
    .io_mem_axi_0_b_ready(uncore_io_mem_axi_0_b_ready),
    .io_mem_axi_0_b_valid(uncore_io_mem_axi_0_b_valid),
    .io_mem_axi_0_b_bits_resp(uncore_io_mem_axi_0_b_bits_resp),
    .io_mem_axi_0_b_bits_id(uncore_io_mem_axi_0_b_bits_id),
    .io_mem_axi_0_b_bits_user(uncore_io_mem_axi_0_b_bits_user),
    .io_mem_axi_0_ar_ready(uncore_io_mem_axi_0_ar_ready),
    .io_mem_axi_0_ar_valid(uncore_io_mem_axi_0_ar_valid),
    .io_mem_axi_0_ar_bits_addr(uncore_io_mem_axi_0_ar_bits_addr),
    .io_mem_axi_0_ar_bits_len(uncore_io_mem_axi_0_ar_bits_len),
    .io_mem_axi_0_ar_bits_size(uncore_io_mem_axi_0_ar_bits_size),
    .io_mem_axi_0_ar_bits_burst(uncore_io_mem_axi_0_ar_bits_burst),
    .io_mem_axi_0_ar_bits_lock(uncore_io_mem_axi_0_ar_bits_lock),
    .io_mem_axi_0_ar_bits_cache(uncore_io_mem_axi_0_ar_bits_cache),
    .io_mem_axi_0_ar_bits_prot(uncore_io_mem_axi_0_ar_bits_prot),
    .io_mem_axi_0_ar_bits_qos(uncore_io_mem_axi_0_ar_bits_qos),
    .io_mem_axi_0_ar_bits_region(uncore_io_mem_axi_0_ar_bits_region),
    .io_mem_axi_0_ar_bits_id(uncore_io_mem_axi_0_ar_bits_id),
    .io_mem_axi_0_ar_bits_user(uncore_io_mem_axi_0_ar_bits_user),
    .io_mem_axi_0_r_ready(uncore_io_mem_axi_0_r_ready),
    .io_mem_axi_0_r_valid(uncore_io_mem_axi_0_r_valid),
    .io_mem_axi_0_r_bits_resp(uncore_io_mem_axi_0_r_bits_resp),
    .io_mem_axi_0_r_bits_data(uncore_io_mem_axi_0_r_bits_data),
    .io_mem_axi_0_r_bits_last(uncore_io_mem_axi_0_r_bits_last),
    .io_mem_axi_0_r_bits_id(uncore_io_mem_axi_0_r_bits_id),
    .io_mem_axi_0_r_bits_user(uncore_io_mem_axi_0_r_bits_user),
    .io_tiles_cached_0_acquire_ready(uncore_io_tiles_cached_0_acquire_ready),
    .io_tiles_cached_0_acquire_valid(uncore_io_tiles_cached_0_acquire_valid),
    .io_tiles_cached_0_acquire_bits_addr_block(uncore_io_tiles_cached_0_acquire_bits_addr_block),
    .io_tiles_cached_0_acquire_bits_client_xact_id(uncore_io_tiles_cached_0_acquire_bits_client_xact_id),
    .io_tiles_cached_0_acquire_bits_addr_beat(uncore_io_tiles_cached_0_acquire_bits_addr_beat),
    .io_tiles_cached_0_acquire_bits_is_builtin_type(uncore_io_tiles_cached_0_acquire_bits_is_builtin_type),
    .io_tiles_cached_0_acquire_bits_a_type(uncore_io_tiles_cached_0_acquire_bits_a_type),
    .io_tiles_cached_0_acquire_bits_union(uncore_io_tiles_cached_0_acquire_bits_union),
    .io_tiles_cached_0_acquire_bits_data(uncore_io_tiles_cached_0_acquire_bits_data),
    .io_tiles_cached_0_probe_ready(uncore_io_tiles_cached_0_probe_ready),
    .io_tiles_cached_0_probe_valid(uncore_io_tiles_cached_0_probe_valid),
    .io_tiles_cached_0_probe_bits_addr_block(uncore_io_tiles_cached_0_probe_bits_addr_block),
    .io_tiles_cached_0_probe_bits_p_type(uncore_io_tiles_cached_0_probe_bits_p_type),
    .io_tiles_cached_0_release_ready(uncore_io_tiles_cached_0_release_ready),
    .io_tiles_cached_0_release_valid(uncore_io_tiles_cached_0_release_valid),
    .io_tiles_cached_0_release_bits_addr_beat(uncore_io_tiles_cached_0_release_bits_addr_beat),
    .io_tiles_cached_0_release_bits_addr_block(uncore_io_tiles_cached_0_release_bits_addr_block),
    .io_tiles_cached_0_release_bits_client_xact_id(uncore_io_tiles_cached_0_release_bits_client_xact_id),
    .io_tiles_cached_0_release_bits_voluntary(uncore_io_tiles_cached_0_release_bits_voluntary),
    .io_tiles_cached_0_release_bits_r_type(uncore_io_tiles_cached_0_release_bits_r_type),
    .io_tiles_cached_0_release_bits_data(uncore_io_tiles_cached_0_release_bits_data),
    .io_tiles_cached_0_grant_ready(uncore_io_tiles_cached_0_grant_ready),
    .io_tiles_cached_0_grant_valid(uncore_io_tiles_cached_0_grant_valid),
    .io_tiles_cached_0_grant_bits_addr_beat(uncore_io_tiles_cached_0_grant_bits_addr_beat),
    .io_tiles_cached_0_grant_bits_client_xact_id(uncore_io_tiles_cached_0_grant_bits_client_xact_id),
    .io_tiles_cached_0_grant_bits_manager_xact_id(uncore_io_tiles_cached_0_grant_bits_manager_xact_id),
    .io_tiles_cached_0_grant_bits_is_builtin_type(uncore_io_tiles_cached_0_grant_bits_is_builtin_type),
    .io_tiles_cached_0_grant_bits_g_type(uncore_io_tiles_cached_0_grant_bits_g_type),
    .io_tiles_cached_0_grant_bits_data(uncore_io_tiles_cached_0_grant_bits_data),
    .io_tiles_cached_0_grant_bits_manager_id(uncore_io_tiles_cached_0_grant_bits_manager_id),
    .io_tiles_cached_0_finish_ready(uncore_io_tiles_cached_0_finish_ready),
    .io_tiles_cached_0_finish_valid(uncore_io_tiles_cached_0_finish_valid),
    .io_tiles_cached_0_finish_bits_manager_xact_id(uncore_io_tiles_cached_0_finish_bits_manager_xact_id),
    .io_tiles_cached_0_finish_bits_manager_id(uncore_io_tiles_cached_0_finish_bits_manager_id),
    .io_tiles_uncached_0_acquire_ready(uncore_io_tiles_uncached_0_acquire_ready),
    .io_tiles_uncached_0_acquire_valid(uncore_io_tiles_uncached_0_acquire_valid),
    .io_tiles_uncached_0_acquire_bits_addr_block(uncore_io_tiles_uncached_0_acquire_bits_addr_block),
    .io_tiles_uncached_0_acquire_bits_client_xact_id(uncore_io_tiles_uncached_0_acquire_bits_client_xact_id),
    .io_tiles_uncached_0_acquire_bits_addr_beat(uncore_io_tiles_uncached_0_acquire_bits_addr_beat),
    .io_tiles_uncached_0_acquire_bits_is_builtin_type(uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type),
    .io_tiles_uncached_0_acquire_bits_a_type(uncore_io_tiles_uncached_0_acquire_bits_a_type),
    .io_tiles_uncached_0_acquire_bits_union(uncore_io_tiles_uncached_0_acquire_bits_union),
    .io_tiles_uncached_0_acquire_bits_data(uncore_io_tiles_uncached_0_acquire_bits_data),
    .io_tiles_uncached_0_grant_ready(uncore_io_tiles_uncached_0_grant_ready),
    .io_tiles_uncached_0_grant_valid(uncore_io_tiles_uncached_0_grant_valid),
    .io_tiles_uncached_0_grant_bits_addr_beat(uncore_io_tiles_uncached_0_grant_bits_addr_beat),
    .io_tiles_uncached_0_grant_bits_client_xact_id(uncore_io_tiles_uncached_0_grant_bits_client_xact_id),
    .io_tiles_uncached_0_grant_bits_manager_xact_id(uncore_io_tiles_uncached_0_grant_bits_manager_xact_id),
    .io_tiles_uncached_0_grant_bits_is_builtin_type(uncore_io_tiles_uncached_0_grant_bits_is_builtin_type),
    .io_tiles_uncached_0_grant_bits_g_type(uncore_io_tiles_uncached_0_grant_bits_g_type),
    .io_tiles_uncached_0_grant_bits_data(uncore_io_tiles_uncached_0_grant_bits_data),
    .io_prci_0_reset(uncore_io_prci_0_reset),
    .io_prci_0_id(uncore_io_prci_0_id),
    .io_prci_0_interrupts_mtip(uncore_io_prci_0_interrupts_mtip),
    .io_prci_0_interrupts_meip(uncore_io_prci_0_interrupts_meip),
    .io_prci_0_interrupts_seip(uncore_io_prci_0_interrupts_seip),
    .io_prci_0_interrupts_debug(uncore_io_prci_0_interrupts_debug),
    .io_prci_0_interrupts_msip(uncore_io_prci_0_interrupts_msip),
    .io_interrupts_0(uncore_io_interrupts_0),
    .io_interrupts_1(uncore_io_interrupts_1),
    .io_debugBus_req_ready(uncore_io_debugBus_req_ready),
    .io_debugBus_req_valid(uncore_io_debugBus_req_valid),
    .io_debugBus_req_bits_addr(uncore_io_debugBus_req_bits_addr),
    .io_debugBus_req_bits_op(uncore_io_debugBus_req_bits_op),
    .io_debugBus_req_bits_data(uncore_io_debugBus_req_bits_data),
    .io_debugBus_resp_ready(uncore_io_debugBus_resp_ready),
    .io_debugBus_resp_valid(uncore_io_debugBus_resp_valid),
    .io_debugBus_resp_bits_resp(uncore_io_debugBus_resp_bits_resp),
    .io_debugBus_resp_bits_data(uncore_io_debugBus_resp_bits_data)
  );
  RocketTile RocketTile_1325 (
    .clk(RocketTile_1325_clk),
    .reset(RocketTile_1325_reset),
    .io_cached_0_acquire_ready(RocketTile_1325_io_cached_0_acquire_ready),
    .io_cached_0_acquire_valid(RocketTile_1325_io_cached_0_acquire_valid),
    .io_cached_0_acquire_bits_addr_block(RocketTile_1325_io_cached_0_acquire_bits_addr_block),
    .io_cached_0_acquire_bits_client_xact_id(RocketTile_1325_io_cached_0_acquire_bits_client_xact_id),
    .io_cached_0_acquire_bits_addr_beat(RocketTile_1325_io_cached_0_acquire_bits_addr_beat),
    .io_cached_0_acquire_bits_is_builtin_type(RocketTile_1325_io_cached_0_acquire_bits_is_builtin_type),
    .io_cached_0_acquire_bits_a_type(RocketTile_1325_io_cached_0_acquire_bits_a_type),
    .io_cached_0_acquire_bits_union(RocketTile_1325_io_cached_0_acquire_bits_union),
    .io_cached_0_acquire_bits_data(RocketTile_1325_io_cached_0_acquire_bits_data),
    .io_cached_0_probe_ready(RocketTile_1325_io_cached_0_probe_ready),
    .io_cached_0_probe_valid(RocketTile_1325_io_cached_0_probe_valid),
    .io_cached_0_probe_bits_addr_block(RocketTile_1325_io_cached_0_probe_bits_addr_block),
    .io_cached_0_probe_bits_p_type(RocketTile_1325_io_cached_0_probe_bits_p_type),
    .io_cached_0_release_ready(RocketTile_1325_io_cached_0_release_ready),
    .io_cached_0_release_valid(RocketTile_1325_io_cached_0_release_valid),
    .io_cached_0_release_bits_addr_beat(RocketTile_1325_io_cached_0_release_bits_addr_beat),
    .io_cached_0_release_bits_addr_block(RocketTile_1325_io_cached_0_release_bits_addr_block),
    .io_cached_0_release_bits_client_xact_id(RocketTile_1325_io_cached_0_release_bits_client_xact_id),
    .io_cached_0_release_bits_voluntary(RocketTile_1325_io_cached_0_release_bits_voluntary),
    .io_cached_0_release_bits_r_type(RocketTile_1325_io_cached_0_release_bits_r_type),
    .io_cached_0_release_bits_data(RocketTile_1325_io_cached_0_release_bits_data),
    .io_cached_0_grant_ready(RocketTile_1325_io_cached_0_grant_ready),
    .io_cached_0_grant_valid(RocketTile_1325_io_cached_0_grant_valid),
    .io_cached_0_grant_bits_addr_beat(RocketTile_1325_io_cached_0_grant_bits_addr_beat),
    .io_cached_0_grant_bits_client_xact_id(RocketTile_1325_io_cached_0_grant_bits_client_xact_id),
    .io_cached_0_grant_bits_manager_xact_id(RocketTile_1325_io_cached_0_grant_bits_manager_xact_id),
    .io_cached_0_grant_bits_is_builtin_type(RocketTile_1325_io_cached_0_grant_bits_is_builtin_type),
    .io_cached_0_grant_bits_g_type(RocketTile_1325_io_cached_0_grant_bits_g_type),
    .io_cached_0_grant_bits_data(RocketTile_1325_io_cached_0_grant_bits_data),
    .io_cached_0_grant_bits_manager_id(RocketTile_1325_io_cached_0_grant_bits_manager_id),
    .io_cached_0_finish_ready(RocketTile_1325_io_cached_0_finish_ready),
    .io_cached_0_finish_valid(RocketTile_1325_io_cached_0_finish_valid),
    .io_cached_0_finish_bits_manager_xact_id(RocketTile_1325_io_cached_0_finish_bits_manager_xact_id),
    .io_cached_0_finish_bits_manager_id(RocketTile_1325_io_cached_0_finish_bits_manager_id),
    .io_uncached_0_acquire_ready(RocketTile_1325_io_uncached_0_acquire_ready),
    .io_uncached_0_acquire_valid(RocketTile_1325_io_uncached_0_acquire_valid),
    .io_uncached_0_acquire_bits_addr_block(RocketTile_1325_io_uncached_0_acquire_bits_addr_block),
    .io_uncached_0_acquire_bits_client_xact_id(RocketTile_1325_io_uncached_0_acquire_bits_client_xact_id),
    .io_uncached_0_acquire_bits_addr_beat(RocketTile_1325_io_uncached_0_acquire_bits_addr_beat),
    .io_uncached_0_acquire_bits_is_builtin_type(RocketTile_1325_io_uncached_0_acquire_bits_is_builtin_type),
    .io_uncached_0_acquire_bits_a_type(RocketTile_1325_io_uncached_0_acquire_bits_a_type),
    .io_uncached_0_acquire_bits_union(RocketTile_1325_io_uncached_0_acquire_bits_union),
    .io_uncached_0_acquire_bits_data(RocketTile_1325_io_uncached_0_acquire_bits_data),
    .io_uncached_0_grant_ready(RocketTile_1325_io_uncached_0_grant_ready),
    .io_uncached_0_grant_valid(RocketTile_1325_io_uncached_0_grant_valid),
    .io_uncached_0_grant_bits_addr_beat(RocketTile_1325_io_uncached_0_grant_bits_addr_beat),
    .io_uncached_0_grant_bits_client_xact_id(RocketTile_1325_io_uncached_0_grant_bits_client_xact_id),
    .io_uncached_0_grant_bits_manager_xact_id(RocketTile_1325_io_uncached_0_grant_bits_manager_xact_id),
    .io_uncached_0_grant_bits_is_builtin_type(RocketTile_1325_io_uncached_0_grant_bits_is_builtin_type),
    .io_uncached_0_grant_bits_g_type(RocketTile_1325_io_uncached_0_grant_bits_g_type),
    .io_uncached_0_grant_bits_data(RocketTile_1325_io_uncached_0_grant_bits_data),
    .io_prci_reset(RocketTile_1325_io_prci_reset),
    .io_prci_id(RocketTile_1325_io_prci_id),
    .io_prci_interrupts_mtip(RocketTile_1325_io_prci_interrupts_mtip),
    .io_prci_interrupts_meip(RocketTile_1325_io_prci_interrupts_meip),
    .io_prci_interrupts_seip(RocketTile_1325_io_prci_interrupts_seip),
    .io_prci_interrupts_debug(RocketTile_1325_io_prci_interrupts_debug),
    .io_prci_interrupts_msip(RocketTile_1325_io_prci_interrupts_msip),
    .io_dma_req_ready(RocketTile_1325_io_dma_req_ready),
    .io_dma_req_valid(RocketTile_1325_io_dma_req_valid),
    .io_dma_req_bits_xact_id(RocketTile_1325_io_dma_req_bits_xact_id),
    .io_dma_req_bits_client_id(RocketTile_1325_io_dma_req_bits_client_id),
    .io_dma_req_bits_cmd(RocketTile_1325_io_dma_req_bits_cmd),
    .io_dma_req_bits_source(RocketTile_1325_io_dma_req_bits_source),
    .io_dma_req_bits_dest(RocketTile_1325_io_dma_req_bits_dest),
    .io_dma_req_bits_length(RocketTile_1325_io_dma_req_bits_length),
    .io_dma_req_bits_size(RocketTile_1325_io_dma_req_bits_size),
    .io_dma_resp_ready(RocketTile_1325_io_dma_resp_ready),
    .io_dma_resp_valid(RocketTile_1325_io_dma_resp_valid),
    .io_dma_resp_bits_xact_id(RocketTile_1325_io_dma_resp_bits_xact_id),
    .io_dma_resp_bits_client_id(RocketTile_1325_io_dma_resp_bits_client_id),
    .io_dma_resp_bits_status(RocketTile_1325_io_dma_resp_bits_status)
  );
  assign io_host_clk = uncore_io_host_clk;
  assign io_host_clk_edge = uncore_io_host_clk_edge;
  assign io_host_in_ready = uncore_io_host_in_ready;
  assign io_host_out_valid = uncore_io_host_out_valid;
  assign io_host_out_bits = uncore_io_host_out_bits;
  assign io_mem_axi_0_aw_valid = uncore_io_mem_axi_0_aw_valid;
  assign io_mem_axi_0_aw_bits_addr = uncore_io_mem_axi_0_aw_bits_addr;
  assign io_mem_axi_0_aw_bits_len = uncore_io_mem_axi_0_aw_bits_len;
  assign io_mem_axi_0_aw_bits_size = uncore_io_mem_axi_0_aw_bits_size;
  assign io_mem_axi_0_aw_bits_burst = uncore_io_mem_axi_0_aw_bits_burst;
  assign io_mem_axi_0_aw_bits_lock = uncore_io_mem_axi_0_aw_bits_lock;
  assign io_mem_axi_0_aw_bits_cache = uncore_io_mem_axi_0_aw_bits_cache;
  assign io_mem_axi_0_aw_bits_prot = uncore_io_mem_axi_0_aw_bits_prot;
  assign io_mem_axi_0_aw_bits_qos = uncore_io_mem_axi_0_aw_bits_qos;
  assign io_mem_axi_0_aw_bits_region = uncore_io_mem_axi_0_aw_bits_region;
  assign io_mem_axi_0_aw_bits_id = uncore_io_mem_axi_0_aw_bits_id;
  assign io_mem_axi_0_aw_bits_user = uncore_io_mem_axi_0_aw_bits_user;
  assign io_mem_axi_0_w_valid = uncore_io_mem_axi_0_w_valid;
  assign io_mem_axi_0_w_bits_data = uncore_io_mem_axi_0_w_bits_data;
  assign io_mem_axi_0_w_bits_last = uncore_io_mem_axi_0_w_bits_last;
  assign io_mem_axi_0_w_bits_id = uncore_io_mem_axi_0_w_bits_id;
  assign io_mem_axi_0_w_bits_strb = uncore_io_mem_axi_0_w_bits_strb;
  assign io_mem_axi_0_w_bits_user = uncore_io_mem_axi_0_w_bits_user;
  assign io_mem_axi_0_b_ready = uncore_io_mem_axi_0_b_ready;
  assign io_mem_axi_0_ar_valid = uncore_io_mem_axi_0_ar_valid;
  assign io_mem_axi_0_ar_bits_addr = uncore_io_mem_axi_0_ar_bits_addr;
  assign io_mem_axi_0_ar_bits_len = uncore_io_mem_axi_0_ar_bits_len;
  assign io_mem_axi_0_ar_bits_size = uncore_io_mem_axi_0_ar_bits_size;
  assign io_mem_axi_0_ar_bits_burst = uncore_io_mem_axi_0_ar_bits_burst;
  assign io_mem_axi_0_ar_bits_lock = uncore_io_mem_axi_0_ar_bits_lock;
  assign io_mem_axi_0_ar_bits_cache = uncore_io_mem_axi_0_ar_bits_cache;
  assign io_mem_axi_0_ar_bits_prot = uncore_io_mem_axi_0_ar_bits_prot;
  assign io_mem_axi_0_ar_bits_qos = uncore_io_mem_axi_0_ar_bits_qos;
  assign io_mem_axi_0_ar_bits_region = uncore_io_mem_axi_0_ar_bits_region;
  assign io_mem_axi_0_ar_bits_id = uncore_io_mem_axi_0_ar_bits_id;
  assign io_mem_axi_0_ar_bits_user = uncore_io_mem_axi_0_ar_bits_user;
  assign io_mem_axi_0_r_ready = uncore_io_mem_axi_0_r_ready;
  assign io_debug_req_ready = uncore_io_debugBus_req_ready;
  assign io_debug_resp_valid = uncore_io_debugBus_resp_valid;
  assign io_debug_resp_bits_resp = uncore_io_debugBus_resp_bits_resp;
  assign io_debug_resp_bits_data = uncore_io_debugBus_resp_bits_data;
  assign uncore_clk = clk;
  assign uncore_reset = reset;
  assign uncore_io_host_in_valid = io_host_in_valid;
  assign uncore_io_host_in_bits = io_host_in_bits;
  assign uncore_io_host_out_ready = io_host_out_ready;
  assign uncore_io_mem_axi_0_aw_ready = io_mem_axi_0_aw_ready;
  assign uncore_io_mem_axi_0_w_ready = io_mem_axi_0_w_ready;
  assign uncore_io_mem_axi_0_b_valid = io_mem_axi_0_b_valid;
  assign uncore_io_mem_axi_0_b_bits_resp = io_mem_axi_0_b_bits_resp;
  assign uncore_io_mem_axi_0_b_bits_id = io_mem_axi_0_b_bits_id;
  assign uncore_io_mem_axi_0_b_bits_user = io_mem_axi_0_b_bits_user;
  assign uncore_io_mem_axi_0_ar_ready = io_mem_axi_0_ar_ready;
  assign uncore_io_mem_axi_0_r_valid = io_mem_axi_0_r_valid;
  assign uncore_io_mem_axi_0_r_bits_resp = io_mem_axi_0_r_bits_resp;
  assign uncore_io_mem_axi_0_r_bits_data = io_mem_axi_0_r_bits_data;
  assign uncore_io_mem_axi_0_r_bits_last = io_mem_axi_0_r_bits_last;
  assign uncore_io_mem_axi_0_r_bits_id = io_mem_axi_0_r_bits_id;
  assign uncore_io_mem_axi_0_r_bits_user = io_mem_axi_0_r_bits_user;
  assign uncore_io_tiles_cached_0_acquire_valid = RocketTile_1325_io_cached_0_acquire_valid;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_block = RocketTile_1325_io_cached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_cached_0_acquire_bits_client_xact_id = RocketTile_1325_io_cached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_acquire_bits_addr_beat = RocketTile_1325_io_cached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_cached_0_acquire_bits_is_builtin_type = RocketTile_1325_io_cached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_cached_0_acquire_bits_a_type = RocketTile_1325_io_cached_0_acquire_bits_a_type;
  assign uncore_io_tiles_cached_0_acquire_bits_union = RocketTile_1325_io_cached_0_acquire_bits_union;
  assign uncore_io_tiles_cached_0_acquire_bits_data = RocketTile_1325_io_cached_0_acquire_bits_data;
  assign uncore_io_tiles_cached_0_probe_ready = RocketTile_1325_io_cached_0_probe_ready;
  assign uncore_io_tiles_cached_0_release_valid = RocketTile_1325_io_cached_0_release_valid;
  assign uncore_io_tiles_cached_0_release_bits_addr_beat = RocketTile_1325_io_cached_0_release_bits_addr_beat;
  assign uncore_io_tiles_cached_0_release_bits_addr_block = RocketTile_1325_io_cached_0_release_bits_addr_block;
  assign uncore_io_tiles_cached_0_release_bits_client_xact_id = RocketTile_1325_io_cached_0_release_bits_client_xact_id;
  assign uncore_io_tiles_cached_0_release_bits_voluntary = RocketTile_1325_io_cached_0_release_bits_voluntary;
  assign uncore_io_tiles_cached_0_release_bits_r_type = RocketTile_1325_io_cached_0_release_bits_r_type;
  assign uncore_io_tiles_cached_0_release_bits_data = RocketTile_1325_io_cached_0_release_bits_data;
  assign uncore_io_tiles_cached_0_grant_ready = RocketTile_1325_io_cached_0_grant_ready;
  assign uncore_io_tiles_cached_0_finish_valid = RocketTile_1325_io_cached_0_finish_valid;
  assign uncore_io_tiles_cached_0_finish_bits_manager_xact_id = RocketTile_1325_io_cached_0_finish_bits_manager_xact_id;
  assign uncore_io_tiles_cached_0_finish_bits_manager_id = RocketTile_1325_io_cached_0_finish_bits_manager_id;
  assign uncore_io_tiles_uncached_0_acquire_valid = RocketTile_1325_io_uncached_0_acquire_valid;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_block = RocketTile_1325_io_uncached_0_acquire_bits_addr_block;
  assign uncore_io_tiles_uncached_0_acquire_bits_client_xact_id = RocketTile_1325_io_uncached_0_acquire_bits_client_xact_id;
  assign uncore_io_tiles_uncached_0_acquire_bits_addr_beat = RocketTile_1325_io_uncached_0_acquire_bits_addr_beat;
  assign uncore_io_tiles_uncached_0_acquire_bits_is_builtin_type = RocketTile_1325_io_uncached_0_acquire_bits_is_builtin_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_a_type = RocketTile_1325_io_uncached_0_acquire_bits_a_type;
  assign uncore_io_tiles_uncached_0_acquire_bits_union = RocketTile_1325_io_uncached_0_acquire_bits_union;
  assign uncore_io_tiles_uncached_0_acquire_bits_data = RocketTile_1325_io_uncached_0_acquire_bits_data;
  assign uncore_io_tiles_uncached_0_grant_ready = RocketTile_1325_io_uncached_0_grant_ready;
  assign uncore_io_interrupts_0 = io_interrupts_0;
  assign uncore_io_interrupts_1 = io_interrupts_1;
  assign uncore_io_debugBus_req_valid = io_debug_req_valid;
  assign uncore_io_debugBus_req_bits_addr = io_debug_req_bits_addr;
  assign uncore_io_debugBus_req_bits_op = io_debug_req_bits_op;
  assign uncore_io_debugBus_req_bits_data = io_debug_req_bits_data;
  assign uncore_io_debugBus_resp_ready = io_debug_resp_ready;
  assign RocketTile_1325_clk = clk;
  assign RocketTile_1325_reset = uncore_io_prci_0_reset;
  assign RocketTile_1325_io_cached_0_acquire_ready = uncore_io_tiles_cached_0_acquire_ready;
  assign RocketTile_1325_io_cached_0_probe_valid = uncore_io_tiles_cached_0_probe_valid;
  assign RocketTile_1325_io_cached_0_probe_bits_addr_block = uncore_io_tiles_cached_0_probe_bits_addr_block;
  assign RocketTile_1325_io_cached_0_probe_bits_p_type = uncore_io_tiles_cached_0_probe_bits_p_type;
  assign RocketTile_1325_io_cached_0_release_ready = uncore_io_tiles_cached_0_release_ready;
  assign RocketTile_1325_io_cached_0_grant_valid = uncore_io_tiles_cached_0_grant_valid;
  assign RocketTile_1325_io_cached_0_grant_bits_addr_beat = uncore_io_tiles_cached_0_grant_bits_addr_beat;
  assign RocketTile_1325_io_cached_0_grant_bits_client_xact_id = uncore_io_tiles_cached_0_grant_bits_client_xact_id;
  assign RocketTile_1325_io_cached_0_grant_bits_manager_xact_id = uncore_io_tiles_cached_0_grant_bits_manager_xact_id;
  assign RocketTile_1325_io_cached_0_grant_bits_is_builtin_type = uncore_io_tiles_cached_0_grant_bits_is_builtin_type;
  assign RocketTile_1325_io_cached_0_grant_bits_g_type = uncore_io_tiles_cached_0_grant_bits_g_type;
  assign RocketTile_1325_io_cached_0_grant_bits_data = uncore_io_tiles_cached_0_grant_bits_data;
  assign RocketTile_1325_io_cached_0_grant_bits_manager_id = uncore_io_tiles_cached_0_grant_bits_manager_id;
  assign RocketTile_1325_io_cached_0_finish_ready = uncore_io_tiles_cached_0_finish_ready;
  assign RocketTile_1325_io_uncached_0_acquire_ready = uncore_io_tiles_uncached_0_acquire_ready;
  assign RocketTile_1325_io_uncached_0_grant_valid = uncore_io_tiles_uncached_0_grant_valid;
  assign RocketTile_1325_io_uncached_0_grant_bits_addr_beat = uncore_io_tiles_uncached_0_grant_bits_addr_beat;
  assign RocketTile_1325_io_uncached_0_grant_bits_client_xact_id = uncore_io_tiles_uncached_0_grant_bits_client_xact_id;
  assign RocketTile_1325_io_uncached_0_grant_bits_manager_xact_id = uncore_io_tiles_uncached_0_grant_bits_manager_xact_id;
  assign RocketTile_1325_io_uncached_0_grant_bits_is_builtin_type = uncore_io_tiles_uncached_0_grant_bits_is_builtin_type;
  assign RocketTile_1325_io_uncached_0_grant_bits_g_type = uncore_io_tiles_uncached_0_grant_bits_g_type;
  assign RocketTile_1325_io_uncached_0_grant_bits_data = uncore_io_tiles_uncached_0_grant_bits_data;
  assign RocketTile_1325_io_prci_reset = uncore_io_prci_0_reset;
  assign RocketTile_1325_io_prci_id = uncore_io_prci_0_id;
  assign RocketTile_1325_io_prci_interrupts_mtip = uncore_io_prci_0_interrupts_mtip;
  assign RocketTile_1325_io_prci_interrupts_meip = uncore_io_prci_0_interrupts_meip;
  assign RocketTile_1325_io_prci_interrupts_seip = uncore_io_prci_0_interrupts_seip;
  assign RocketTile_1325_io_prci_interrupts_debug = uncore_io_prci_0_interrupts_debug;
  assign RocketTile_1325_io_prci_interrupts_msip = uncore_io_prci_0_interrupts_msip;
  assign RocketTile_1325_io_dma_req_ready = GEN_0;
  assign RocketTile_1325_io_dma_resp_valid = GEN_1;
  assign RocketTile_1325_io_dma_resp_bits_xact_id = GEN_2;
  assign RocketTile_1325_io_dma_resp_bits_client_id = GEN_3;
  assign RocketTile_1325_io_dma_resp_bits_status = GEN_4;
`ifndef SYNTHESIS
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  GEN_5 = {1{$random}};
  GEN_0 = GEN_5[0:0];
  GEN_6 = {1{$random}};
  GEN_1 = GEN_6[0:0];
  GEN_7 = {1{$random}};
  GEN_2 = GEN_7[1:0];
  GEN_8 = {1{$random}};
  GEN_3 = GEN_8[0:0];
  GEN_9 = {1{$random}};
  GEN_4 = GEN_9[1:0];
  end
`endif
endmodule
